
module ALU_WIDTH32_RADIX4_OPCODE6 ( A, B, .OP({\OP[4] , \OP[3] , \OP[2] , 
        \OP[1] , \OP[0] }), Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input \OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] ;
  wire   s_SIGN, N21, N22, N25, N27, N28, N29, N30, N31, N33, N34, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N62, N63, N66, N67, N87, N89, N91,
         N92, \ADD_SUB/carry_ST[0] , \MULT/SHIFTERi_0/N19 , n1, n24, n26, n87,
         n88, n89, n93, n96, n105, n107, n110, n118, n119, n122, n127, n900,
         n1119, n1155, n1616, n1617, n1618, n1619, n3308, n3309, n3314, n3331,
         n3332, n3333, n3432, n4840, n4841, n4842, n4843, \intadd_0/B[7] ,
         \intadd_0/B[6] , \intadd_0/B[5] , \intadd_0/B[4] , \intadd_0/B[3] ,
         \intadd_0/B[2] , \intadd_0/B[1] , \intadd_0/B[0] , \intadd_0/CI ,
         \intadd_0/SUM[7] , \intadd_0/SUM[6] , \intadd_0/SUM[5] ,
         \intadd_0/SUM[4] , \intadd_0/SUM[3] , \intadd_0/SUM[2] ,
         \intadd_0/SUM[1] , \intadd_0/SUM[0] , \intadd_0/n8 , \intadd_0/n7 ,
         \intadd_0/n6 , \intadd_0/n5 , \intadd_0/n4 , \intadd_0/n3 ,
         \intadd_0/n2 , \intadd_0/n1 , \intadd_1/B[7] , \intadd_1/B[6] ,
         \intadd_1/B[5] , \intadd_1/B[4] , \intadd_1/B[3] , \intadd_1/B[2] ,
         \intadd_1/B[1] , \intadd_1/B[0] , \intadd_1/CI , \intadd_1/SUM[7] ,
         \intadd_1/SUM[6] , \intadd_1/SUM[5] , \intadd_1/SUM[4] ,
         \intadd_1/SUM[3] , \intadd_1/SUM[2] , \intadd_1/SUM[1] ,
         \intadd_1/SUM[0] , \intadd_1/n8 , \intadd_1/n7 , \intadd_1/n6 ,
         \intadd_1/n5 , \intadd_1/n4 , \intadd_1/n3 , \intadd_1/n2 ,
         \intadd_1/n1 , \intadd_2/A[3] , \intadd_2/A[2] , \intadd_2/A[1] ,
         \intadd_2/A[0] , \intadd_2/B[3] , \intadd_2/B[2] , \intadd_2/B[1] ,
         \intadd_2/B[0] , \intadd_2/CI , \intadd_2/SUM[3] , \intadd_2/SUM[2] ,
         \intadd_2/SUM[1] , \intadd_2/SUM[0] , \intadd_2/n4 , \intadd_2/n3 ,
         \intadd_2/n2 , \intadd_2/n1 , \intadd_3/A[3] , \intadd_3/A[2] ,
         \intadd_3/A[1] , \intadd_3/A[0] , \intadd_3/B[3] , \intadd_3/B[2] ,
         \intadd_3/B[1] , \intadd_3/B[0] , \intadd_3/CI , \intadd_3/SUM[3] ,
         \intadd_3/SUM[2] , \intadd_3/SUM[1] , \intadd_3/SUM[0] ,
         \intadd_3/n4 , \intadd_3/n3 , \intadd_3/n2 , \intadd_3/n1 ,
         \intadd_4/A[3] , \intadd_4/A[2] , \intadd_4/A[1] , \intadd_4/A[0] ,
         \intadd_4/B[3] , \intadd_4/B[2] , \intadd_4/B[1] , \intadd_4/B[0] ,
         \intadd_4/CI , \intadd_4/SUM[3] , \intadd_4/n4 , \intadd_4/n3 ,
         \intadd_4/n2 , \intadd_4/n1 , \intadd_5/A[2] , \intadd_5/A[0] ,
         \intadd_5/B[1] , \intadd_5/B[0] , \intadd_5/CI , \intadd_5/SUM[2] ,
         \intadd_5/SUM[1] , \intadd_5/SUM[0] , \intadd_5/n3 , \intadd_5/n2 ,
         \intadd_5/n1 , \intadd_6/A[2] , \intadd_6/A[1] , \intadd_6/A[0] ,
         \intadd_6/B[0] , \intadd_6/CI , \intadd_6/n3 , \intadd_6/n2 ,
         \intadd_6/n1 , \intadd_7/A[2] , \intadd_7/A[1] , \intadd_7/A[0] ,
         \intadd_7/B[2] , \intadd_7/B[1] , \intadd_7/B[0] , \intadd_7/CI ,
         \intadd_7/n3 , \intadd_7/n2 , \intadd_7/n1 , \intadd_8/A[2] ,
         \intadd_8/A[1] , \intadd_8/A[0] , \intadd_8/B[2] , \intadd_8/B[1] ,
         \intadd_8/B[0] , \intadd_8/CI , \intadd_8/SUM[2] , \intadd_8/n3 ,
         \intadd_8/n2 , \intadd_8/n1 , \intadd_9/A[1] , \intadd_9/B[2] ,
         \intadd_9/B[1] , \intadd_9/B[0] , \intadd_9/CI , \intadd_9/SUM[2] ,
         \intadd_9/n3 , \intadd_9/n2 , \intadd_9/n1 , \intadd_10/A[2] ,
         \intadd_10/A[0] , \intadd_10/B[1] , \intadd_10/B[0] , \intadd_10/CI ,
         \intadd_10/SUM[2] , \intadd_10/SUM[1] , \intadd_10/SUM[0] ,
         \intadd_10/n3 , \intadd_10/n2 , \intadd_10/n1 , \intadd_11/A[2] ,
         \intadd_11/A[1] , \intadd_11/A[0] , \intadd_11/B[2] ,
         \intadd_11/B[1] , \intadd_11/B[0] , \intadd_11/CI ,
         \intadd_11/SUM[2] , \intadd_11/SUM[1] , \intadd_11/SUM[0] ,
         \intadd_11/n3 , \intadd_11/n2 , \intadd_11/n1 , \intadd_12/A[2] ,
         \intadd_12/A[1] , \intadd_12/A[0] , \intadd_12/B[0] , \intadd_12/CI ,
         \intadd_12/SUM[2] , \intadd_12/SUM[1] , \intadd_12/SUM[0] ,
         \intadd_12/n3 , \intadd_12/n2 , \intadd_12/n1 , n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6329, n6330, n6331, n6333, n6334,
         n6336, n6337, n6339, n6346, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6451, n7619, n7620, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n14, n15, n17, n18, n19, n20, n21, n22, n23, n25, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n80, n81, n82, n83, n84, n85, n86, n90,
         n91, n92, n94, n95, n97, n98, n99, n100, n101, n102, n103, n104, n106,
         n108, n109, n111, n112, n113, n114, n115, n116, n117, n120, n121,
         n123, n124, n125, n126, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n434, n436, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n450, n451, n452, n454, n456, n457, n458, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537;
  wire   [4:0] OP;
  wire   [31:0] s_A_ADDER;
  wire   [31:0] S_B_ADDER;
  wire   [31:0] s_A_LOGIC;
  wire   [31:0] S_B_LOGIC;
  wire   [3:0] s_LOGIC;
  wire   [31:0] s_A_SHIFT;
  wire   [31:0] S_B_SHIFT;
  wire   [1:0] s_SHIFT;
  wire   [15:0] s_A_MULT;
  wire   [15:0] S_B_MULT;
  wire   [15:0] S_B_LHI;

  DLH_X1 s_SIGN_reg ( .G(N91), .D(N92), .Q(s_SIGN) );
  DLH_X1 \S_B_ADDER_reg[5]  ( .G(n80), .D(N59), .Q(S_B_ADDER[5]) );
  DLH_X1 \S_B_ADDER_reg[4]  ( .G(N21), .D(N58), .Q(S_B_ADDER[4]) );
  DLH_X1 \S_B_ADDER_reg[3]  ( .G(N21), .D(N57), .Q(S_B_ADDER[3]) );
  DLH_X1 \S_B_ADDER_reg[2]  ( .G(n80), .D(N56), .Q(S_B_ADDER[2]) );
  DLH_X1 \S_B_ADDER_reg[1]  ( .G(N21), .D(N55), .Q(S_B_ADDER[1]) );
  DLH_X1 \S_B_ADDER_reg[0]  ( .G(n80), .D(N54), .Q(S_B_ADDER[0]) );
  DLH_X1 s_ADD_SUB_reg ( .G(n80), .D(n3432), .Q(\ADD_SUB/carry_ST[0] ) );
  DLH_X1 \s_A_LOGIC_reg[31]  ( .G(n78), .D(A[31]), .Q(s_A_LOGIC[31]) );
  DLH_X1 \s_A_LOGIC_reg[30]  ( .G(n1525), .D(A[30]), .Q(s_A_LOGIC[30]) );
  DLH_X1 \s_A_LOGIC_reg[29]  ( .G(n1535), .D(A[29]), .Q(s_A_LOGIC[29]) );
  DLH_X1 \s_A_LOGIC_reg[28]  ( .G(n1535), .D(A[28]), .Q(s_A_LOGIC[28]) );
  DLH_X1 \s_A_LOGIC_reg[27]  ( .G(n78), .D(A[27]), .Q(s_A_LOGIC[27]) );
  DLH_X1 \s_A_LOGIC_reg[26]  ( .G(n1535), .D(A[26]), .Q(s_A_LOGIC[26]) );
  DLH_X1 \s_A_LOGIC_reg[25]  ( .G(n1525), .D(A[25]), .Q(s_A_LOGIC[25]) );
  DLH_X1 \s_A_LOGIC_reg[24]  ( .G(n1535), .D(A[24]), .Q(s_A_LOGIC[24]) );
  DLH_X1 \s_A_LOGIC_reg[23]  ( .G(n78), .D(A[23]), .Q(s_A_LOGIC[23]) );
  DLH_X1 \s_A_LOGIC_reg[22]  ( .G(n78), .D(A[22]), .Q(s_A_LOGIC[22]) );
  DLH_X1 \s_A_LOGIC_reg[21]  ( .G(n1535), .D(A[21]), .Q(s_A_LOGIC[21]) );
  DLH_X1 \s_A_LOGIC_reg[20]  ( .G(n1527), .D(A[20]), .Q(s_A_LOGIC[20]) );
  DLH_X1 \s_A_LOGIC_reg[19]  ( .G(n1535), .D(A[19]), .Q(s_A_LOGIC[19]) );
  DLH_X1 \s_A_LOGIC_reg[18]  ( .G(n1535), .D(A[18]), .Q(s_A_LOGIC[18]) );
  DLH_X1 \s_A_LOGIC_reg[17]  ( .G(n1525), .D(A[17]), .Q(s_A_LOGIC[17]) );
  DLH_X1 \s_A_LOGIC_reg[16]  ( .G(n1535), .D(A[16]), .Q(s_A_LOGIC[16]) );
  DLH_X1 \s_A_LOGIC_reg[15]  ( .G(n78), .D(A[15]), .Q(s_A_LOGIC[15]) );
  DLH_X1 \s_A_LOGIC_reg[14]  ( .G(n78), .D(A[14]), .Q(s_A_LOGIC[14]) );
  DLH_X1 \s_A_LOGIC_reg[13]  ( .G(n78), .D(A[13]), .Q(s_A_LOGIC[13]) );
  DLH_X1 \s_A_LOGIC_reg[12]  ( .G(n1527), .D(A[12]), .Q(s_A_LOGIC[12]) );
  DLH_X1 \s_A_LOGIC_reg[11]  ( .G(n1535), .D(A[11]), .Q(s_A_LOGIC[11]) );
  DLH_X1 \s_A_LOGIC_reg[10]  ( .G(n1535), .D(A[10]), .Q(s_A_LOGIC[10]) );
  DLH_X1 \s_A_LOGIC_reg[9]  ( .G(n1527), .D(A[9]), .Q(s_A_LOGIC[9]) );
  DLH_X1 \s_A_LOGIC_reg[8]  ( .G(n1527), .D(A[8]), .Q(s_A_LOGIC[8]) );
  DLH_X1 \s_A_LOGIC_reg[7]  ( .G(n1535), .D(A[7]), .Q(s_A_LOGIC[7]) );
  DLH_X1 \s_A_LOGIC_reg[6]  ( .G(n1527), .D(A[6]), .Q(s_A_LOGIC[6]) );
  DLH_X1 \s_A_LOGIC_reg[5]  ( .G(n1527), .D(A[5]), .Q(s_A_LOGIC[5]) );
  DLH_X1 \s_A_LOGIC_reg[4]  ( .G(n1527), .D(A[4]), .Q(s_A_LOGIC[4]) );
  DLH_X1 \s_A_LOGIC_reg[3]  ( .G(n1535), .D(A[3]), .Q(s_A_LOGIC[3]) );
  DLH_X1 \s_A_LOGIC_reg[2]  ( .G(n1527), .D(A[2]), .Q(s_A_LOGIC[2]) );
  DLH_X1 \s_A_LOGIC_reg[1]  ( .G(n1527), .D(A[1]), .Q(s_A_LOGIC[1]) );
  DLH_X1 \s_A_LOGIC_reg[0]  ( .G(n78), .D(A[0]), .Q(s_A_LOGIC[0]) );
  DLH_X1 \S_B_LOGIC_reg[31]  ( .G(n1535), .D(B[31]), .Q(S_B_LOGIC[31]) );
  DLH_X1 \S_B_LOGIC_reg[30]  ( .G(n1535), .D(B[30]), .Q(S_B_LOGIC[30]) );
  DLH_X1 \S_B_LOGIC_reg[29]  ( .G(n78), .D(B[29]), .Q(S_B_LOGIC[29]) );
  DLH_X1 \S_B_LOGIC_reg[28]  ( .G(n78), .D(B[28]), .Q(S_B_LOGIC[28]) );
  DLH_X1 \S_B_LOGIC_reg[27]  ( .G(n1527), .D(B[27]), .Q(S_B_LOGIC[27]) );
  DLH_X1 \S_B_LOGIC_reg[26]  ( .G(n1527), .D(B[26]), .Q(S_B_LOGIC[26]) );
  DLH_X1 \S_B_LOGIC_reg[25]  ( .G(n78), .D(B[25]), .Q(S_B_LOGIC[25]) );
  DLH_X1 \S_B_LOGIC_reg[24]  ( .G(n78), .D(B[24]), .Q(S_B_LOGIC[24]) );
  DLH_X1 \S_B_LOGIC_reg[23]  ( .G(n1527), .D(B[23]), .Q(S_B_LOGIC[23]) );
  DLH_X1 \S_B_LOGIC_reg[22]  ( .G(n78), .D(B[22]), .Q(S_B_LOGIC[22]) );
  DLH_X1 \S_B_LOGIC_reg[21]  ( .G(n1535), .D(B[21]), .Q(S_B_LOGIC[21]) );
  DLH_X1 \S_B_LOGIC_reg[20]  ( .G(n78), .D(B[20]), .Q(S_B_LOGIC[20]) );
  DLH_X1 \S_B_LOGIC_reg[19]  ( .G(n78), .D(B[19]), .Q(S_B_LOGIC[19]) );
  DLH_X1 \S_B_LOGIC_reg[18]  ( .G(n78), .D(B[18]), .Q(S_B_LOGIC[18]) );
  DLH_X1 \S_B_LOGIC_reg[17]  ( .G(n78), .D(B[17]), .Q(S_B_LOGIC[17]) );
  DLH_X1 \S_B_LOGIC_reg[16]  ( .G(n78), .D(B[16]), .Q(S_B_LOGIC[16]) );
  DLH_X1 \S_B_LOGIC_reg[15]  ( .G(n78), .D(B[15]), .Q(S_B_LOGIC[15]) );
  DLH_X1 \S_B_LOGIC_reg[14]  ( .G(n78), .D(B[14]), .Q(S_B_LOGIC[14]) );
  DLH_X1 \S_B_LOGIC_reg[13]  ( .G(n1535), .D(B[13]), .Q(S_B_LOGIC[13]) );
  DLH_X1 \S_B_LOGIC_reg[12]  ( .G(n78), .D(B[12]), .Q(S_B_LOGIC[12]) );
  DLH_X1 \S_B_LOGIC_reg[11]  ( .G(n78), .D(B[11]), .Q(S_B_LOGIC[11]) );
  DLH_X1 \S_B_LOGIC_reg[10]  ( .G(n78), .D(B[10]), .Q(S_B_LOGIC[10]) );
  DLH_X1 \S_B_LOGIC_reg[9]  ( .G(n1535), .D(B[9]), .Q(S_B_LOGIC[9]) );
  DLH_X1 \S_B_LOGIC_reg[8]  ( .G(n78), .D(B[8]), .Q(S_B_LOGIC[8]) );
  DLH_X1 \S_B_LOGIC_reg[7]  ( .G(n1527), .D(B[7]), .Q(S_B_LOGIC[7]) );
  DLH_X1 \S_B_LOGIC_reg[6]  ( .G(n1535), .D(B[6]), .Q(S_B_LOGIC[6]) );
  DLH_X1 \S_B_LOGIC_reg[5]  ( .G(n78), .D(B[5]), .Q(S_B_LOGIC[5]) );
  DLH_X1 \S_B_LOGIC_reg[4]  ( .G(n78), .D(B[4]), .Q(S_B_LOGIC[4]) );
  DLH_X1 \S_B_LOGIC_reg[3]  ( .G(n1535), .D(B[3]), .Q(S_B_LOGIC[3]) );
  DLH_X1 \S_B_LOGIC_reg[2]  ( .G(n1535), .D(B[2]), .Q(S_B_LOGIC[2]) );
  DLH_X1 \S_B_LOGIC_reg[1]  ( .G(n1535), .D(B[1]), .Q(S_B_LOGIC[1]) );
  DLH_X1 \S_B_LOGIC_reg[0]  ( .G(n78), .D(B[0]), .Q(S_B_LOGIC[0]) );
  DLH_X1 \s_LOGIC_reg[3]  ( .G(n1527), .D(N89), .Q(s_LOGIC[3]) );
  DLH_X1 \s_LOGIC_reg[1]  ( .G(n1535), .D(n4843), .Q(s_LOGIC[1]) );
  DLH_X1 \s_A_SHIFT_reg[31]  ( .G(n6451), .D(A[31]), .Q(s_A_SHIFT[31]) );
  DLH_X1 \s_A_SHIFT_reg[30]  ( .G(n71), .D(A[30]), .Q(s_A_SHIFT[30]) );
  DLH_X1 \s_A_SHIFT_reg[29]  ( .G(n71), .D(A[29]), .Q(s_A_SHIFT[29]) );
  DLH_X1 \s_A_SHIFT_reg[28]  ( .G(n71), .D(A[28]), .Q(s_A_SHIFT[28]) );
  DLH_X1 \s_A_SHIFT_reg[27]  ( .G(n71), .D(A[27]), .Q(s_A_SHIFT[27]) );
  DLH_X1 \s_A_SHIFT_reg[26]  ( .G(n71), .D(A[26]), .Q(s_A_SHIFT[26]) );
  DLH_X1 \s_A_SHIFT_reg[25]  ( .G(n71), .D(A[25]), .Q(s_A_SHIFT[25]) );
  DLH_X1 \s_A_SHIFT_reg[24]  ( .G(n71), .D(A[24]), .Q(s_A_SHIFT[24]) );
  DLH_X1 \s_A_SHIFT_reg[23]  ( .G(n71), .D(A[23]), .Q(s_A_SHIFT[23]) );
  DLH_X1 \s_A_SHIFT_reg[22]  ( .G(n71), .D(A[22]), .Q(s_A_SHIFT[22]) );
  DLH_X1 \s_A_SHIFT_reg[21]  ( .G(n71), .D(A[21]), .Q(s_A_SHIFT[21]) );
  DLH_X1 \s_A_SHIFT_reg[20]  ( .G(n1404), .D(A[20]), .Q(s_A_SHIFT[20]) );
  DLH_X1 \s_A_SHIFT_reg[19]  ( .G(n71), .D(A[19]), .Q(s_A_SHIFT[19]) );
  DLH_X1 \s_A_SHIFT_reg[18]  ( .G(n1404), .D(A[18]), .Q(s_A_SHIFT[18]) );
  DLH_X1 \s_A_SHIFT_reg[17]  ( .G(n6451), .D(A[17]), .Q(s_A_SHIFT[17]) );
  DLH_X1 \s_A_SHIFT_reg[16]  ( .G(n71), .D(A[16]), .Q(s_A_SHIFT[16]) );
  DLH_X1 \s_A_SHIFT_reg[15]  ( .G(n71), .D(A[15]), .Q(s_A_SHIFT[15]) );
  DLH_X1 \s_A_SHIFT_reg[14]  ( .G(n1404), .D(A[14]), .Q(s_A_SHIFT[14]) );
  DLH_X1 \s_A_SHIFT_reg[13]  ( .G(n6451), .D(A[13]), .Q(s_A_SHIFT[13]) );
  DLH_X1 \s_A_SHIFT_reg[12]  ( .G(n71), .D(A[12]), .Q(s_A_SHIFT[12]) );
  DLH_X1 \s_A_SHIFT_reg[11]  ( .G(n71), .D(A[11]), .Q(s_A_SHIFT[11]) );
  DLH_X1 \s_A_SHIFT_reg[10]  ( .G(n1404), .D(A[10]), .Q(s_A_SHIFT[10]) );
  DLH_X1 \s_A_SHIFT_reg[9]  ( .G(n6451), .D(A[9]), .Q(s_A_SHIFT[9]) );
  DLH_X1 \s_A_SHIFT_reg[8]  ( .G(n71), .D(A[8]), .Q(s_A_SHIFT[8]) );
  DLH_X1 \s_A_SHIFT_reg[7]  ( .G(n71), .D(A[7]), .Q(s_A_SHIFT[7]) );
  DLH_X1 \s_A_SHIFT_reg[6]  ( .G(n1404), .D(A[6]), .Q(s_A_SHIFT[6]) );
  DLH_X1 \s_A_SHIFT_reg[5]  ( .G(n1404), .D(A[5]), .Q(s_A_SHIFT[5]) );
  DLH_X1 \s_A_SHIFT_reg[4]  ( .G(n1404), .D(A[4]), .Q(s_A_SHIFT[4]) );
  DLH_X1 \s_A_SHIFT_reg[3]  ( .G(n1404), .D(A[3]), .Q(s_A_SHIFT[3]) );
  DLH_X1 \s_A_SHIFT_reg[2]  ( .G(n6451), .D(A[2]), .Q(s_A_SHIFT[2]) );
  DLH_X1 \s_A_SHIFT_reg[1]  ( .G(n6451), .D(A[1]), .Q(s_A_SHIFT[1]) );
  DLH_X1 \s_A_SHIFT_reg[0]  ( .G(n71), .D(A[0]), .Q(s_A_SHIFT[0]) );
  DLH_X1 \S_B_SHIFT_reg[4]  ( .G(n6451), .D(B[4]), .Q(S_B_SHIFT[4]) );
  DLH_X1 \S_B_SHIFT_reg[3]  ( .G(n6451), .D(B[3]), .Q(S_B_SHIFT[3]) );
  DLH_X1 \S_B_SHIFT_reg[2]  ( .G(n71), .D(B[2]), .Q(S_B_SHIFT[2]) );
  DLH_X1 \S_B_SHIFT_reg[1]  ( .G(n6451), .D(B[1]), .Q(S_B_SHIFT[1]) );
  DLH_X1 \S_B_SHIFT_reg[0]  ( .G(n6451), .D(B[0]), .Q(S_B_SHIFT[0]) );
  DLH_X1 \s_SHIFT_reg[1]  ( .G(n71), .D(n1618), .Q(s_SHIFT[1]) );
  DLH_X1 \s_SHIFT_reg[0]  ( .G(n71), .D(n1619), .Q(s_SHIFT[0]) );
  DLH_X1 \s_A_MULT_reg[13]  ( .G(n72), .D(A[13]), .Q(s_A_MULT[13]) );
  DLH_X1 \s_A_MULT_reg[6]  ( .G(n72), .D(A[6]), .Q(s_A_MULT[6]) );
  DLH_X1 \s_A_MULT_reg[4]  ( .G(n72), .D(A[4]), .Q(s_A_MULT[4]) );
  DLH_X1 \s_A_MULT_reg[3]  ( .G(n72), .D(A[3]), .Q(s_A_MULT[3]) );
  DLH_X1 \s_A_MULT_reg[2]  ( .G(n72), .D(A[2]), .Q(s_A_MULT[2]) );
  DLH_X1 \S_B_MULT_reg[15]  ( .G(n72), .D(B[15]), .Q(S_B_MULT[15]) );
  DLH_X1 \S_B_MULT_reg[14]  ( .G(n72), .D(B[14]), .Q(S_B_MULT[14]) );
  DLH_X1 \S_B_MULT_reg[13]  ( .G(n1617), .D(B[13]), .Q(S_B_MULT[13]) );
  DLH_X1 \S_B_MULT_reg[12]  ( .G(n72), .D(B[12]), .Q(S_B_MULT[12]) );
  DLH_X1 \S_B_MULT_reg[10]  ( .G(n1617), .D(B[10]), .Q(S_B_MULT[10]) );
  DLH_X1 \S_B_MULT_reg[9]  ( .G(n1617), .D(B[9]), .Q(S_B_MULT[9]) );
  DLH_X1 \S_B_MULT_reg[8]  ( .G(n72), .D(B[8]), .Q(S_B_MULT[8]) );
  DLH_X1 \S_B_MULT_reg[7]  ( .G(n1617), .D(B[7]), .Q(S_B_MULT[7]) );
  DLH_X1 \S_B_MULT_reg[6]  ( .G(n72), .D(B[6]), .Q(S_B_MULT[6]) );
  DLH_X1 \S_B_MULT_reg[5]  ( .G(n1617), .D(B[5]), .Q(S_B_MULT[5]) );
  DLH_X1 \S_B_MULT_reg[4]  ( .G(n1617), .D(B[4]), .Q(S_B_MULT[4]) );
  DLH_X1 \S_B_MULT_reg[3]  ( .G(n1617), .D(B[3]), .Q(S_B_MULT[3]) );
  DLH_X1 \S_B_MULT_reg[2]  ( .G(n1617), .D(B[2]), .Q(S_B_MULT[2]) );
  DLH_X1 \S_B_MULT_reg[1]  ( .G(n1617), .D(B[1]), .Q(S_B_MULT[1]) );
  DLH_X1 \S_B_MULT_reg[0]  ( .G(n72), .D(B[0]), .Q(S_B_MULT[0]) );
  DLH_X1 \s_A_ADDER_reg[0]  ( .G(N21), .D(N22), .Q(s_A_ADDER[0]) );
  DLH_X1 \S_B_ADDER_reg[17]  ( .G(n80), .D(n6330), .Q(S_B_ADDER[17]) );
  DLH_X1 \s_A_ADDER_reg[16]  ( .G(N21), .D(n6331), .Q(s_A_ADDER[16]) );
  DLH_X1 \S_B_ADDER_reg[16]  ( .G(n80), .D(n6333), .Q(S_B_ADDER[16]) );
  DLH_X1 \s_A_ADDER_reg[15]  ( .G(N21), .D(n127), .Q(s_A_ADDER[15]) );
  DLH_X1 \S_B_ADDER_reg[15]  ( .G(n80), .D(n3332), .Q(S_B_ADDER[15]) );
  DLH_X1 \s_A_ADDER_reg[14]  ( .G(n80), .D(n3333), .Q(s_A_ADDER[14]) );
  DLH_X1 \S_B_ADDER_reg[14]  ( .G(n80), .D(n6334), .Q(S_B_ADDER[14]) );
  DLH_X1 \s_A_ADDER_reg[13]  ( .G(n80), .D(n3331), .Q(s_A_ADDER[13]) );
  DLH_X1 \s_A_ADDER_reg[12]  ( .G(N21), .D(N34), .Q(s_A_ADDER[12]) );
  DLH_X1 \S_B_ADDER_reg[13]  ( .G(n80), .D(N67), .Q(S_B_ADDER[13]) );
  DLH_X1 \S_B_ADDER_reg[12]  ( .G(N21), .D(N66), .Q(S_B_ADDER[12]) );
  DLH_X1 \s_A_ADDER_reg[11]  ( .G(n80), .D(N33), .Q(s_A_ADDER[11]) );
  DLH_X1 \S_B_ADDER_reg[11]  ( .G(N21), .D(n6337), .Q(S_B_ADDER[11]) );
  DLH_X1 \s_A_ADDER_reg[10]  ( .G(N21), .D(n6336), .Q(s_A_ADDER[10]) );
  DLH_X1 \S_B_ADDER_reg[10]  ( .G(N21), .D(n6339), .Q(S_B_ADDER[10]) );
  DLH_X1 \s_A_ADDER_reg[9]  ( .G(n80), .D(N31), .Q(s_A_ADDER[9]) );
  DLH_X1 \s_A_ADDER_reg[8]  ( .G(n80), .D(N30), .Q(s_A_ADDER[8]) );
  DLH_X1 \S_B_ADDER_reg[9]  ( .G(N21), .D(N63), .Q(S_B_ADDER[9]) );
  DLH_X1 \S_B_ADDER_reg[8]  ( .G(N21), .D(N62), .Q(S_B_ADDER[8]) );
  DLH_X1 \s_A_ADDER_reg[7]  ( .G(n80), .D(N29), .Q(s_A_ADDER[7]) );
  DLH_X1 \S_B_ADDER_reg[7]  ( .G(n80), .D(N61), .Q(S_B_ADDER[7]) );
  DLH_X1 \s_A_ADDER_reg[6]  ( .G(N21), .D(N28), .Q(s_A_ADDER[6]) );
  DLH_X1 \S_B_ADDER_reg[6]  ( .G(N21), .D(N60), .Q(S_B_ADDER[6]) );
  DLH_X1 \s_A_ADDER_reg[5]  ( .G(n80), .D(N27), .Q(s_A_ADDER[5]) );
  DLH_X1 \s_A_ADDER_reg[4]  ( .G(n80), .D(n4841), .Q(s_A_ADDER[4]) );
  DLH_X1 \s_A_ADDER_reg[3]  ( .G(N21), .D(N25), .Q(s_A_ADDER[3]) );
  DLH_X1 \s_A_ADDER_reg[2]  ( .G(n80), .D(n4842), .Q(s_A_ADDER[2]) );
  DLH_X1 \s_A_ADDER_reg[1]  ( .G(n80), .D(n6346), .Q(s_A_ADDER[1]) );
  DLH_X1 \s_A_ADDER_reg[31]  ( .G(N21), .D(N53), .Q(s_A_ADDER[31]) );
  DLH_X1 \S_B_ADDER_reg[31]  ( .G(n80), .D(n88), .Q(S_B_ADDER[31]) );
  DLH_X1 \s_A_ADDER_reg[30]  ( .G(n80), .D(n87), .Q(s_A_ADDER[30]) );
  DLH_X1 \S_B_ADDER_reg[30]  ( .G(n80), .D(n89), .Q(S_B_ADDER[30]) );
  DLH_X1 \s_A_ADDER_reg[29]  ( .G(N21), .D(n900), .Q(n1) );
  DLH_X1 \S_B_ADDER_reg[29]  ( .G(n80), .D(n6321), .Q(S_B_ADDER[29]) );
  DLH_X1 \s_A_ADDER_reg[28]  ( .G(n80), .D(n7620), .Q(s_A_ADDER[28]) );
  DLH_X1 \s_A_ADDER_reg[27]  ( .G(N21), .D(n93), .Q(s_A_ADDER[27]) );
  DLH_X1 \S_B_ADDER_reg[28]  ( .G(n80), .D(n6320), .Q(S_B_ADDER[28]) );
  DLH_X1 \s_A_ADDER_reg[26]  ( .G(n80), .D(n96), .Q(s_A_ADDER[26]) );
  DLH_X1 \S_B_ADDER_reg[27]  ( .G(N21), .D(n6322), .Q(S_B_ADDER[27]) );
  DLH_X1 \s_A_ADDER_reg[25]  ( .G(n80), .D(n4840), .Q(s_A_ADDER[25]) );
  DLH_X1 \S_B_ADDER_reg[26]  ( .G(N21), .D(n6323), .Q(S_B_ADDER[26]) );
  DLH_X1 \S_B_ADDER_reg[25]  ( .G(N21), .D(n6327), .Q(S_B_ADDER[25]) );
  DLH_X1 \s_A_ADDER_reg[24]  ( .G(N21), .D(n105), .Q(s_A_ADDER[24]) );
  DLH_X1 \S_B_ADDER_reg[24]  ( .G(N21), .D(n6324), .Q(S_B_ADDER[24]) );
  DLH_X1 \s_A_ADDER_reg[23]  ( .G(N21), .D(n107), .Q(s_A_ADDER[23]) );
  DLH_X1 \S_B_ADDER_reg[23]  ( .G(N21), .D(n6325), .Q(S_B_ADDER[23]) );
  DLH_X1 \s_A_ADDER_reg[22]  ( .G(n80), .D(n110), .Q(s_A_ADDER[22]) );
  DLH_X1 \S_B_ADDER_reg[18]  ( .G(N21), .D(n3309), .Q(S_B_ADDER[18]) );
  DLH_X1 \s_A_ADDER_reg[17]  ( .G(N21), .D(n122), .Q(s_A_ADDER[17]) );
  DLH_X1 \S_B_ADDER_reg[19]  ( .G(N21), .D(n3308), .Q(S_B_ADDER[19]) );
  DLH_X1 \s_A_ADDER_reg[18]  ( .G(n80), .D(n119), .Q(s_A_ADDER[18]) );
  DLH_X1 \S_B_ADDER_reg[22]  ( .G(N21), .D(n6326), .Q(S_B_ADDER[22]) );
  DLH_X1 \s_A_ADDER_reg[21]  ( .G(n80), .D(n3314), .Q(s_A_ADDER[21]) );
  DLH_X1 \S_B_ADDER_reg[21]  ( .G(N21), .D(n6329), .Q(S_B_ADDER[21]) );
  DLH_X1 \s_A_ADDER_reg[20]  ( .G(n80), .D(n1119), .Q(n24) );
  DLH_X1 \S_B_ADDER_reg[20]  ( .G(N21), .D(n118), .Q(S_B_ADDER[20]) );
  DLH_X1 \s_A_ADDER_reg[19]  ( .G(n80), .D(n1155), .Q(n26) );
  DLH_X1 \S_B_LHI_reg[15]  ( .G(n75), .D(B[15]), .Q(S_B_LHI[15]) );
  DLH_X1 \S_B_LHI_reg[14]  ( .G(n75), .D(B[14]), .Q(S_B_LHI[14]) );
  DLH_X1 \S_B_LHI_reg[13]  ( .G(n75), .D(B[13]), .Q(S_B_LHI[13]) );
  DLH_X1 \S_B_LHI_reg[12]  ( .G(n75), .D(B[12]), .Q(S_B_LHI[12]) );
  DLH_X1 \S_B_LHI_reg[11]  ( .G(n75), .D(B[11]), .Q(S_B_LHI[11]) );
  DLH_X1 \S_B_LHI_reg[10]  ( .G(n75), .D(B[10]), .Q(S_B_LHI[10]) );
  DLH_X1 \S_B_LHI_reg[9]  ( .G(n75), .D(B[9]), .Q(S_B_LHI[9]) );
  DLH_X1 \S_B_LHI_reg[8]  ( .G(n75), .D(B[8]), .Q(S_B_LHI[8]) );
  DLH_X1 \S_B_LHI_reg[7]  ( .G(n75), .D(B[7]), .Q(S_B_LHI[7]) );
  DLH_X1 \S_B_LHI_reg[6]  ( .G(n75), .D(B[6]), .Q(S_B_LHI[6]) );
  DLH_X1 \S_B_LHI_reg[5]  ( .G(n75), .D(B[5]), .Q(S_B_LHI[5]) );
  DLH_X1 \S_B_LHI_reg[4]  ( .G(n1616), .D(B[4]), .Q(S_B_LHI[4]) );
  DLH_X1 \S_B_LHI_reg[3]  ( .G(n75), .D(B[3]), .Q(S_B_LHI[3]) );
  DLH_X1 \S_B_LHI_reg[2]  ( .G(n1616), .D(B[2]), .Q(S_B_LHI[2]) );
  DLH_X1 \S_B_LHI_reg[1]  ( .G(n75), .D(B[1]), .Q(S_B_LHI[1]) );
  DLH_X1 \S_B_LHI_reg[0]  ( .G(n1616), .D(B[0]), .Q(S_B_LHI[0]) );
  FA_X1 \intadd_0/U9  ( .A(s_A_ADDER[24]), .B(\intadd_0/B[0] ), .CI(
        \intadd_0/CI ), .CO(\intadd_0/n8 ), .S(\intadd_0/SUM[0] ) );
  FA_X1 \intadd_0/U8  ( .A(s_A_ADDER[25]), .B(\intadd_0/B[1] ), .CI(
        \intadd_0/n8 ), .CO(\intadd_0/n7 ), .S(\intadd_0/SUM[1] ) );
  FA_X1 \intadd_0/U7  ( .A(s_A_ADDER[26]), .B(\intadd_0/B[2] ), .CI(
        \intadd_0/n7 ), .CO(\intadd_0/n6 ), .S(\intadd_0/SUM[2] ) );
  FA_X1 \intadd_0/U6  ( .A(s_A_ADDER[27]), .B(\intadd_0/B[3] ), .CI(
        \intadd_0/n6 ), .CO(\intadd_0/n5 ), .S(\intadd_0/SUM[3] ) );
  FA_X1 \intadd_0/U5  ( .A(s_A_ADDER[28]), .B(\intadd_0/B[4] ), .CI(
        \intadd_0/n5 ), .CO(\intadd_0/n4 ), .S(\intadd_0/SUM[4] ) );
  FA_X1 \intadd_0/U4  ( .A(n6433), .B(\intadd_0/B[5] ), .CI(\intadd_0/n4 ), 
        .CO(\intadd_0/n3 ), .S(\intadd_0/SUM[5] ) );
  FA_X1 \intadd_0/U3  ( .A(s_A_ADDER[30]), .B(\intadd_0/B[6] ), .CI(
        \intadd_0/n3 ), .CO(\intadd_0/n2 ), .S(\intadd_0/SUM[6] ) );
  FA_X1 \intadd_0/U2  ( .A(s_A_ADDER[31]), .B(\intadd_0/B[7] ), .CI(
        \intadd_0/n2 ), .CO(\intadd_0/n1 ), .S(\intadd_0/SUM[7] ) );
  FA_X1 \intadd_1/U9  ( .A(n6432), .B(\intadd_1/B[0] ), .CI(\intadd_1/CI ), 
        .CO(\intadd_1/n8 ), .S(\intadd_1/SUM[0] ) );
  FA_X1 \intadd_1/U8  ( .A(n6431), .B(\intadd_1/B[1] ), .CI(\intadd_1/n8 ), 
        .CO(\intadd_1/n7 ), .S(\intadd_1/SUM[1] ) );
  FA_X1 \intadd_1/U7  ( .A(n6430), .B(\intadd_1/B[2] ), .CI(\intadd_1/n7 ), 
        .CO(\intadd_1/n6 ), .S(\intadd_1/SUM[2] ) );
  FA_X1 \intadd_1/U6  ( .A(n6429), .B(\intadd_1/B[3] ), .CI(\intadd_1/n6 ), 
        .CO(\intadd_1/n5 ), .S(\intadd_1/SUM[3] ) );
  FA_X1 \intadd_1/U5  ( .A(n6428), .B(\intadd_1/B[4] ), .CI(\intadd_1/n5 ), 
        .CO(\intadd_1/n4 ), .S(\intadd_1/SUM[4] ) );
  FA_X1 \intadd_1/U4  ( .A(n6427), .B(\intadd_1/B[5] ), .CI(\intadd_1/n4 ), 
        .CO(\intadd_1/n3 ), .S(\intadd_1/SUM[5] ) );
  FA_X1 \intadd_1/U3  ( .A(n6426), .B(\intadd_1/B[6] ), .CI(\intadd_1/n3 ), 
        .CO(\intadd_1/n2 ), .S(\intadd_1/SUM[6] ) );
  FA_X1 \intadd_1/U2  ( .A(n6425), .B(\intadd_1/B[7] ), .CI(\intadd_1/n2 ), 
        .CO(\intadd_1/n1 ), .S(\intadd_1/SUM[7] ) );
  FA_X1 \intadd_2/U5  ( .A(\intadd_2/A[0] ), .B(\intadd_2/B[0] ), .CI(
        \intadd_2/CI ), .CO(\intadd_2/n4 ), .S(\intadd_2/SUM[0] ) );
  FA_X1 \intadd_2/U4  ( .A(\intadd_2/A[1] ), .B(\intadd_2/B[1] ), .CI(
        \intadd_2/n4 ), .CO(\intadd_2/n3 ), .S(\intadd_2/SUM[1] ) );
  FA_X1 \intadd_2/U3  ( .A(\intadd_2/A[2] ), .B(\intadd_2/B[2] ), .CI(
        \intadd_2/n3 ), .CO(\intadd_2/n2 ), .S(\intadd_2/SUM[2] ) );
  FA_X1 \intadd_2/U2  ( .A(\intadd_2/A[3] ), .B(\intadd_2/B[3] ), .CI(
        \intadd_2/n2 ), .CO(\intadd_2/n1 ), .S(\intadd_2/SUM[3] ) );
  FA_X1 \intadd_3/U5  ( .A(\intadd_3/A[0] ), .B(\intadd_3/B[0] ), .CI(
        \intadd_3/CI ), .CO(\intadd_3/n4 ), .S(\intadd_3/SUM[0] ) );
  FA_X1 \intadd_3/U4  ( .A(\intadd_3/A[1] ), .B(\intadd_3/B[1] ), .CI(
        \intadd_3/n4 ), .CO(\intadd_3/n3 ), .S(\intadd_3/SUM[1] ) );
  FA_X1 \intadd_3/U3  ( .A(\intadd_3/A[2] ), .B(\intadd_3/B[2] ), .CI(
        \intadd_3/n3 ), .CO(\intadd_3/n2 ), .S(\intadd_3/SUM[2] ) );
  FA_X1 \intadd_3/U2  ( .A(\intadd_3/A[3] ), .B(\intadd_3/B[3] ), .CI(
        \intadd_3/n2 ), .CO(\intadd_3/n1 ), .S(\intadd_3/SUM[3] ) );
  FA_X1 \intadd_4/U5  ( .A(\intadd_4/A[0] ), .B(\intadd_4/B[0] ), .CI(
        \intadd_4/CI ), .CO(\intadd_4/n4 ), .S(\intadd_3/A[1] ) );
  FA_X1 \intadd_4/U4  ( .A(\intadd_4/A[1] ), .B(\intadd_4/B[1] ), .CI(
        \intadd_4/n4 ), .CO(\intadd_4/n3 ), .S(\intadd_3/B[2] ) );
  FA_X1 \intadd_4/U3  ( .A(\intadd_4/A[2] ), .B(\intadd_4/B[2] ), .CI(
        \intadd_4/n3 ), .CO(\intadd_4/n2 ), .S(\intadd_3/A[3] ) );
  FA_X1 \intadd_4/U2  ( .A(\intadd_4/A[3] ), .B(\intadd_4/B[3] ), .CI(
        \intadd_4/n2 ), .CO(\intadd_4/n1 ), .S(\intadd_4/SUM[3] ) );
  FA_X1 \intadd_5/U4  ( .A(\intadd_5/A[0] ), .B(\intadd_5/B[0] ), .CI(
        \intadd_5/CI ), .CO(\intadd_5/n3 ), .S(\intadd_5/SUM[0] ) );
  FA_X1 \intadd_5/U3  ( .A(\intadd_3/SUM[0] ), .B(\intadd_5/B[1] ), .CI(
        \intadd_5/n3 ), .CO(\intadd_5/n2 ), .S(\intadd_5/SUM[1] ) );
  FA_X1 \intadd_5/U2  ( .A(\intadd_5/A[2] ), .B(\intadd_3/SUM[1] ), .CI(
        \intadd_5/n2 ), .CO(\intadd_5/n1 ), .S(\intadd_5/SUM[2] ) );
  FA_X1 \intadd_6/U4  ( .A(\intadd_6/A[0] ), .B(\intadd_6/B[0] ), .CI(
        \intadd_6/CI ), .CO(\intadd_6/n3 ), .S(\intadd_2/B[1] ) );
  FA_X1 \intadd_6/U3  ( .A(\intadd_6/A[1] ), .B(\intadd_5/SUM[0] ), .CI(
        \intadd_6/n3 ), .CO(\intadd_6/n2 ), .S(\intadd_2/B[2] ) );
  FA_X1 \intadd_6/U2  ( .A(\intadd_6/A[2] ), .B(\intadd_5/SUM[1] ), .CI(
        \intadd_6/n2 ), .CO(\intadd_6/n1 ), .S(\intadd_2/A[3] ) );
  FA_X1 \intadd_7/U4  ( .A(\intadd_7/A[0] ), .B(\intadd_7/B[0] ), .CI(
        \intadd_7/CI ), .CO(\intadd_7/n3 ), .S(\intadd_4/B[1] ) );
  FA_X1 \intadd_7/U3  ( .A(\intadd_7/A[1] ), .B(\intadd_7/B[1] ), .CI(
        \intadd_7/n3 ), .CO(\intadd_7/n2 ), .S(\intadd_4/B[2] ) );
  FA_X1 \intadd_7/U2  ( .A(\intadd_7/A[2] ), .B(\intadd_7/B[2] ), .CI(
        \intadd_7/n2 ), .CO(\intadd_7/n1 ), .S(\intadd_4/A[3] ) );
  FA_X1 \intadd_8/U4  ( .A(\intadd_8/A[0] ), .B(\intadd_8/B[0] ), .CI(
        \intadd_8/CI ), .CO(\intadd_8/n3 ), .S(\intadd_7/B[1] ) );
  FA_X1 \intadd_8/U3  ( .A(\intadd_8/A[1] ), .B(\intadd_8/B[1] ), .CI(
        \intadd_8/n3 ), .CO(\intadd_8/n2 ), .S(\intadd_7/B[2] ) );
  FA_X1 \intadd_8/U2  ( .A(\intadd_8/A[2] ), .B(\intadd_8/B[2] ), .CI(
        \intadd_8/n2 ), .CO(\intadd_8/n1 ), .S(\intadd_8/SUM[2] ) );
  FA_X1 \intadd_9/U4  ( .A(\intadd_8/B[0] ), .B(\intadd_9/B[0] ), .CI(
        \intadd_9/CI ), .CO(\intadd_9/n3 ), .S(\intadd_8/A[1] ) );
  FA_X1 \intadd_9/U3  ( .A(\intadd_9/A[1] ), .B(\intadd_9/B[1] ), .CI(
        \intadd_9/n3 ), .CO(\intadd_9/n2 ), .S(\intadd_8/A[2] ) );
  FA_X1 \intadd_9/U2  ( .A(n7619), .B(\intadd_9/B[2] ), .CI(\intadd_9/n2 ), 
        .CO(\intadd_9/n1 ), .S(\intadd_9/SUM[2] ) );
  FA_X1 \intadd_10/U4  ( .A(\intadd_10/A[0] ), .B(\intadd_10/B[0] ), .CI(
        \intadd_10/CI ), .CO(\intadd_10/n3 ), .S(\intadd_10/SUM[0] ) );
  FA_X1 \intadd_10/U3  ( .A(\intadd_2/SUM[0] ), .B(\intadd_10/B[1] ), .CI(
        \intadd_10/n3 ), .CO(\intadd_10/n2 ), .S(\intadd_10/SUM[1] ) );
  FA_X1 \intadd_10/U2  ( .A(\intadd_10/A[2] ), .B(\intadd_2/SUM[1] ), .CI(
        \intadd_10/n2 ), .CO(\intadd_10/n1 ), .S(\intadd_10/SUM[2] ) );
  FA_X1 \intadd_11/U4  ( .A(\intadd_11/A[0] ), .B(\intadd_11/B[0] ), .CI(
        \intadd_11/CI ), .CO(\intadd_11/n3 ), .S(\intadd_11/SUM[0] ) );
  FA_X1 \intadd_11/U3  ( .A(\intadd_11/A[1] ), .B(\intadd_11/B[1] ), .CI(
        \intadd_11/n3 ), .CO(\intadd_11/n2 ), .S(\intadd_11/SUM[1] ) );
  FA_X1 \intadd_11/U2  ( .A(\intadd_11/A[2] ), .B(\intadd_11/B[2] ), .CI(
        \intadd_11/n2 ), .CO(\intadd_11/n1 ), .S(\intadd_11/SUM[2] ) );
  FA_X1 \intadd_12/U4  ( .A(\intadd_12/A[0] ), .B(\intadd_12/B[0] ), .CI(
        \intadd_12/CI ), .CO(\intadd_12/n3 ), .S(\intadd_12/SUM[0] ) );
  FA_X1 \intadd_12/U3  ( .A(\intadd_12/A[1] ), .B(\intadd_11/SUM[0] ), .CI(
        \intadd_12/n3 ), .CO(\intadd_12/n2 ), .S(\intadd_12/SUM[1] ) );
  FA_X1 \intadd_12/U2  ( .A(\intadd_12/A[2] ), .B(\intadd_11/SUM[1] ), .CI(
        \intadd_12/n2 ), .CO(\intadd_12/n1 ), .S(\intadd_12/SUM[2] ) );
  DLH_X1 \s_A_MULT_reg[5]  ( .G(n72), .D(A[5]), .Q(s_A_MULT[5]) );
  DLH_X1 \s_A_MULT_reg[8]  ( .G(n72), .D(A[8]), .Q(s_A_MULT[8]) );
  DLH_X1 \s_A_MULT_reg[15]  ( .G(n1617), .D(A[15]), .Q(s_A_MULT[15]) );
  DLH_X1 \s_A_MULT_reg[11]  ( .G(n72), .D(A[11]), .Q(s_A_MULT[11]) );
  DLH_X1 \s_A_MULT_reg[14]  ( .G(n72), .D(A[14]), .Q(s_A_MULT[14]) );
  DLH_X1 \s_A_MULT_reg[7]  ( .G(n1617), .D(A[7]), .Q(s_A_MULT[7]) );
  DLH_X1 \S_B_MULT_reg[11]  ( .G(n72), .D(B[11]), .Q(S_B_MULT[11]) );
  DLH_X1 \s_A_MULT_reg[12]  ( .G(n1617), .D(A[12]), .Q(s_A_MULT[12]) );
  DLH_X1 \s_A_MULT_reg[9]  ( .G(n72), .D(A[9]), .Q(s_A_MULT[9]) );
  DLH_X1 \s_A_MULT_reg[10]  ( .G(n72), .D(A[10]), .Q(s_A_MULT[10]) );
  DLH_X1 \s_A_MULT_reg[1]  ( .G(n72), .D(A[1]), .Q(s_A_MULT[1]) );
  DLH_X1 \s_A_MULT_reg[0]  ( .G(n1617), .D(A[0]), .Q(\MULT/SHIFTERi_0/N19 ) );
  AOI22_X1 U3449 ( .A1(n643), .A2(s_A_SHIFT[23]), .B1(n644), .B2(s_A_SHIFT[15]), .ZN(n2) );
  OAI211_X1 U3450 ( .C1(n57), .C2(n646), .A(n645), .B(n2), .ZN(n3) );
  AOI22_X1 U3451 ( .A1(n1433), .A2(n3), .B1(n648), .B2(n647), .ZN(n4) );
  AOI22_X1 U3453 ( .A1(n649), .A2(\intadd_0/SUM[7] ), .B1(n1616), .B2(
        S_B_LHI[15]), .ZN(n6) );
  NAND2_X1 U3454 ( .A1(s_A_LOGIC[31]), .A2(S_B_LOGIC[31]), .ZN(n7) );
  OAI221_X1 U3456 ( .B1(n7), .B2(n1403), .C1(s_A_LOGIC[31]), .C2(S_B_LOGIC[31]), .A(n8), .ZN(n9) );
  NAND4_X1 U3457 ( .A1(n4), .A2(n5), .A3(n6), .A4(n9), .ZN(Y[31]) );
  INV_X1 U3458 ( .A(S_B_LOGIC[19]), .ZN(n10) );
  OAI22_X1 U3462 ( .A1(n1406), .A2(n463), .B1(n1421), .B2(n464), .ZN(n14) );
  OAI22_X1 U3463 ( .A1(n726), .A2(n532), .B1(n1423), .B2(n502), .ZN(n15) );
  OAI221_X1 U3465 ( .B1(S_B_LOGIC[19]), .B2(n1428), .C1(n10), .C2(n1403), .A(
        s_A_LOGIC[19]), .ZN(n17) );
  INV_X1 U3467 ( .A(S_B_LOGIC[17]), .ZN(n18) );
  AOI22_X1 U3469 ( .A1(n75), .A2(S_B_LHI[1]), .B1(n649), .B2(n446), .ZN(n20)
         );
  OAI21_X1 U3470 ( .B1(n695), .B2(n454), .A(n20), .ZN(n21) );
  OAI22_X1 U3471 ( .A1(n730), .A2(n532), .B1(n614), .B2(n444), .ZN(n22) );
  OAI22_X1 U3472 ( .A1(n726), .A2(n502), .B1(n678), .B2(n464), .ZN(n23) );
  NOR4_X1 U3473 ( .A1(n19), .A2(n21), .A3(n22), .A4(n23), .ZN(n25) );
  OAI221_X1 U3474 ( .B1(S_B_LOGIC[17]), .B2(n1399), .C1(n18), .C2(n1403), .A(
        s_A_LOGIC[17]), .ZN(n27) );
  OAI211_X1 U3475 ( .C1(n728), .C2(n460), .A(n25), .B(n27), .ZN(Y[17]) );
  NAND2_X1 U3476 ( .A1(n329), .A2(n331), .ZN(n28) );
  AOI22_X1 U3477 ( .A1(n1441), .A2(n329), .B1(n1400), .B2(n28), .ZN(n29) );
  INV_X1 U3478 ( .A(n311), .ZN(n30) );
  OAI221_X1 U3479 ( .B1(n478), .B2(n688), .C1(n478), .C2(n663), .A(n6451), 
        .ZN(n31) );
  AOI211_X1 U3480 ( .C1(n475), .C2(n663), .A(n323), .B(n322), .ZN(n32) );
  AOI21_X1 U3481 ( .B1(n711), .B2(n31), .A(n32), .ZN(n33) );
  OAI21_X1 U3482 ( .B1(S_B_LOGIC[0]), .B2(s_A_LOGIC[0]), .A(n324), .ZN(n34) );
  OAI22_X1 U3483 ( .A1(n1420), .A2(n324), .B1(n1435), .B2(n34), .ZN(n35) );
  XNOR2_X1 U3485 ( .A(n329), .B(n1401), .ZN(n37) );
  NOR2_X1 U3486 ( .A1(n325), .A2(n326), .ZN(n38) );
  AOI21_X1 U3487 ( .B1(n329), .B2(n331), .A(n327), .ZN(n39) );
  AOI21_X1 U3488 ( .B1(n331), .B2(n38), .A(n39), .ZN(n40) );
  OAI22_X1 U3489 ( .A1(n1157), .A2(n37), .B1(n1452), .B2(n40), .ZN(n41) );
  NOR2_X1 U3490 ( .A1(n1441), .A2(n1454), .ZN(n42) );
  AOI222_X1 U3491 ( .A1(n28), .A2(n1454), .B1(n331), .B2(n42), .C1(n1441), 
        .C2(n329), .ZN(n43) );
  AOI22_X1 U3492 ( .A1(n1430), .A2(n41), .B1(n332), .B2(n43), .ZN(n44) );
  OAI211_X1 U3493 ( .C1(n333), .C2(n29), .A(n36), .B(n44), .ZN(Y[0]) );
  AOI22_X1 U3496 ( .A1(n1433), .A2(n717), .B1(n718), .B2(n721), .ZN(n47) );
  NAND2_X1 U3497 ( .A1(s_A_LOGIC[8]), .A2(S_B_LOGIC[8]), .ZN(n48) );
  OAI22_X1 U3498 ( .A1(s_A_LOGIC[8]), .A2(S_B_LOGIC[8]), .B1(n737), .B2(n48), 
        .ZN(n49) );
  OAI22_X1 U3500 ( .A1(n714), .A2(n715), .B1(n713), .B2(n725), .ZN(n51) );
  AOI211_X1 U3501 ( .C1(n719), .C2(n1418), .A(n50), .B(n51), .ZN(n52) );
  OAI211_X1 U3502 ( .C1(n1406), .C2(\intadd_1/SUM[6] ), .A(n47), .B(n52), .ZN(
        Y[8]) );
  OR4_X1 U3503 ( .A1(S_B_MULT[7]), .A2(S_B_MULT[8]), .A3(n204), .A4(n176), 
        .ZN(n53) );
  OR3_X1 U3504 ( .A1(n204), .A2(S_B_MULT[0]), .A3(n942), .ZN(n54) );
  AOI211_X2 U3505 ( .C1(n66), .C2(s_A_SHIFT[27]), .A(n484), .B(n483), .ZN(n569) );
  INV_X1 U3506 ( .A(n54), .ZN(n55) );
  AOI211_X2 U3507 ( .C1(s_A_SHIFT[2]), .C2(n643), .A(n431), .B(n346), .ZN(n444) );
  AOI211_X2 U3508 ( .C1(s_A_SHIFT[8]), .C2(n643), .A(n431), .B(n430), .ZN(n532) );
  AOI211_X2 U3509 ( .C1(s_A_SHIFT[4]), .C2(n643), .A(n431), .B(n380), .ZN(n464) );
  INV_X1 U3510 ( .A(n53), .ZN(n56) );
  NOR3_X2 U3511 ( .A1(n174), .A2(n176), .A3(n204), .ZN(n1069) );
  NOR3_X2 U3512 ( .A1(n204), .A2(n203), .A3(n205), .ZN(n1258) );
  NOR2_X2 U3513 ( .A1(n317), .A2(n315), .ZN(n702) );
  NOR2_X2 U3514 ( .A1(n318), .A2(n317), .ZN(n663) );
  NOR2_X2 U3515 ( .A1(n204), .A2(n1001), .ZN(n1159) );
  NOR2_X2 U3516 ( .A1(S_B_MULT[11]), .A2(n179), .ZN(n1085) );
  NOR2_X2 U3517 ( .A1(S_B_MULT[9]), .A2(n174), .ZN(n1070) );
  NOR2_X2 U3518 ( .A1(S_B_MULT[5]), .A2(n113), .ZN(n968) );
  NOR2_X2 U3519 ( .A1(n204), .A2(n972), .ZN(n967) );
  NOR2_X2 U3520 ( .A1(n850), .A2(s_A_MULT[15]), .ZN(n204) );
  NOR2_X2 U3521 ( .A1(n314), .A2(n440), .ZN(n616) );
  NOR2_X2 U3522 ( .A1(S_B_MULT[7]), .A2(n150), .ZN(n1076) );
  NOR2_X2 U3523 ( .A1(S_B_MULT[7]), .A2(n133), .ZN(n1048) );
  NOR2_X2 U3524 ( .A1(S_B_MULT[5]), .A2(n106), .ZN(n966) );
  AOI211_X2 U3525 ( .C1(n66), .C2(s_A_SHIFT[25]), .A(n484), .B(n448), .ZN(n557) );
  AOI211_X2 U3526 ( .C1(s_A_SHIFT[6]), .C2(n643), .A(n431), .B(n404), .ZN(n502) );
  AOI221_X4 U3527 ( .B1(n325), .B2(n1401), .C1(n1432), .C2(n1157), .A(n1430), 
        .ZN(n649) );
  NOR2_X2 U3528 ( .A1(S_B_MULT[13]), .A2(n206), .ZN(n1259) );
  NOR2_X2 U3530 ( .A1(S_B_MULT[11]), .A2(n200), .ZN(n1160) );
  NOR2_X2 U3531 ( .A1(S_B_MULT[15]), .A2(n214), .ZN(n1246) );
  NOR2_X2 U3532 ( .A1(S_B_MULT[9]), .A2(n175), .ZN(n1073) );
  NOR2_X2 U3533 ( .A1(n427), .A2(n440), .ZN(n644) );
  NOR4_X4 U3534 ( .A1(S_B_MULT[6]), .A2(n204), .A3(S_B_MULT[5]), .A4(n1043), 
        .ZN(n1075) );
  BUF_X1 U3536 ( .A(N21), .Z(n80) );
  NAND2_X1 U3537 ( .A1(n1156), .A2(n1405), .ZN(N21) );
  BUF_X1 U3539 ( .A(n1527), .Z(n78) );
  INV_X1 U3540 ( .A(n197), .ZN(n221) );
  INV_X1 U3541 ( .A(n72), .ZN(n73) );
  INV_X1 U3542 ( .A(n72), .ZN(n74) );
  INV_X1 U3543 ( .A(s_A_MULT[15]), .ZN(n1164) );
  INV_X1 U3544 ( .A(n838), .ZN(n1307) );
  INV_X1 U3545 ( .A(n1231), .ZN(n1260) );
  NOR2_X1 U3546 ( .A1(n1515), .A2(n83), .ZN(n1617) );
  INV_X1 U3547 ( .A(n855), .ZN(n1309) );
  INV_X1 U3548 ( .A(n856), .ZN(n1308) );
  INV_X1 U3549 ( .A(n204), .ZN(n816) );
  INV_X1 U3550 ( .A(s_A_MULT[13]), .ZN(n1236) );
  INV_X1 U3551 ( .A(s_A_MULT[14]), .ZN(n1079) );
  BUF_X1 U3552 ( .A(n1396), .Z(n70) );
  INV_X1 U3553 ( .A(n1374), .ZN(n1396) );
  INV_X1 U3554 ( .A(N91), .ZN(n1156) );
  OR2_X1 U3557 ( .A1(n1454), .A2(n424), .ZN(n333) );
  INV_X1 U3559 ( .A(n77), .ZN(n76) );
  INV_X1 U3560 ( .A(\ADD_SUB/carry_ST[0] ), .ZN(n77) );
  INV_X1 U3567 ( .A(n736), .ZN(n695) );
  INV_X1 U3569 ( .A(OP[4]), .ZN(n1154) );
  INV_X1 U3571 ( .A(OP[1]), .ZN(n328) );
  INV_X1 U3573 ( .A(n698), .ZN(n686) );
  INV_X1 U3574 ( .A(n704), .ZN(n687) );
  INV_X1 U3575 ( .A(n57), .ZN(n67) );
  INV_X1 U3576 ( .A(n59), .ZN(n66) );
  OR3_X1 U3577 ( .A1(S_B_SHIFT[4]), .A2(S_B_SHIFT[3]), .A3(n314), .ZN(n59) );
  NOR2_X2 U3578 ( .A1(S_B_MULT[3]), .A2(n91), .ZN(n948) );
  NOR2_X2 U3579 ( .A1(S_B_MULT[15]), .A2(n213), .ZN(n1247) );
  NOR2_X2 U3580 ( .A1(S_B_MULT[13]), .A2(n205), .ZN(n1262) );
  NAND2_X1 U3581 ( .A1(n81), .A2(n1452), .ZN(n83) );
  NOR2_X2 U3582 ( .A1(n427), .A2(n441), .ZN(n643) );
  NOR2_X2 U3583 ( .A1(n314), .A2(n441), .ZN(n617) );
  NOR2_X1 U3584 ( .A1(n1247), .A2(n1246), .ZN(n60) );
  NOR2_X1 U3585 ( .A1(n1262), .A2(n1259), .ZN(n62) );
  NOR2_X1 U3586 ( .A1(n1085), .A2(n1160), .ZN(n64) );
  OR3_X1 U3587 ( .A1(S_B_SHIFT[4]), .A2(S_B_SHIFT[3]), .A3(n427), .ZN(n57) );
  INV_X1 U3588 ( .A(n1258), .ZN(n63) );
  INV_X1 U3589 ( .A(n1159), .ZN(n65) );
  INV_X1 U3590 ( .A(n1239), .ZN(n61) );
  BUF_X1 U3591 ( .A(n1617), .Z(n72) );
  MUX2_X1 U3592 ( .A(n60), .B(n61), .S(n1164), .Z(n222) );
  MUX2_X1 U3593 ( .A(n62), .B(n63), .S(n1164), .Z(n1216) );
  MUX2_X1 U3594 ( .A(n64), .B(n65), .S(n1164), .Z(n1251) );
  INV_X1 U3595 ( .A(n58), .ZN(n68) );
  OAI221_X1 U3597 ( .B1(n1454), .B2(n1441), .C1(n1454), .C2(n1432), .A(n1430), 
        .ZN(n82) );
  NAND2_X1 U3599 ( .A1(n1154), .A2(OP[0]), .ZN(n1136) );
  INV_X1 U3600 ( .A(n1451), .ZN(n81) );
  INV_X1 U3601 ( .A(n83), .ZN(n332) );
  NAND2_X1 U3602 ( .A1(n332), .A2(n1515), .ZN(n245) );
  OAI211_X1 U3603 ( .C1(n1452), .C2(n82), .A(n333), .B(n245), .ZN(N91) );
  INV_X1 U3606 ( .A(A[0]), .ZN(n85) );
  NOR3_X1 U3607 ( .A1(s_A_MULT[1]), .A2(\MULT/SHIFTERi_0/N19 ), .A3(
        s_A_MULT[2]), .ZN(n97) );
  INV_X1 U3608 ( .A(s_A_MULT[3]), .ZN(n137) );
  NAND2_X1 U3609 ( .A1(n97), .A2(n137), .ZN(n104) );
  NOR2_X1 U3610 ( .A1(s_A_MULT[4]), .A2(n104), .ZN(n120) );
  INV_X1 U3611 ( .A(s_A_MULT[5]), .ZN(n787) );
  NAND2_X1 U3612 ( .A1(n120), .A2(n787), .ZN(n140) );
  NOR2_X1 U3613 ( .A1(s_A_MULT[6]), .A2(n140), .ZN(n169) );
  INV_X1 U3614 ( .A(s_A_MULT[7]), .ZN(n766) );
  NAND2_X1 U3615 ( .A1(n169), .A2(n766), .ZN(n173) );
  NOR2_X1 U3616 ( .A1(s_A_MULT[8]), .A2(n173), .ZN(n172) );
  INV_X1 U3617 ( .A(s_A_MULT[9]), .ZN(n915) );
  NAND2_X1 U3618 ( .A1(n172), .A2(n915), .ZN(n779) );
  NOR2_X1 U3619 ( .A1(s_A_MULT[10]), .A2(n779), .ZN(n824) );
  INV_X1 U3620 ( .A(s_A_MULT[11]), .ZN(n840) );
  NAND2_X1 U3621 ( .A1(n824), .A2(n840), .ZN(n841) );
  NOR2_X1 U3622 ( .A1(s_A_MULT[12]), .A2(n841), .ZN(n853) );
  NAND2_X1 U3623 ( .A1(n853), .A2(n1236), .ZN(n852) );
  INV_X1 U3624 ( .A(n852), .ZN(n851) );
  NAND2_X1 U3625 ( .A1(n1079), .A2(n851), .ZN(n850) );
  NAND3_X1 U3626 ( .A1(S_B_MULT[1]), .A2(S_B_MULT[0]), .A3(n816), .ZN(n856) );
  INV_X1 U3627 ( .A(S_B_MULT[1]), .ZN(n942) );
  NAND2_X1 U3628 ( .A1(S_B_MULT[0]), .A2(n942), .ZN(n855) );
  OAI211_X1 U3629 ( .C1(n1308), .C2(n1309), .A(\MULT/SHIFTERi_0/N19 ), .B(n72), 
        .ZN(n84) );
  OAI21_X1 U3630 ( .B1(n70), .B2(n85), .A(n84), .ZN(N22) );
  INV_X1 U3631 ( .A(A[3]), .ZN(n101) );
  INV_X1 U3632 ( .A(s_A_MULT[1]), .ZN(n910) );
  INV_X1 U3633 ( .A(\MULT/SHIFTERi_0/N19 ), .ZN(n797) );
  NAND2_X1 U3634 ( .A1(n910), .A2(n797), .ZN(n86) );
  AOI21_X1 U3635 ( .B1(s_A_MULT[2]), .B2(n86), .A(n97), .ZN(n908) );
  OAI21_X1 U3636 ( .B1(n797), .B2(n910), .A(n86), .ZN(n838) );
  AOI222_X1 U3637 ( .A1(s_A_MULT[2]), .A2(n1309), .B1(n1308), .B2(n908), .C1(
        n1307), .C2(n55), .ZN(n1194) );
  INV_X1 U3638 ( .A(S_B_MULT[2]), .ZN(n90) );
  AOI22_X1 U3639 ( .A1(S_B_MULT[1]), .A2(n90), .B1(S_B_MULT[2]), .B2(n942), 
        .ZN(n91) );
  INV_X1 U3640 ( .A(S_B_MULT[3]), .ZN(n92) );
  NOR2_X1 U3641 ( .A1(n92), .A2(n91), .ZN(n939) );
  NAND2_X1 U3642 ( .A1(n939), .A2(n816), .ZN(n941) );
  INV_X1 U3643 ( .A(n941), .ZN(n94) );
  OAI21_X1 U3644 ( .B1(n948), .B2(n94), .A(\MULT/SHIFTERi_0/N19 ), .ZN(n1193)
         );
  NOR2_X1 U3645 ( .A1(n1194), .A2(n1193), .ZN(n1192) );
  NAND3_X1 U3646 ( .A1(S_B_MULT[2]), .A2(S_B_MULT[1]), .A3(n92), .ZN(n945) );
  NOR2_X1 U3647 ( .A1(S_B_MULT[2]), .A2(n92), .ZN(n943) );
  NAND3_X1 U3648 ( .A1(n943), .A2(n816), .A3(n942), .ZN(n936) );
  NAND2_X1 U3649 ( .A1(n945), .A2(n936), .ZN(n95) );
  AOI222_X1 U3650 ( .A1(n95), .A2(\MULT/SHIFTERi_0/N19 ), .B1(n94), .B2(n1307), 
        .C1(s_A_MULT[1]), .C2(n948), .ZN(n124) );
  OAI21_X1 U3651 ( .B1(n97), .B2(n137), .A(n104), .ZN(n934) );
  INV_X1 U3652 ( .A(n934), .ZN(n899) );
  AOI222_X1 U3653 ( .A1(n899), .A2(n1308), .B1(n1309), .B2(s_A_MULT[3]), .C1(
        n908), .C2(n55), .ZN(n98) );
  INV_X1 U3654 ( .A(n98), .ZN(n125) );
  XNOR2_X1 U3655 ( .A(n124), .B(n125), .ZN(n99) );
  NAND2_X1 U3656 ( .A1(n1192), .A2(n99), .ZN(n1186) );
  OAI211_X1 U3657 ( .C1(n1192), .C2(n99), .A(n72), .B(n1186), .ZN(n100) );
  OAI21_X1 U3658 ( .B1(n70), .B2(n101), .A(n100), .ZN(N25) );
  INV_X1 U3659 ( .A(A[5]), .ZN(n129) );
  NOR2_X1 U3660 ( .A1(n910), .A2(n945), .ZN(n103) );
  INV_X1 U3661 ( .A(n908), .ZN(n902) );
  OAI22_X1 U3662 ( .A1(n941), .A2(n902), .B1(n838), .B2(n936), .ZN(n102) );
  AOI211_X1 U3663 ( .C1(n948), .C2(s_A_MULT[2]), .A(n103), .B(n102), .ZN(n112)
         );
  AOI21_X1 U3664 ( .B1(s_A_MULT[4]), .B2(n104), .A(n120), .ZN(n959) );
  AOI222_X1 U3665 ( .A1(s_A_MULT[4]), .A2(n1309), .B1(n1308), .B2(n959), .C1(
        n899), .C2(n55), .ZN(n111) );
  NOR2_X1 U3666 ( .A1(S_B_MULT[3]), .A2(S_B_MULT[4]), .ZN(n969) );
  AOI21_X1 U3667 ( .B1(S_B_MULT[4]), .B2(S_B_MULT[3]), .A(n969), .ZN(n108) );
  INV_X1 U3668 ( .A(n108), .ZN(n106) );
  NAND2_X1 U3669 ( .A1(S_B_MULT[5]), .A2(n108), .ZN(n972) );
  OAI21_X1 U3670 ( .B1(n966), .B2(n967), .A(\MULT/SHIFTERi_0/N19 ), .ZN(n109)
         );
  NOR2_X1 U3671 ( .A1(n1189), .A2(n1186), .ZN(n231) );
  FA_X1 U3672 ( .A(n112), .B(n111), .CI(n109), .CO(n123), .S(n1189) );
  NAND2_X1 U3673 ( .A1(S_B_MULT[3]), .A2(S_B_MULT[4]), .ZN(n113) );
  INV_X1 U3674 ( .A(n968), .ZN(n973) );
  NAND3_X1 U3675 ( .A1(S_B_MULT[5]), .A2(n969), .A3(n816), .ZN(n1056) );
  NAND2_X1 U3676 ( .A1(n973), .A2(n1056), .ZN(n114) );
  AOI222_X1 U3677 ( .A1(n114), .A2(\MULT/SHIFTERi_0/N19 ), .B1(n967), .B2(
        n1307), .C1(s_A_MULT[1]), .C2(n966), .ZN(n132) );
  INV_X1 U3678 ( .A(s_A_MULT[2]), .ZN(n115) );
  NOR2_X1 U3679 ( .A1(n115), .A2(n945), .ZN(n117) );
  OAI22_X1 U3680 ( .A1(n941), .A2(n934), .B1(n902), .B2(n936), .ZN(n116) );
  AOI211_X1 U3681 ( .C1(n948), .C2(s_A_MULT[3]), .A(n117), .B(n116), .ZN(n131)
         );
  OAI21_X1 U3682 ( .B1(n120), .B2(n787), .A(n140), .ZN(n988) );
  INV_X1 U3683 ( .A(n988), .ZN(n831) );
  AOI222_X1 U3684 ( .A1(s_A_MULT[5]), .A2(n1309), .B1(n1308), .B2(n831), .C1(
        n959), .C2(n55), .ZN(n130) );
  NOR2_X1 U3685 ( .A1(n121), .A2(n123), .ZN(n141) );
  AOI21_X1 U3686 ( .B1(n123), .B2(n121), .A(n141), .ZN(n1385) );
  INV_X1 U3687 ( .A(n124), .ZN(n126) );
  NAND2_X1 U3688 ( .A1(n126), .A2(n125), .ZN(n1187) );
  NOR2_X1 U3689 ( .A1(n1189), .A2(n1187), .ZN(n1384) );
  XOR2_X1 U3690 ( .A(n1385), .B(n1384), .Z(n230) );
  XNOR2_X1 U3691 ( .A(n231), .B(n230), .ZN(n128) );
  OAI22_X1 U3692 ( .A1(n70), .A2(n129), .B1(n73), .B2(n128), .ZN(N27) );
  INV_X1 U3693 ( .A(A[6]), .ZN(n146) );
  FA_X1 U3694 ( .A(n132), .B(n131), .CI(n130), .CO(n149), .S(n121) );
  NAND2_X1 U3695 ( .A1(S_B_MULT[6]), .A2(S_B_MULT[5]), .ZN(n150) );
  OAI21_X1 U3696 ( .B1(S_B_MULT[6]), .B2(S_B_MULT[5]), .A(n150), .ZN(n133) );
  INV_X1 U3697 ( .A(S_B_MULT[7]), .ZN(n1043) );
  NOR2_X1 U3698 ( .A1(n1043), .A2(n133), .ZN(n1081) );
  NAND2_X1 U3699 ( .A1(n1081), .A2(n816), .ZN(n1046) );
  INV_X1 U3700 ( .A(n1046), .ZN(n134) );
  OAI21_X1 U3701 ( .B1(n1048), .B2(n134), .A(\MULT/SHIFTERi_0/N19 ), .ZN(n148)
         );
  AOI22_X1 U3702 ( .A1(s_A_MULT[2]), .A2(n966), .B1(n967), .B2(n908), .ZN(n135) );
  OAI21_X1 U3703 ( .B1(n838), .B2(n1056), .A(n135), .ZN(n136) );
  AOI21_X1 U3704 ( .B1(s_A_MULT[1]), .B2(n968), .A(n136), .ZN(n154) );
  NOR2_X1 U3705 ( .A1(n137), .A2(n945), .ZN(n139) );
  INV_X1 U3706 ( .A(n959), .ZN(n833) );
  OAI22_X1 U3707 ( .A1(n941), .A2(n833), .B1(n934), .B2(n936), .ZN(n138) );
  AOI211_X1 U3708 ( .C1(n948), .C2(s_A_MULT[4]), .A(n139), .B(n138), .ZN(n153)
         );
  AOI21_X1 U3709 ( .B1(s_A_MULT[6]), .B2(n140), .A(n169), .ZN(n1089) );
  AOI222_X1 U3710 ( .A1(s_A_MULT[6]), .A2(n1309), .B1(n1308), .B2(n1089), .C1(
        n831), .C2(n55), .ZN(n152) );
  INV_X1 U3711 ( .A(n141), .ZN(n142) );
  NOR2_X1 U3712 ( .A1(n143), .A2(n142), .ZN(n235) );
  AOI21_X1 U3713 ( .B1(n143), .B2(n142), .A(n235), .ZN(n1383) );
  NAND2_X1 U3714 ( .A1(n1385), .A2(n1384), .ZN(n144) );
  XOR2_X1 U3715 ( .A(n1383), .B(n144), .Z(n145) );
  OAI22_X1 U3716 ( .A1(n70), .A2(n146), .B1(n73), .B2(n145), .ZN(N28) );
  INV_X1 U3717 ( .A(A[7]), .ZN(n158) );
  FA_X1 U3718 ( .A(n149), .B(n148), .CI(n147), .CO(n156), .S(n143) );
  INV_X1 U3719 ( .A(n1048), .ZN(n1078) );
  OAI22_X1 U3720 ( .A1(n910), .A2(n1078), .B1(n1046), .B2(n838), .ZN(n151) );
  AOI221_X1 U3721 ( .B1(n1076), .B2(\MULT/SHIFTERi_0/N19 ), .C1(n1075), .C2(
        \MULT/SHIFTERi_0/N19 ), .A(n151), .ZN(n160) );
  FA_X1 U3722 ( .A(n154), .B(n153), .CI(n152), .CO(n159), .S(n147) );
  NOR2_X1 U3723 ( .A1(n155), .A2(n156), .ZN(n1389) );
  AOI21_X1 U3724 ( .B1(n156), .B2(n155), .A(n1389), .ZN(n234) );
  XNOR2_X1 U3725 ( .A(n235), .B(n234), .ZN(n157) );
  OAI22_X1 U3726 ( .A1(n70), .A2(n158), .B1(n73), .B2(n157), .ZN(N29) );
  INV_X1 U3727 ( .A(A[8]), .ZN(n163) );
  FA_X1 U3728 ( .A(\intadd_12/SUM[0] ), .B(n160), .CI(n159), .CO(n161), .S(
        n155) );
  NOR2_X1 U3729 ( .A1(n161), .A2(\intadd_12/SUM[1] ), .ZN(n1313) );
  AOI21_X1 U3730 ( .B1(\intadd_12/SUM[1] ), .B2(n161), .A(n1313), .ZN(n1388)
         );
  XNOR2_X1 U3731 ( .A(n1389), .B(n1388), .ZN(n162) );
  OAI22_X1 U3732 ( .A1(n70), .A2(n163), .B1(n73), .B2(n162), .ZN(N30) );
  INV_X1 U3733 ( .A(A[9]), .ZN(n165) );
  XOR2_X1 U3734 ( .A(n1313), .B(\intadd_12/SUM[2] ), .Z(n164) );
  OAI22_X1 U3735 ( .A1(n70), .A2(n165), .B1(n73), .B2(n164), .ZN(N31) );
  INV_X1 U3736 ( .A(A[11]), .ZN(n189) );
  INV_X1 U3737 ( .A(\intadd_10/SUM[1] ), .ZN(n192) );
  AOI22_X1 U3738 ( .A1(s_A_MULT[4]), .A2(n968), .B1(n967), .B2(n831), .ZN(n166) );
  OAI21_X1 U3739 ( .B1(n833), .B2(n1056), .A(n166), .ZN(n167) );
  AOI21_X1 U3740 ( .B1(s_A_MULT[5]), .B2(n966), .A(n167), .ZN(n792) );
  INV_X1 U3741 ( .A(s_A_MULT[6]), .ZN(n168) );
  NOR2_X1 U3742 ( .A1(n168), .A2(n945), .ZN(n171) );
  OAI21_X1 U3743 ( .B1(n169), .B2(n766), .A(n173), .ZN(n1087) );
  INV_X1 U3744 ( .A(n1089), .ZN(n922) );
  OAI22_X1 U3745 ( .A1(n941), .A2(n1087), .B1(n922), .B2(n936), .ZN(n170) );
  AOI211_X1 U3746 ( .C1(n948), .C2(s_A_MULT[7]), .A(n171), .B(n170), .ZN(n791)
         );
  OAI21_X1 U3747 ( .B1(n172), .B2(n915), .A(n779), .ZN(n1083) );
  INV_X1 U3748 ( .A(n1083), .ZN(n979) );
  AOI21_X1 U3749 ( .B1(s_A_MULT[8]), .B2(n173), .A(n172), .ZN(n1068) );
  AOI222_X1 U3750 ( .A1(s_A_MULT[9]), .A2(n1309), .B1(n1308), .B2(n979), .C1(
        n55), .C2(n1068), .ZN(n790) );
  NAND2_X1 U3751 ( .A1(S_B_MULT[8]), .A2(S_B_MULT[7]), .ZN(n175) );
  OAI21_X1 U3752 ( .B1(S_B_MULT[8]), .B2(S_B_MULT[7]), .A(n175), .ZN(n174) );
  INV_X1 U3753 ( .A(S_B_MULT[9]), .ZN(n176) );
  AOI22_X1 U3754 ( .A1(n1070), .A2(s_A_MULT[2]), .B1(n1069), .B2(n908), .ZN(
        n178) );
  AOI22_X1 U3755 ( .A1(n1073), .A2(s_A_MULT[1]), .B1(n1307), .B2(n56), .ZN(
        n177) );
  NAND2_X1 U3756 ( .A1(n178), .A2(n177), .ZN(n187) );
  NOR2_X1 U3757 ( .A1(S_B_MULT[9]), .A2(S_B_MULT[10]), .ZN(n1161) );
  AOI21_X1 U3758 ( .B1(S_B_MULT[10]), .B2(S_B_MULT[9]), .A(n1161), .ZN(n180)
         );
  INV_X1 U3759 ( .A(n180), .ZN(n179) );
  INV_X1 U3760 ( .A(n1085), .ZN(n1165) );
  NAND2_X1 U3761 ( .A1(S_B_MULT[11]), .A2(n180), .ZN(n1001) );
  AOI21_X1 U3762 ( .B1(n1165), .B2(n65), .A(n797), .ZN(n186) );
  AOI22_X1 U3763 ( .A1(s_A_MULT[4]), .A2(n1048), .B1(s_A_MULT[3]), .B2(n1076), 
        .ZN(n182) );
  NAND2_X1 U3764 ( .A1(n899), .A2(n1075), .ZN(n181) );
  OAI211_X1 U3765 ( .C1(n833), .C2(n1046), .A(n182), .B(n181), .ZN(n185) );
  INV_X1 U3766 ( .A(n183), .ZN(n785) );
  INV_X1 U3767 ( .A(n184), .ZN(n191) );
  FA_X1 U3768 ( .A(n187), .B(n186), .CI(n185), .CO(n190), .S(n183) );
  XOR2_X1 U3769 ( .A(\intadd_11/n1 ), .B(n1393), .Z(n188) );
  OAI22_X1 U3770 ( .A1(n70), .A2(n189), .B1(n73), .B2(n188), .ZN(N33) );
  INV_X1 U3771 ( .A(A[12]), .ZN(n194) );
  FA_X1 U3772 ( .A(n192), .B(n191), .CI(n190), .CO(n239), .S(n1393) );
  XOR2_X1 U3773 ( .A(\intadd_10/SUM[2] ), .B(n239), .Z(n193) );
  OAI22_X1 U3774 ( .A1(n70), .A2(n194), .B1(n73), .B2(n193), .ZN(N34) );
  NAND2_X1 U3775 ( .A1(n1164), .A2(n816), .ZN(n197) );
  AOI22_X1 U3776 ( .A1(s_A_MULT[15]), .A2(n855), .B1(n856), .B2(n1164), .ZN(
        n940) );
  AOI21_X1 U3777 ( .B1(n221), .B2(S_B_MULT[1]), .A(n940), .ZN(\intadd_8/B[0] )
         );
  INV_X1 U3778 ( .A(A[31]), .ZN(n243) );
  NOR2_X1 U3779 ( .A1(n197), .A2(S_B_MULT[8]), .ZN(n196) );
  INV_X1 U3780 ( .A(n1069), .ZN(n1041) );
  OAI21_X1 U3781 ( .B1(n1070), .B2(n1073), .A(s_A_MULT[15]), .ZN(n195) );
  OAI21_X1 U3782 ( .B1(s_A_MULT[15]), .B2(n1041), .A(n195), .ZN(n1005) );
  AOI21_X1 U3783 ( .B1(n196), .B2(S_B_MULT[9]), .A(n1005), .ZN(n202) );
  NOR2_X1 U3784 ( .A1(n197), .A2(S_B_MULT[6]), .ZN(n199) );
  OAI21_X1 U3785 ( .B1(n1076), .B2(n1048), .A(s_A_MULT[15]), .ZN(n198) );
  OAI21_X1 U3786 ( .B1(s_A_MULT[15]), .B2(n1046), .A(n198), .ZN(n1014) );
  AOI21_X1 U3787 ( .B1(n199), .B2(S_B_MULT[7]), .A(n1014), .ZN(n1170) );
  NOR2_X1 U3788 ( .A1(n202), .A2(n1170), .ZN(n1255) );
  NAND2_X1 U3789 ( .A1(n221), .A2(S_B_MULT[11]), .ZN(n201) );
  NAND2_X1 U3790 ( .A1(S_B_MULT[9]), .A2(S_B_MULT[10]), .ZN(n200) );
  OAI21_X1 U3791 ( .B1(S_B_MULT[10]), .B2(n201), .A(n1251), .ZN(n217) );
  NAND2_X1 U3792 ( .A1(n202), .A2(n1170), .ZN(n1254) );
  OAI21_X1 U3793 ( .B1(n1255), .B2(n217), .A(n1254), .ZN(n1220) );
  NAND2_X1 U3794 ( .A1(n221), .A2(S_B_MULT[13]), .ZN(n207) );
  INV_X1 U3795 ( .A(S_B_MULT[13]), .ZN(n203) );
  NAND2_X1 U3796 ( .A1(S_B_MULT[11]), .A2(S_B_MULT[12]), .ZN(n206) );
  OAI21_X1 U3797 ( .B1(S_B_MULT[11]), .B2(S_B_MULT[12]), .A(n206), .ZN(n205)
         );
  OAI21_X1 U3798 ( .B1(S_B_MULT[12]), .B2(n207), .A(n1216), .ZN(n208) );
  INV_X1 U3799 ( .A(n208), .ZN(n209) );
  NAND2_X1 U3800 ( .A1(n1220), .A2(n209), .ZN(n1205) );
  INV_X1 U3801 ( .A(n1205), .ZN(n210) );
  NOR2_X1 U3802 ( .A1(n209), .A2(n1220), .ZN(n1203) );
  NOR2_X1 U3803 ( .A1(n210), .A2(n1203), .ZN(n1201) );
  NAND2_X1 U3804 ( .A1(n850), .A2(s_A_MULT[15]), .ZN(n1257) );
  INV_X1 U3805 ( .A(n1257), .ZN(n1253) );
  NOR2_X1 U3806 ( .A1(S_B_MULT[13]), .A2(S_B_MULT[14]), .ZN(n211) );
  NAND3_X1 U3807 ( .A1(S_B_MULT[15]), .A2(n211), .A3(n816), .ZN(n1242) );
  NAND2_X1 U3808 ( .A1(S_B_MULT[15]), .A2(n816), .ZN(n212) );
  NAND2_X1 U3809 ( .A1(S_B_MULT[13]), .A2(S_B_MULT[14]), .ZN(n214) );
  OAI21_X1 U3810 ( .B1(S_B_MULT[13]), .B2(S_B_MULT[14]), .A(n214), .ZN(n213)
         );
  NOR2_X1 U3811 ( .A1(n212), .A2(n213), .ZN(n1239) );
  OAI21_X1 U3812 ( .B1(n1253), .B2(n1242), .A(n222), .ZN(n215) );
  INV_X1 U3813 ( .A(n215), .ZN(n224) );
  XOR2_X1 U3814 ( .A(n1201), .B(n224), .Z(n1198) );
  INV_X1 U3815 ( .A(n1254), .ZN(n216) );
  NOR2_X1 U3816 ( .A1(n216), .A2(n1255), .ZN(n1266) );
  XNOR2_X1 U3817 ( .A(n1266), .B(n217), .ZN(n1268) );
  NAND2_X1 U3818 ( .A1(S_B_MULT[5]), .A2(n221), .ZN(n218) );
  OAI21_X1 U3819 ( .B1(n218), .B2(S_B_MULT[4]), .A(n1055), .ZN(n1054) );
  NOR2_X1 U3820 ( .A1(n948), .A2(n1164), .ZN(n219) );
  AOI22_X1 U3821 ( .A1(n219), .A2(n945), .B1(n1164), .B2(n941), .ZN(n993) );
  AOI21_X1 U3822 ( .B1(n221), .B2(n943), .A(n993), .ZN(n220) );
  NAND2_X1 U3823 ( .A1(\intadd_8/B[0] ), .A2(n220), .ZN(n1103) );
  NOR2_X1 U3824 ( .A1(n1054), .A2(n1103), .ZN(n1269) );
  NAND2_X1 U3825 ( .A1(n1268), .A2(n1269), .ZN(n1223) );
  NOR2_X1 U3826 ( .A1(\intadd_8/B[0] ), .A2(n220), .ZN(n1101) );
  NAND2_X1 U3827 ( .A1(n1101), .A2(n1054), .ZN(n1267) );
  NOR2_X1 U3828 ( .A1(n1268), .A2(n1267), .ZN(n1221) );
  AOI21_X1 U3829 ( .B1(n1198), .B2(n1223), .A(n1221), .ZN(n228) );
  NAND2_X1 U3830 ( .A1(S_B_MULT[15]), .A2(n221), .ZN(n223) );
  OAI21_X1 U3831 ( .B1(n223), .B2(S_B_MULT[14]), .A(n222), .ZN(n226) );
  OAI21_X1 U3832 ( .B1(n1203), .B2(n224), .A(n1205), .ZN(n225) );
  XOR2_X1 U3833 ( .A(n226), .B(n225), .Z(n227) );
  XNOR2_X1 U3834 ( .A(n228), .B(n227), .ZN(n229) );
  OAI22_X1 U3835 ( .A1(n1396), .A2(n243), .B1(n73), .B2(n229), .ZN(N53) );
  AND2_X1 U3836 ( .A1(n1416), .A2(B[0]), .ZN(N54) );
  AND2_X1 U3837 ( .A1(n1416), .A2(B[1]), .ZN(N55) );
  AND2_X1 U3838 ( .A1(n1416), .A2(B[2]), .ZN(N56) );
  AND2_X1 U3839 ( .A1(n1416), .A2(B[3]), .ZN(N57) );
  AND2_X1 U3840 ( .A1(n1416), .A2(B[4]), .ZN(N58) );
  AND2_X1 U3841 ( .A1(n1416), .A2(B[5]), .ZN(N59) );
  INV_X1 U3842 ( .A(B[6]), .ZN(n233) );
  NAND3_X1 U3843 ( .A1(n72), .A2(n231), .A3(n230), .ZN(n232) );
  OAI21_X1 U3844 ( .B1(n70), .B2(n233), .A(n232), .ZN(N60) );
  INV_X1 U3845 ( .A(B[8]), .ZN(n237) );
  NAND2_X1 U3846 ( .A1(n235), .A2(n234), .ZN(n236) );
  OAI22_X1 U3847 ( .A1(n1396), .A2(n237), .B1(n73), .B2(n236), .ZN(N62) );
  INV_X1 U3848 ( .A(B[13]), .ZN(n241) );
  INV_X1 U3849 ( .A(\intadd_10/SUM[2] ), .ZN(n238) );
  NAND2_X1 U3850 ( .A1(n239), .A2(n238), .ZN(n240) );
  OAI22_X1 U3851 ( .A1(n1396), .A2(n241), .B1(n73), .B2(n240), .ZN(N67) );
  NOR2_X1 U3852 ( .A1(OP[4]), .A2(OP[3]), .ZN(n246) );
  INV_X1 U3854 ( .A(n242), .ZN(n4843) );
  OAI22_X1 U3855 ( .A1(n1401), .A2(n242), .B1(n1526), .B2(n1451), .ZN(N89) );
  NAND2_X1 U3856 ( .A1(OP[2]), .A2(OP[1]), .ZN(n1135) );
  INV_X1 U3857 ( .A(n1135), .ZN(n247) );
  INV_X1 U3858 ( .A(B[31]), .ZN(n1212) );
  AOI22_X1 U3859 ( .A1(A[31]), .A2(n1212), .B1(B[31]), .B2(n243), .ZN(n244) );
  AOI221_X1 U3860 ( .B1(n247), .B2(n333), .C1(n245), .C2(n333), .A(n244), .ZN(
        N92) );
  XOR2_X1 U3863 ( .A(n76), .B(S_B_ADDER[20]), .Z(n749) );
  XNOR2_X1 U3864 ( .A(n749), .B(n24), .ZN(n259) );
  XOR2_X1 U3865 ( .A(n76), .B(S_B_ADDER[17]), .Z(n248) );
  NAND2_X1 U3866 ( .A1(n248), .A2(s_A_ADDER[17]), .ZN(n281) );
  INV_X1 U3867 ( .A(n281), .ZN(n249) );
  NOR2_X1 U3868 ( .A1(n248), .A2(s_A_ADDER[17]), .ZN(n280) );
  NOR2_X1 U3869 ( .A1(n249), .A2(n280), .ZN(n268) );
  XOR2_X1 U3870 ( .A(n76), .B(S_B_ADDER[16]), .Z(n254) );
  NAND2_X1 U3871 ( .A1(n254), .A2(s_A_ADDER[16]), .ZN(n265) );
  INV_X1 U3872 ( .A(n265), .ZN(n255) );
  XOR2_X1 U3873 ( .A(n76), .B(S_B_ADDER[18]), .Z(n307) );
  AOI22_X1 U3874 ( .A1(n268), .A2(n255), .B1(s_A_ADDER[18]), .B2(n307), .ZN(
        n250) );
  NOR2_X1 U3875 ( .A1(s_A_ADDER[18]), .A2(n307), .ZN(n257) );
  AOI21_X1 U3876 ( .B1(n250), .B2(n281), .A(n257), .ZN(n253) );
  XNOR2_X1 U3877 ( .A(n76), .B(S_B_ADDER[19]), .ZN(n256) );
  NAND2_X1 U3878 ( .A1(n26), .A2(n256), .ZN(n252) );
  NOR2_X1 U3879 ( .A1(n26), .A2(n256), .ZN(n251) );
  AOI21_X1 U3880 ( .B1(n253), .B2(n252), .A(n251), .ZN(n746) );
  NOR2_X1 U3881 ( .A1(n254), .A2(s_A_ADDER[16]), .ZN(n267) );
  NOR2_X1 U3882 ( .A1(n255), .A2(n267), .ZN(n260) );
  INV_X1 U3883 ( .A(s_A_ADDER[15]), .ZN(n285) );
  XNOR2_X1 U3884 ( .A(\ADD_SUB/carry_ST[0] ), .B(S_B_ADDER[15]), .ZN(n284) );
  INV_X1 U3885 ( .A(s_A_ADDER[14]), .ZN(n275) );
  XNOR2_X1 U3886 ( .A(n76), .B(S_B_ADDER[14]), .ZN(n274) );
  INV_X1 U3887 ( .A(s_A_ADDER[13]), .ZN(n278) );
  XNOR2_X1 U3888 ( .A(n76), .B(S_B_ADDER[13]), .ZN(n277) );
  INV_X1 U3889 ( .A(s_A_ADDER[12]), .ZN(n295) );
  XNOR2_X1 U3890 ( .A(n76), .B(S_B_ADDER[12]), .ZN(n294) );
  INV_X1 U3891 ( .A(s_A_ADDER[11]), .ZN(n298) );
  XNOR2_X1 U3892 ( .A(\ADD_SUB/carry_ST[0] ), .B(S_B_ADDER[11]), .ZN(n297) );
  INV_X1 U3893 ( .A(s_A_ADDER[10]), .ZN(n300) );
  XNOR2_X1 U3894 ( .A(\ADD_SUB/carry_ST[0] ), .B(S_B_ADDER[10]), .ZN(n299) );
  XNOR2_X1 U3895 ( .A(n26), .B(n256), .ZN(n309) );
  NOR3_X1 U3896 ( .A1(n257), .A2(n266), .A3(n309), .ZN(n258) );
  NAND3_X1 U3897 ( .A1(n268), .A2(n260), .A3(n258), .ZN(n745) );
  NAND2_X1 U3898 ( .A1(n746), .A2(n745), .ZN(n270) );
  XNOR2_X1 U3899 ( .A(n259), .B(n270), .ZN(n489) );
  XOR2_X1 U3900 ( .A(n260), .B(n266), .Z(n434) );
  XOR2_X1 U3901 ( .A(n76), .B(S_B_ADDER[1]), .Z(n765) );
  INV_X1 U3902 ( .A(n765), .ZN(n262) );
  NAND2_X1 U3903 ( .A1(s_A_ADDER[0]), .A2(n262), .ZN(n261) );
  OAI211_X1 U3904 ( .C1(s_A_ADDER[0]), .C2(n262), .A(S_B_ADDER[0]), .B(n261), 
        .ZN(n263) );
  OAI21_X1 U3905 ( .B1(S_B_ADDER[1]), .B2(S_B_ADDER[0]), .A(n263), .ZN(n264)
         );
  XNOR2_X1 U3906 ( .A(n264), .B(s_A_ADDER[1]), .ZN(n469) );
  OAI21_X1 U3907 ( .B1(n267), .B2(n266), .A(n265), .ZN(n279) );
  XOR2_X1 U3908 ( .A(n268), .B(n279), .Z(n446) );
  NOR4_X1 U3909 ( .A1(\intadd_0/SUM[5] ), .A2(\intadd_0/SUM[4] ), .A3(
        \intadd_0/SUM[3] ), .A4(\intadd_0/SUM[2] ), .ZN(n290) );
  NAND2_X1 U3910 ( .A1(\intadd_1/SUM[0] ), .A2(\intadd_1/SUM[1] ), .ZN(n269)
         );
  NOR3_X1 U3911 ( .A1(\intadd_0/SUM[6] ), .A2(\intadd_0/SUM[7] ), .A3(n269), 
        .ZN(n289) );
  INV_X1 U3912 ( .A(s_A_ADDER[22]), .ZN(n744) );
  XOR2_X1 U3913 ( .A(n76), .B(S_B_ADDER[22]), .Z(n757) );
  INV_X1 U3914 ( .A(n757), .ZN(n743) );
  INV_X1 U3915 ( .A(s_A_ADDER[21]), .ZN(n753) );
  XNOR2_X1 U3916 ( .A(\ADD_SUB/carry_ST[0] ), .B(S_B_ADDER[21]), .ZN(n754) );
  INV_X1 U3917 ( .A(n24), .ZN(n748) );
  INV_X1 U3918 ( .A(n749), .ZN(n747) );
  NAND2_X1 U3919 ( .A1(n24), .A2(n747), .ZN(n271) );
  AOI22_X1 U3920 ( .A1(n749), .A2(n748), .B1(n271), .B2(n270), .ZN(n272) );
  FA_X1 U3921 ( .A(n753), .B(n754), .CI(n272), .CO(n291), .S(n498) );
  FA_X1 U3922 ( .A(n275), .B(n274), .CI(n273), .CO(n283), .S(n410) );
  FA_X1 U3923 ( .A(n278), .B(n277), .CI(n276), .CO(n273), .S(n399) );
  AND4_X1 U3924 ( .A1(n514), .A2(n498), .A3(n410), .A4(n399), .ZN(n288) );
  INV_X1 U3925 ( .A(n279), .ZN(n282) );
  AOI21_X1 U3926 ( .B1(n282), .B2(n281), .A(n280), .ZN(n306) );
  FA_X1 U3927 ( .A(n285), .B(n284), .CI(n283), .CO(n266), .S(n286) );
  INV_X1 U3928 ( .A(n286), .ZN(n420) );
  NOR4_X1 U3929 ( .A1(\intadd_0/SUM[1] ), .A2(\intadd_0/SUM[0] ), .A3(n450), 
        .A4(n420), .ZN(n287) );
  NAND4_X1 U3930 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(n305) );
  FA_X1 U3931 ( .A(n744), .B(n743), .CI(n291), .CO(n292), .S(n514) );
  XOR2_X1 U3932 ( .A(n76), .B(S_B_ADDER[23]), .Z(n758) );
  XNOR2_X1 U3933 ( .A(n758), .B(s_A_ADDER[23]), .ZN(n761) );
  XNOR2_X1 U3934 ( .A(n292), .B(n761), .ZN(n531) );
  FA_X1 U3935 ( .A(n295), .B(n294), .CI(n293), .CO(n276), .S(n387) );
  FA_X1 U3936 ( .A(n298), .B(n297), .CI(n296), .CO(n293), .S(n376) );
  NAND4_X1 U3937 ( .A1(\intadd_1/SUM[5] ), .A2(\intadd_1/SUM[4] ), .A3(
        \intadd_1/SUM[3] ), .A4(\intadd_1/SUM[2] ), .ZN(n302) );
  INV_X1 U3938 ( .A(S_B_ADDER[0]), .ZN(n763) );
  NOR2_X1 U3939 ( .A1(s_A_ADDER[0]), .A2(n763), .ZN(n762) );
  AOI21_X1 U3940 ( .B1(s_A_ADDER[0]), .B2(n763), .A(n762), .ZN(n311) );
  FA_X1 U3941 ( .A(n300), .B(\intadd_1/n1 ), .CI(n299), .CO(n296), .S(n357) );
  NAND4_X1 U3942 ( .A1(n311), .A2(\intadd_1/SUM[7] ), .A3(\intadd_1/SUM[6] ), 
        .A4(n357), .ZN(n301) );
  NOR2_X1 U3943 ( .A1(n302), .A2(n301), .ZN(n303) );
  NAND4_X1 U3944 ( .A1(n531), .A2(n387), .A3(n376), .A4(n303), .ZN(n304) );
  NOR4_X1 U3945 ( .A1(n469), .A2(n446), .A3(n305), .A4(n304), .ZN(n310) );
  FA_X1 U3946 ( .A(s_A_ADDER[18]), .B(n307), .CI(n306), .CO(n308), .S(n450) );
  XOR2_X1 U3947 ( .A(n309), .B(n308), .Z(n463) );
  NAND4_X1 U3948 ( .A1(n489), .A2(n434), .A3(n310), .A4(n463), .ZN(n331) );
  XOR2_X1 U3949 ( .A(\intadd_0/n1 ), .B(s_SIGN), .Z(n329) );
  INV_X1 U3950 ( .A(s_SHIFT[0]), .ZN(n344) );
  INV_X1 U3951 ( .A(s_SHIFT[1]), .ZN(n312) );
  NAND2_X1 U3952 ( .A1(n344), .A2(n312), .ZN(n427) );
  XOR2_X1 U3953 ( .A(n427), .B(S_B_SHIFT[0]), .Z(n334) );
  XOR2_X1 U3955 ( .A(n427), .B(S_B_SHIFT[1]), .Z(n317) );
  XNOR2_X1 U3956 ( .A(n427), .B(S_B_SHIFT[2]), .ZN(n315) );
  INV_X1 U3957 ( .A(n702), .ZN(n677) );
  OAI21_X1 U3958 ( .B1(n312), .B2(n344), .A(n427), .ZN(n314) );
  INV_X1 U3959 ( .A(S_B_SHIFT[3]), .ZN(n313) );
  OR2_X1 U3960 ( .A1(n313), .A2(S_B_SHIFT[4]), .ZN(n441) );
  NAND2_X1 U3961 ( .A1(S_B_SHIFT[4]), .A2(n313), .ZN(n440) );
  AOI222_X1 U3962 ( .A1(n66), .A2(s_A_SHIFT[3]), .B1(n617), .B2(s_A_SHIFT[11]), 
        .C1(n616), .C2(s_A_SHIFT[19]), .ZN(n620) );
  NAND2_X1 U3963 ( .A1(n315), .A2(n317), .ZN(n698) );
  AOI222_X1 U3964 ( .A1(n66), .A2(s_A_SHIFT[5]), .B1(n617), .B2(s_A_SHIFT[13]), 
        .C1(n616), .C2(s_A_SHIFT[21]), .ZN(n662) );
  INV_X1 U3965 ( .A(n315), .ZN(n318) );
  NAND2_X1 U3966 ( .A1(n318), .A2(n317), .ZN(n704) );
  AOI222_X1 U3967 ( .A1(n66), .A2(s_A_SHIFT[1]), .B1(n617), .B2(s_A_SHIFT[9]), 
        .C1(n616), .C2(s_A_SHIFT[17]), .ZN(n316) );
  OAI222_X1 U3968 ( .A1(n677), .A2(n620), .B1(n698), .B2(n662), .C1(n704), 
        .C2(n316), .ZN(n478) );
  AOI22_X1 U3969 ( .A1(n66), .A2(s_A_SHIFT[7]), .B1(n616), .B2(s_A_SHIFT[23]), 
        .ZN(n320) );
  AOI22_X1 U3970 ( .A1(s_A_SHIFT[0]), .A2(n67), .B1(n617), .B2(s_A_SHIFT[15]), 
        .ZN(n319) );
  NAND2_X1 U3971 ( .A1(n320), .A2(n319), .ZN(n688) );
  AOI222_X1 U3972 ( .A1(s_A_SHIFT[22]), .A2(n616), .B1(s_A_SHIFT[6]), .B2(n66), 
        .C1(s_A_SHIFT[14]), .C2(n617), .ZN(n674) );
  INV_X1 U3973 ( .A(n674), .ZN(n475) );
  AOI222_X1 U3974 ( .A1(n66), .A2(s_A_SHIFT[4]), .B1(n617), .B2(s_A_SHIFT[12]), 
        .C1(n616), .C2(s_A_SHIFT[20]), .ZN(n653) );
  OAI21_X1 U3975 ( .B1(n653), .B2(n698), .A(n334), .ZN(n323) );
  AOI222_X1 U3976 ( .A1(n66), .A2(s_A_SHIFT[0]), .B1(n617), .B2(s_A_SHIFT[8]), 
        .C1(n616), .C2(s_A_SHIFT[16]), .ZN(n321) );
  AOI222_X1 U3977 ( .A1(n66), .A2(s_A_SHIFT[2]), .B1(n617), .B2(s_A_SHIFT[10]), 
        .C1(n616), .C2(s_A_SHIFT[18]), .ZN(n477) );
  OAI22_X1 U3978 ( .A1(n321), .A2(n704), .B1(n477), .B2(n677), .ZN(n322) );
  NAND2_X1 U3979 ( .A1(S_B_LOGIC[0]), .A2(s_A_LOGIC[0]), .ZN(n324) );
  NOR2_X1 U3981 ( .A1(n329), .A2(n1432), .ZN(n326) );
  NAND3_X1 U3982 ( .A1(n1417), .A2(n1441), .A3(n1432), .ZN(n327) );
  INV_X1 U3984 ( .A(n617), .ZN(n369) );
  INV_X1 U3985 ( .A(s_A_SHIFT[21]), .ZN(n603) );
  AOI22_X1 U3986 ( .A1(n66), .A2(s_A_SHIFT[13]), .B1(n616), .B2(s_A_SHIFT[29]), 
        .ZN(n336) );
  OAI21_X1 U3987 ( .B1(n369), .B2(n603), .A(n336), .ZN(n337) );
  AOI21_X1 U3988 ( .B1(s_A_SHIFT[6]), .B2(n67), .A(n337), .ZN(n725) );
  AOI22_X1 U3990 ( .A1(n66), .A2(s_A_SHIFT[11]), .B1(s_A_SHIFT[4]), .B2(n67), 
        .ZN(n339) );
  AOI22_X1 U3991 ( .A1(n617), .A2(s_A_SHIFT[19]), .B1(n616), .B2(s_A_SHIFT[27]), .ZN(n338) );
  NAND2_X1 U3992 ( .A1(n339), .A2(n338), .ZN(n723) );
  INV_X1 U3993 ( .A(n723), .ZN(n715) );
  OAI22_X1 U3994 ( .A1(n714), .A2(n725), .B1(n538), .B2(n715), .ZN(n340) );
  INV_X1 U3995 ( .A(n340), .ZN(n364) );
  NAND2_X1 U3996 ( .A1(n686), .A2(n736), .ZN(n713) );
  INV_X1 U3997 ( .A(n713), .ZN(n648) );
  INV_X1 U3998 ( .A(n616), .ZN(n343) );
  INV_X1 U3999 ( .A(s_A_SHIFT[31]), .ZN(n646) );
  AOI22_X1 U4000 ( .A1(s_A_SHIFT[0]), .A2(n643), .B1(s_A_SHIFT[8]), .B2(n67), 
        .ZN(n342) );
  AOI22_X1 U4001 ( .A1(n66), .A2(s_A_SHIFT[15]), .B1(n617), .B2(s_A_SHIFT[23]), 
        .ZN(n341) );
  OAI211_X1 U4002 ( .C1(n343), .C2(n646), .A(n342), .B(n341), .ZN(n717) );
  INV_X1 U4004 ( .A(n728), .ZN(n716) );
  NAND3_X1 U4005 ( .A1(s_SHIFT[1]), .A2(s_A_SHIFT[31]), .A3(n344), .ZN(n551)
         );
  NOR2_X1 U4006 ( .A1(n440), .A2(n551), .ZN(n431) );
  INV_X1 U4007 ( .A(s_A_SHIFT[17]), .ZN(n553) );
  AOI22_X1 U4008 ( .A1(n617), .A2(s_A_SHIFT[25]), .B1(s_A_SHIFT[10]), .B2(n67), 
        .ZN(n345) );
  OAI21_X1 U4009 ( .B1(n59), .B2(n553), .A(n345), .ZN(n346) );
  INV_X1 U4010 ( .A(n444), .ZN(n415) );
  AOI22_X1 U4011 ( .A1(n648), .A2(n717), .B1(n716), .B2(n415), .ZN(n363) );
  INV_X1 U4012 ( .A(s_A_SHIFT[20]), .ZN(n590) );
  AOI22_X1 U4013 ( .A1(n66), .A2(s_A_SHIFT[12]), .B1(s_A_SHIFT[5]), .B2(n67), 
        .ZN(n347) );
  OAI21_X1 U4014 ( .B1(n369), .B2(n590), .A(n347), .ZN(n348) );
  AOI21_X1 U4015 ( .B1(n616), .B2(s_A_SHIFT[28]), .A(n348), .ZN(n699) );
  INV_X1 U4016 ( .A(s_A_SHIFT[14]), .ZN(n403) );
  AOI22_X1 U4017 ( .A1(n616), .A2(s_A_SHIFT[30]), .B1(n67), .B2(s_A_SHIFT[7]), 
        .ZN(n349) );
  OAI21_X1 U4018 ( .B1(n59), .B2(n403), .A(n349), .ZN(n350) );
  AOI21_X1 U4019 ( .B1(n617), .B2(s_A_SHIFT[22]), .A(n350), .ZN(n697) );
  AOI22_X1 U4020 ( .A1(n66), .A2(s_A_SHIFT[10]), .B1(s_A_SHIFT[3]), .B2(n67), 
        .ZN(n352) );
  AOI22_X1 U4021 ( .A1(n617), .A2(s_A_SHIFT[18]), .B1(n616), .B2(s_A_SHIFT[26]), .ZN(n351) );
  NAND2_X1 U4022 ( .A1(n352), .A2(n351), .ZN(n701) );
  INV_X1 U4023 ( .A(n701), .ZN(n353) );
  OAI222_X1 U4024 ( .A1(n677), .A2(n699), .B1(n698), .B2(n697), .C1(n704), 
        .C2(n353), .ZN(n735) );
  INV_X1 U4025 ( .A(S_B_LOGIC[10]), .ZN(n360) );
  NOR3_X1 U4026 ( .A1(s_A_LOGIC[10]), .A2(n360), .A3(n1436), .ZN(n359) );
  INV_X1 U4027 ( .A(s_A_SHIFT[16]), .ZN(n355) );
  AOI22_X1 U4028 ( .A1(s_A_SHIFT[1]), .A2(n643), .B1(s_A_SHIFT[9]), .B2(n67), 
        .ZN(n354) );
  OAI21_X1 U4029 ( .B1(n59), .B2(n355), .A(n354), .ZN(n356) );
  AOI211_X1 U4030 ( .C1(n617), .C2(s_A_SHIFT[24]), .A(n431), .B(n356), .ZN(
        n727) );
  OAI22_X1 U4032 ( .A1(n1406), .A2(n357), .B1(n727), .B2(n1427), .ZN(n358) );
  AOI211_X1 U4033 ( .C1(n1418), .C2(n735), .A(n359), .B(n358), .ZN(n362) );
  OAI221_X1 U4034 ( .B1(S_B_LOGIC[10]), .B2(n1428), .C1(n360), .C2(n1403), .A(
        s_A_LOGIC[10]), .ZN(n361) );
  NAND4_X1 U4035 ( .A1(n364), .A2(n363), .A3(n362), .A4(n361), .ZN(Y[10]) );
  NAND2_X1 U4036 ( .A1(S_B_LOGIC[11]), .A2(s_A_LOGIC[11]), .ZN(n366) );
  OAI221_X1 U4038 ( .B1(n366), .B2(n1402), .C1(S_B_LOGIC[11]), .C2(
        s_A_LOGIC[11]), .A(n365), .ZN(n375) );
  OAI22_X1 U4040 ( .A1(n444), .A2(n1427), .B1(n715), .B2(n1421), .ZN(n373) );
  INV_X1 U4041 ( .A(s_A_SHIFT[26]), .ZN(n565) );
  AOI21_X1 U4042 ( .B1(s_A_SHIFT[3]), .B2(n643), .A(n431), .ZN(n368) );
  AOI22_X1 U4043 ( .A1(n66), .A2(s_A_SHIFT[18]), .B1(s_A_SHIFT[11]), .B2(n67), 
        .ZN(n367) );
  OAI211_X1 U4044 ( .C1(n369), .C2(n565), .A(n368), .B(n367), .ZN(n445) );
  INV_X1 U4045 ( .A(n445), .ZN(n394) );
  OAI22_X1 U4046 ( .A1(n394), .A2(n728), .B1(n697), .B2(n714), .ZN(n372) );
  INV_X1 U4047 ( .A(n717), .ZN(n731) );
  OAI22_X1 U4049 ( .A1(n699), .A2(n538), .B1(n731), .B2(n726), .ZN(n371) );
  OAI22_X1 U4051 ( .A1(n725), .A2(n678), .B1(n727), .B2(n713), .ZN(n370) );
  NOR4_X1 U4052 ( .A1(n373), .A2(n372), .A3(n371), .A4(n370), .ZN(n374) );
  OAI211_X1 U4053 ( .C1(n1405), .C2(n376), .A(n375), .B(n374), .ZN(Y[11]) );
  NAND2_X1 U4054 ( .A1(S_B_LOGIC[12]), .A2(s_A_LOGIC[12]), .ZN(n378) );
  OAI221_X1 U4056 ( .B1(n378), .B2(n1403), .C1(S_B_LOGIC[12]), .C2(
        s_A_LOGIC[12]), .A(n377), .ZN(n386) );
  OAI22_X1 U4057 ( .A1(n394), .A2(n1427), .B1(n699), .B2(n1421), .ZN(n384) );
  INV_X1 U4058 ( .A(s_A_SHIFT[19]), .ZN(n578) );
  AOI22_X1 U4059 ( .A1(n617), .A2(s_A_SHIFT[27]), .B1(s_A_SHIFT[12]), .B2(n67), 
        .ZN(n379) );
  OAI21_X1 U4060 ( .B1(n59), .B2(n578), .A(n379), .ZN(n380) );
  OAI22_X1 U4061 ( .A1(n464), .A2(n728), .B1(n731), .B2(n714), .ZN(n383) );
  OAI22_X1 U4062 ( .A1(n725), .A2(n538), .B1(n727), .B2(n726), .ZN(n382) );
  OAI22_X1 U4063 ( .A1(n444), .A2(n713), .B1(n697), .B2(n678), .ZN(n381) );
  OAI211_X1 U4065 ( .C1(n1406), .C2(n387), .A(n386), .B(n385), .ZN(Y[12]) );
  NAND2_X1 U4066 ( .A1(S_B_LOGIC[13]), .A2(s_A_LOGIC[13]), .ZN(n389) );
  OAI221_X1 U4068 ( .B1(n389), .B2(n1402), .C1(S_B_LOGIC[13]), .C2(
        s_A_LOGIC[13]), .A(n388), .ZN(n398) );
  AOI21_X1 U4069 ( .B1(s_A_SHIFT[5]), .B2(n643), .A(n431), .ZN(n391) );
  AOI22_X1 U4070 ( .A1(n617), .A2(s_A_SHIFT[28]), .B1(s_A_SHIFT[13]), .B2(n67), 
        .ZN(n390) );
  OAI211_X1 U4071 ( .C1(n59), .C2(n590), .A(n391), .B(n390), .ZN(n465) );
  OAI22_X1 U4072 ( .A1(n697), .A2(n704), .B1(n727), .B2(n677), .ZN(n392) );
  AOI21_X1 U4073 ( .B1(n663), .B2(n465), .A(n392), .ZN(n393) );
  OAI21_X1 U4074 ( .B1(n394), .B2(n698), .A(n393), .ZN(n407) );
  OAI22_X1 U4075 ( .A1(n444), .A2(n726), .B1(n731), .B2(n1423), .ZN(n396) );
  OAI22_X1 U4076 ( .A1(n464), .A2(n1427), .B1(n725), .B2(n614), .ZN(n395) );
  AOI211_X1 U4077 ( .C1(n1434), .C2(n407), .A(n396), .B(n395), .ZN(n397) );
  OAI211_X1 U4078 ( .C1(n1406), .C2(n399), .A(n398), .B(n397), .ZN(Y[13]) );
  NAND2_X1 U4079 ( .A1(S_B_LOGIC[14]), .A2(s_A_LOGIC[14]), .ZN(n401) );
  OAI221_X1 U4081 ( .B1(n401), .B2(n1403), .C1(S_B_LOGIC[14]), .C2(
        s_A_LOGIC[14]), .A(n400), .ZN(n409) );
  OAI22_X1 U4082 ( .A1(n464), .A2(n713), .B1(n731), .B2(n538), .ZN(n406) );
  AOI22_X1 U4083 ( .A1(n66), .A2(s_A_SHIFT[21]), .B1(n617), .B2(s_A_SHIFT[29]), 
        .ZN(n402) );
  OAI21_X1 U4084 ( .B1(n403), .B2(n57), .A(n402), .ZN(n404) );
  OAI22_X1 U4085 ( .A1(n502), .A2(n728), .B1(n444), .B2(n714), .ZN(n405) );
  OAI211_X1 U4087 ( .C1(n1406), .C2(n410), .A(n409), .B(n408), .ZN(Y[14]) );
  INV_X1 U4088 ( .A(s_A_SHIFT[22]), .ZN(n629) );
  AOI21_X1 U4089 ( .B1(s_A_SHIFT[7]), .B2(n643), .A(n431), .ZN(n412) );
  AOI22_X1 U4090 ( .A1(n617), .A2(s_A_SHIFT[30]), .B1(n67), .B2(s_A_SHIFT[15]), 
        .ZN(n411) );
  OAI211_X1 U4091 ( .C1(n59), .C2(n629), .A(n412), .B(n411), .ZN(n495) );
  AOI22_X1 U4092 ( .A1(n702), .A2(n445), .B1(n686), .B2(n465), .ZN(n413) );
  OAI21_X1 U4093 ( .B1(n727), .B2(n704), .A(n413), .ZN(n414) );
  AOI21_X1 U4094 ( .B1(n663), .B2(n495), .A(n414), .ZN(n439) );
  INV_X1 U4095 ( .A(n1423), .ZN(n724) );
  INV_X1 U4097 ( .A(n464), .ZN(n451) );
  AOI22_X1 U4098 ( .A1(n724), .A2(n415), .B1(n654), .B2(n451), .ZN(n422) );
  OAI22_X1 U4099 ( .A1(n502), .A2(n1427), .B1(n731), .B2(n614), .ZN(n419) );
  NAND2_X1 U4100 ( .A1(S_B_LOGIC[15]), .A2(s_A_LOGIC[15]), .ZN(n417) );
  OAI211_X1 U4101 ( .C1(S_B_LOGIC[15]), .C2(s_A_LOGIC[15]), .A(n1428), .B(n417), .ZN(n416) );
  OAI21_X1 U4102 ( .B1(n1420), .B2(n417), .A(n416), .ZN(n418) );
  AOI211_X1 U4103 ( .C1(n649), .C2(n420), .A(n419), .B(n418), .ZN(n421) );
  OAI211_X1 U4104 ( .C1(n439), .C2(n695), .A(n422), .B(n421), .ZN(Y[15]) );
  NAND2_X1 U4105 ( .A1(n1398), .A2(S_B_LOGIC[16]), .ZN(n425) );
  OAI22_X1 U4106 ( .A1(n464), .A2(n714), .B1(s_A_LOGIC[16]), .B2(n425), .ZN(
        n426) );
  AOI21_X1 U4107 ( .B1(n75), .B2(S_B_LHI[0]), .A(n426), .ZN(n438) );
  AOI22_X1 U4108 ( .A1(s_A_SHIFT[0]), .A2(n644), .B1(s_A_SHIFT[16]), .B2(n67), 
        .ZN(n429) );
  AOI22_X1 U4109 ( .A1(n66), .A2(s_A_SHIFT[23]), .B1(n617), .B2(s_A_SHIFT[31]), 
        .ZN(n428) );
  NAND2_X1 U4110 ( .A1(n429), .A2(n428), .ZN(n430) );
  INV_X1 U4111 ( .A(n532), .ZN(n517) );
  OAI22_X1 U4112 ( .A1(n502), .A2(n713), .B1(n444), .B2(n538), .ZN(n436) );
  INV_X1 U4113 ( .A(S_B_LOGIC[16]), .ZN(n432) );
  AOI22_X1 U4118 ( .A1(s_A_SHIFT[1]), .A2(n644), .B1(s_A_SHIFT[9]), .B2(n643), 
        .ZN(n443) );
  AOI22_X1 U4119 ( .A1(n66), .A2(s_A_SHIFT[24]), .B1(s_A_SHIFT[17]), .B2(n67), 
        .ZN(n442) );
  AOI21_X1 U4120 ( .B1(n441), .B2(n440), .A(n551), .ZN(n484) );
  INV_X1 U4121 ( .A(n484), .ZN(n539) );
  NAND3_X1 U4122 ( .A1(n443), .A2(n442), .A3(n539), .ZN(n524) );
  INV_X1 U4123 ( .A(n524), .ZN(n460) );
  AOI222_X1 U4124 ( .A1(n445), .A2(n687), .B1(n465), .B2(n702), .C1(n495), 
        .C2(n686), .ZN(n454) );
  INV_X1 U4125 ( .A(s_A_SHIFT[18]), .ZN(n566) );
  AOI22_X1 U4126 ( .A1(s_A_SHIFT[2]), .A2(n644), .B1(s_A_SHIFT[10]), .B2(n643), 
        .ZN(n447) );
  OAI21_X1 U4127 ( .B1(n566), .B2(n57), .A(n447), .ZN(n448) );
  INV_X1 U4128 ( .A(n557), .ZN(n466) );
  OAI22_X1 U4129 ( .A1(n532), .A2(n713), .B1(n502), .B2(n714), .ZN(n456) );
  INV_X1 U4132 ( .A(n538), .ZN(n718) );
  AOI22_X1 U4133 ( .A1(n718), .A2(n451), .B1(n450), .B2(n649), .ZN(n452) );
  INV_X1 U4136 ( .A(S_B_LOGIC[18]), .ZN(n457) );
  OAI221_X1 U4137 ( .B1(S_B_LOGIC[18]), .B2(n58), .C1(n457), .C2(n1402), .A(
        s_A_LOGIC[18]), .ZN(n458) );
  AOI22_X1 U4139 ( .A1(s_A_SHIFT[3]), .A2(n644), .B1(s_A_SHIFT[11]), .B2(n643), 
        .ZN(n461) );
  OAI21_X1 U4140 ( .B1(n578), .B2(n57), .A(n461), .ZN(n462) );
  AOI211_X1 U4141 ( .C1(n66), .C2(s_A_SHIFT[26]), .A(n484), .B(n462), .ZN(n556) );
  AOI222_X1 U4142 ( .A1(n465), .A2(n687), .B1(n495), .B2(n702), .C1(n524), 
        .C2(n686), .ZN(n488) );
  NOR2_X1 U4144 ( .A1(s_A_LOGIC[1]), .A2(n68), .ZN(n467) );
  AOI22_X1 U4145 ( .A1(n467), .A2(S_B_LOGIC[1]), .B1(n666), .B2(n688), .ZN(
        n481) );
  INV_X1 U4146 ( .A(S_B_LOGIC[1]), .ZN(n468) );
  AOI22_X1 U4148 ( .A1(s_A_LOGIC[1]), .A2(n470), .B1(n469), .B2(n649), .ZN(
        n480) );
  INV_X1 U4149 ( .A(s_A_SHIFT[8]), .ZN(n472) );
  AOI22_X1 U4150 ( .A1(n616), .A2(s_A_SHIFT[24]), .B1(s_A_SHIFT[1]), .B2(n67), 
        .ZN(n471) );
  OAI21_X1 U4151 ( .B1(n59), .B2(n472), .A(n471), .ZN(n473) );
  AOI21_X1 U4152 ( .B1(n617), .B2(s_A_SHIFT[16]), .A(n473), .ZN(n705) );
  INV_X1 U4153 ( .A(n663), .ZN(n696) );
  OAI22_X1 U4154 ( .A1(n653), .A2(n677), .B1(n705), .B2(n696), .ZN(n474) );
  AOI21_X1 U4155 ( .B1(n686), .B2(n475), .A(n474), .ZN(n476) );
  OAI21_X1 U4156 ( .B1(n477), .B2(n704), .A(n476), .ZN(n624) );
  AOI22_X1 U4157 ( .A1(n1418), .A2(n478), .B1(n1434), .B2(n624), .ZN(n479) );
  NAND3_X1 U4158 ( .A1(n481), .A2(n480), .A3(n479), .ZN(Y[1]) );
  INV_X1 U4159 ( .A(S_B_LOGIC[20]), .ZN(n487) );
  NOR3_X1 U4160 ( .A1(s_A_LOGIC[20]), .A2(n487), .A3(n1435), .ZN(n486) );
  AOI22_X1 U4161 ( .A1(s_A_SHIFT[4]), .A2(n644), .B1(s_A_SHIFT[12]), .B2(n643), 
        .ZN(n482) );
  OAI21_X1 U4162 ( .B1(n590), .B2(n57), .A(n482), .ZN(n483) );
  OAI22_X1 U4163 ( .A1(n569), .A2(n728), .B1(n556), .B2(n1427), .ZN(n485) );
  AOI211_X1 U4164 ( .C1(S_B_LHI[4]), .C2(n1616), .A(n486), .B(n485), .ZN(n494)
         );
  OAI22_X1 U4166 ( .A1(n532), .A2(n714), .B1(n502), .B2(n538), .ZN(n491) );
  OAI22_X1 U4167 ( .A1(n1405), .A2(n489), .B1(n488), .B2(n711), .ZN(n490) );
  AOI211_X1 U4168 ( .C1(s_A_LOGIC[20]), .C2(n492), .A(n491), .B(n490), .ZN(
        n493) );
  OAI211_X1 U4169 ( .C1(n557), .C2(n713), .A(n494), .B(n493), .ZN(Y[20]) );
  INV_X1 U4170 ( .A(n556), .ZN(n523) );
  AOI222_X1 U4171 ( .A1(n495), .A2(n687), .B1(n524), .B2(n702), .C1(n523), 
        .C2(n686), .ZN(n520) );
  INV_X1 U4172 ( .A(S_B_LOGIC[21]), .ZN(n501) );
  NOR3_X1 U4173 ( .A1(s_A_LOGIC[21]), .A2(n501), .A3(n1435), .ZN(n500) );
  AOI22_X1 U4174 ( .A1(s_A_SHIFT[5]), .A2(n644), .B1(s_A_SHIFT[13]), .B2(n643), 
        .ZN(n497) );
  AOI22_X1 U4175 ( .A1(n66), .A2(s_A_SHIFT[28]), .B1(s_A_SHIFT[21]), .B2(n67), 
        .ZN(n496) );
  NAND3_X1 U4176 ( .A1(n497), .A2(n496), .A3(n539), .ZN(n592) );
  INV_X1 U4177 ( .A(n592), .ZN(n526) );
  OAI22_X1 U4178 ( .A1(n1405), .A2(n498), .B1(n526), .B2(n728), .ZN(n499) );
  AOI211_X1 U4179 ( .C1(S_B_LHI[5]), .C2(n1616), .A(n500), .B(n499), .ZN(n507)
         );
  OAI22_X1 U4181 ( .A1(n569), .A2(n730), .B1(n557), .B2(n726), .ZN(n504) );
  OAI22_X1 U4182 ( .A1(n502), .A2(n614), .B1(n532), .B2(n1423), .ZN(n503) );
  AOI211_X1 U4183 ( .C1(s_A_LOGIC[21]), .C2(n505), .A(n504), .B(n503), .ZN(
        n506) );
  OAI211_X1 U4184 ( .C1(n520), .C2(n695), .A(n507), .B(n506), .ZN(Y[21]) );
  AOI22_X1 U4185 ( .A1(s_A_SHIFT[6]), .A2(n644), .B1(s_A_SHIFT[14]), .B2(n643), 
        .ZN(n508) );
  OAI211_X1 U4186 ( .C1(n57), .C2(n629), .A(n508), .B(n539), .ZN(n509) );
  AOI21_X1 U4187 ( .B1(n66), .B2(s_A_SHIFT[29]), .A(n509), .ZN(n615) );
  INV_X1 U4188 ( .A(n615), .ZN(n594) );
  AOI22_X1 U4189 ( .A1(n716), .A2(n594), .B1(n666), .B2(n592), .ZN(n519) );
  OAI22_X1 U4190 ( .A1(n557), .A2(n714), .B1(n569), .B2(n713), .ZN(n516) );
  NAND2_X1 U4191 ( .A1(S_B_LOGIC[22]), .A2(s_A_LOGIC[22]), .ZN(n511) );
  OAI221_X1 U4193 ( .B1(n511), .B2(n1402), .C1(S_B_LOGIC[22]), .C2(
        s_A_LOGIC[22]), .A(n510), .ZN(n513) );
  NAND2_X1 U4194 ( .A1(n75), .A2(S_B_LHI[6]), .ZN(n512) );
  OAI211_X1 U4195 ( .C1(n1405), .C2(n514), .A(n513), .B(n512), .ZN(n515) );
  OAI211_X1 U4197 ( .C1(n520), .C2(n711), .A(n519), .B(n518), .ZN(Y[22]) );
  AOI22_X1 U4198 ( .A1(s_A_SHIFT[15]), .A2(n643), .B1(s_A_SHIFT[7]), .B2(n644), 
        .ZN(n522) );
  AOI22_X1 U4199 ( .A1(n66), .A2(s_A_SHIFT[30]), .B1(n67), .B2(s_A_SHIFT[23]), 
        .ZN(n521) );
  NAND3_X1 U4200 ( .A1(n522), .A2(n521), .A3(n539), .ZN(n604) );
  AOI22_X1 U4201 ( .A1(n687), .A2(n524), .B1(n702), .B2(n523), .ZN(n525) );
  OAI21_X1 U4202 ( .B1(n526), .B2(n698), .A(n525), .ZN(n527) );
  AOI21_X1 U4203 ( .B1(n663), .B2(n604), .A(n527), .ZN(n550) );
  NAND2_X1 U4204 ( .A1(n1399), .A2(s_A_LOGIC[23]), .ZN(n528) );
  OAI22_X1 U4205 ( .A1(S_B_LOGIC[23]), .A2(n528), .B1(n557), .B2(n1423), .ZN(
        n529) );
  AOI21_X1 U4206 ( .B1(n1616), .B2(S_B_LHI[7]), .A(n529), .ZN(n537) );
  INV_X1 U4207 ( .A(s_A_LOGIC[23]), .ZN(n530) );
  AOI22_X1 U4208 ( .A1(s_A_LOGIC[23]), .A2(n1420), .B1(n68), .B2(n530), .ZN(
        n535) );
  OAI22_X1 U4209 ( .A1(n569), .A2(n726), .B1(n615), .B2(n730), .ZN(n534) );
  OAI22_X1 U4210 ( .A1(n532), .A2(n1421), .B1(n732), .B2(n531), .ZN(n533) );
  AOI211_X1 U4211 ( .C1(S_B_LOGIC[23]), .C2(n535), .A(n534), .B(n533), .ZN(
        n536) );
  OAI211_X1 U4212 ( .C1(n550), .C2(n695), .A(n537), .B(n536), .ZN(Y[23]) );
  OAI22_X1 U4213 ( .A1(n557), .A2(n538), .B1(n615), .B2(n713), .ZN(n548) );
  AOI22_X1 U4214 ( .A1(s_A_SHIFT[8]), .A2(n644), .B1(s_A_SHIFT[16]), .B2(n643), 
        .ZN(n540) );
  OAI211_X1 U4215 ( .C1(n646), .C2(n59), .A(n540), .B(n539), .ZN(n541) );
  AOI21_X1 U4216 ( .B1(n67), .B2(s_A_SHIFT[24]), .A(n541), .ZN(n588) );
  OAI22_X1 U4217 ( .A1(n569), .A2(n714), .B1(n588), .B2(n728), .ZN(n547) );
  NAND2_X1 U4218 ( .A1(s_A_LOGIC[24]), .A2(S_B_LOGIC[24]), .ZN(n545) );
  AOI22_X1 U4219 ( .A1(S_B_LHI[8]), .A2(n1616), .B1(\intadd_0/SUM[0] ), .B2(
        n649), .ZN(n543) );
  OAI211_X1 U4220 ( .C1(s_A_LOGIC[24]), .C2(S_B_LOGIC[24]), .A(n1399), .B(n545), .ZN(n542) );
  OAI211_X1 U4221 ( .C1(n545), .C2(n1420), .A(n543), .B(n542), .ZN(n546) );
  NOR3_X1 U4222 ( .A1(n548), .A2(n547), .A3(n546), .ZN(n549) );
  OAI21_X1 U4223 ( .B1(n550), .B2(n711), .A(n549), .ZN(Y[24]) );
  AOI22_X1 U4224 ( .A1(S_B_LHI[9]), .A2(n1616), .B1(\intadd_0/SUM[1] ), .B2(
        n649), .ZN(n564) );
  AOI22_X1 U4225 ( .A1(n702), .A2(n592), .B1(n686), .B2(n604), .ZN(n555) );
  INV_X1 U4226 ( .A(n643), .ZN(n630) );
  AOI22_X1 U4227 ( .A1(s_A_SHIFT[9]), .A2(n644), .B1(n67), .B2(s_A_SHIFT[25]), 
        .ZN(n552) );
  AOI21_X1 U4228 ( .B1(S_B_SHIFT[4]), .B2(S_B_SHIFT[3]), .A(n551), .ZN(n568)
         );
  INV_X1 U4229 ( .A(n568), .ZN(n645) );
  OAI211_X1 U4230 ( .C1(n630), .C2(n553), .A(n552), .B(n645), .ZN(n651) );
  NAND2_X1 U4231 ( .A1(n663), .A2(n651), .ZN(n554) );
  OAI211_X1 U4232 ( .C1(n556), .C2(n704), .A(n555), .B(n554), .ZN(n570) );
  OAI22_X1 U4233 ( .A1(n615), .A2(n726), .B1(n569), .B2(n678), .ZN(n559) );
  OAI22_X1 U4234 ( .A1(n557), .A2(n1421), .B1(n588), .B2(n1427), .ZN(n558) );
  AOI211_X1 U4235 ( .C1(n1434), .C2(n570), .A(n559), .B(n558), .ZN(n563) );
  NAND2_X1 U4236 ( .A1(s_A_LOGIC[25]), .A2(S_B_LOGIC[25]), .ZN(n560) );
  OAI211_X1 U4237 ( .C1(s_A_LOGIC[25]), .C2(S_B_LOGIC[25]), .A(n1428), .B(n560), .ZN(n562) );
  NAND3_X1 U4238 ( .A1(n1403), .A2(s_A_LOGIC[25]), .A3(S_B_LOGIC[25]), .ZN(
        n561) );
  NAND4_X1 U4239 ( .A1(n564), .A2(n563), .A3(n562), .A4(n561), .ZN(Y[25]) );
  AND2_X1 U4240 ( .A1(s_A_LOGIC[26]), .A2(S_B_LOGIC[26]), .ZN(n576) );
  OAI21_X1 U4241 ( .B1(s_A_LOGIC[26]), .B2(S_B_LOGIC[26]), .A(n1399), .ZN(n575) );
  OAI22_X1 U4242 ( .A1(n566), .A2(n630), .B1(n57), .B2(n565), .ZN(n567) );
  AOI211_X1 U4243 ( .C1(n644), .C2(s_A_SHIFT[10]), .A(n568), .B(n567), .ZN(
        n591) );
  AOI22_X1 U4244 ( .A1(S_B_LHI[10]), .A2(n1616), .B1(\intadd_0/SUM[2] ), .B2(
        n649), .ZN(n572) );
  OAI222_X1 U4245 ( .A1(n677), .A2(n615), .B1(n698), .B2(n588), .C1(n704), 
        .C2(n569), .ZN(n582) );
  AOI22_X1 U4246 ( .A1(n1418), .A2(n570), .B1(n1434), .B2(n582), .ZN(n571) );
  OAI211_X1 U4247 ( .C1(n591), .C2(n728), .A(n572), .B(n571), .ZN(n573) );
  AOI21_X1 U4248 ( .B1(n1402), .B2(n576), .A(n573), .ZN(n574) );
  OAI21_X1 U4249 ( .B1(n576), .B2(n575), .A(n574), .ZN(Y[26]) );
  INV_X1 U4250 ( .A(n714), .ZN(n665) );
  AOI22_X1 U4251 ( .A1(n665), .A2(n604), .B1(n718), .B2(n592), .ZN(n587) );
  AOI22_X1 U4252 ( .A1(s_A_SHIFT[11]), .A2(n644), .B1(n67), .B2(s_A_SHIFT[27]), 
        .ZN(n577) );
  OAI211_X1 U4253 ( .C1(n630), .C2(n578), .A(n577), .B(n645), .ZN(n650) );
  AOI22_X1 U4254 ( .A1(n648), .A2(n651), .B1(n1433), .B2(n650), .ZN(n586) );
  INV_X1 U4255 ( .A(S_B_LOGIC[27]), .ZN(n583) );
  NOR3_X1 U4256 ( .A1(s_A_LOGIC[27]), .A2(n583), .A3(n68), .ZN(n581) );
  AOI22_X1 U4257 ( .A1(S_B_LHI[11]), .A2(n75), .B1(\intadd_0/SUM[3] ), .B2(
        n649), .ZN(n579) );
  OAI21_X1 U4258 ( .B1(n591), .B2(n1427), .A(n579), .ZN(n580) );
  AOI211_X1 U4259 ( .C1(n1419), .C2(n582), .A(n581), .B(n580), .ZN(n585) );
  OAI221_X1 U4260 ( .B1(S_B_LOGIC[27]), .B2(n1428), .C1(n583), .C2(n1402), .A(
        s_A_LOGIC[27]), .ZN(n584) );
  NAND4_X1 U4261 ( .A1(n587), .A2(n586), .A3(n585), .A4(n584), .ZN(Y[27]) );
  INV_X1 U4262 ( .A(n588), .ZN(n634) );
  AOI22_X1 U4263 ( .A1(s_A_SHIFT[12]), .A2(n644), .B1(n67), .B2(s_A_SHIFT[28]), 
        .ZN(n589) );
  OAI211_X1 U4264 ( .C1(n630), .C2(n590), .A(n589), .B(n645), .ZN(n631) );
  INV_X1 U4265 ( .A(n591), .ZN(n633) );
  AOI222_X1 U4266 ( .A1(n634), .A2(n702), .B1(n631), .B2(n663), .C1(n633), 
        .C2(n686), .ZN(n611) );
  INV_X1 U4267 ( .A(n1421), .ZN(n722) );
  AOI22_X1 U4268 ( .A1(n722), .A2(n592), .B1(n724), .B2(n604), .ZN(n601) );
  NAND2_X1 U4269 ( .A1(s_A_LOGIC[28]), .A2(S_B_LOGIC[28]), .ZN(n595) );
  INV_X1 U4270 ( .A(n595), .ZN(n593) );
  AOI22_X1 U4271 ( .A1(n1403), .A2(n593), .B1(n666), .B2(n650), .ZN(n599) );
  AOI22_X1 U4272 ( .A1(S_B_LHI[12]), .A2(n1616), .B1(\intadd_0/SUM[4] ), .B2(
        n649), .ZN(n598) );
  AOI22_X1 U4273 ( .A1(n718), .A2(n594), .B1(n654), .B2(n651), .ZN(n597) );
  OAI211_X1 U4274 ( .C1(s_A_LOGIC[28]), .C2(S_B_LOGIC[28]), .A(n1399), .B(n595), .ZN(n596) );
  AND4_X1 U4275 ( .A1(n599), .A2(n598), .A3(n597), .A4(n596), .ZN(n600) );
  OAI211_X1 U4276 ( .C1(n611), .C2(n695), .A(n601), .B(n600), .ZN(Y[28]) );
  AOI22_X1 U4277 ( .A1(s_A_SHIFT[13]), .A2(n644), .B1(n67), .B2(s_A_SHIFT[29]), 
        .ZN(n602) );
  OAI211_X1 U4278 ( .C1(n630), .C2(n603), .A(n602), .B(n645), .ZN(n647) );
  AOI22_X1 U4279 ( .A1(n663), .A2(n647), .B1(n686), .B2(n650), .ZN(n606) );
  AOI22_X1 U4280 ( .A1(n687), .A2(n604), .B1(n702), .B2(n651), .ZN(n605) );
  NAND2_X1 U4281 ( .A1(n606), .A2(n605), .ZN(n637) );
  AOI22_X1 U4282 ( .A1(S_B_LHI[13]), .A2(n75), .B1(\intadd_0/SUM[5] ), .B2(
        n649), .ZN(n610) );
  NAND2_X1 U4283 ( .A1(S_B_LOGIC[29]), .A2(s_A_LOGIC[29]), .ZN(n608) );
  OAI221_X1 U4285 ( .B1(n608), .B2(n1402), .C1(S_B_LOGIC[29]), .C2(
        s_A_LOGIC[29]), .A(n607), .ZN(n609) );
  OAI211_X1 U4286 ( .C1(n611), .C2(n711), .A(n610), .B(n609), .ZN(n612) );
  AOI21_X1 U4287 ( .B1(n1434), .B2(n637), .A(n612), .ZN(n613) );
  OAI21_X1 U4288 ( .B1(n615), .B2(n1421), .A(n613), .ZN(Y[29]) );
  AOI22_X1 U4289 ( .A1(n66), .A2(s_A_SHIFT[9]), .B1(s_A_SHIFT[2]), .B2(n67), 
        .ZN(n619) );
  AOI22_X1 U4290 ( .A1(n617), .A2(s_A_SHIFT[17]), .B1(n616), .B2(s_A_SHIFT[25]), .ZN(n618) );
  NAND2_X1 U4291 ( .A1(n619), .A2(n618), .ZN(n721) );
  OAI22_X1 U4292 ( .A1(n662), .A2(n677), .B1(n620), .B2(n704), .ZN(n621) );
  AOI21_X1 U4293 ( .B1(n663), .B2(n721), .A(n621), .ZN(n661) );
  INV_X1 U4294 ( .A(S_B_LOGIC[2]), .ZN(n625) );
  NOR3_X1 U4295 ( .A1(s_A_LOGIC[2]), .A2(n625), .A3(n1436), .ZN(n623) );
  INV_X1 U4296 ( .A(n688), .ZN(n679) );
  OAI22_X1 U4297 ( .A1(n679), .A2(n713), .B1(n732), .B2(\intadd_1/SUM[0] ), 
        .ZN(n622) );
  AOI211_X1 U4298 ( .C1(n1419), .C2(n624), .A(n623), .B(n622), .ZN(n627) );
  OAI221_X1 U4299 ( .B1(S_B_LOGIC[2]), .B2(n1428), .C1(n625), .C2(n1402), .A(
        s_A_LOGIC[2]), .ZN(n626) );
  OAI211_X1 U4300 ( .C1(n661), .C2(n1397), .A(n627), .B(n626), .ZN(Y[2]) );
  AOI22_X1 U4301 ( .A1(S_B_LHI[14]), .A2(n1616), .B1(\intadd_0/SUM[6] ), .B2(
        n649), .ZN(n642) );
  AOI22_X1 U4302 ( .A1(s_A_SHIFT[14]), .A2(n644), .B1(n67), .B2(s_A_SHIFT[30]), 
        .ZN(n628) );
  OAI211_X1 U4303 ( .C1(n630), .C2(n629), .A(n628), .B(n645), .ZN(n632) );
  AOI22_X1 U4304 ( .A1(n663), .A2(n632), .B1(n686), .B2(n631), .ZN(n636) );
  AOI22_X1 U4305 ( .A1(n687), .A2(n634), .B1(n702), .B2(n633), .ZN(n635) );
  NAND2_X1 U4306 ( .A1(n636), .A2(n635), .ZN(n652) );
  AOI22_X1 U4307 ( .A1(n1419), .A2(n637), .B1(n1434), .B2(n652), .ZN(n641) );
  INV_X1 U4308 ( .A(S_B_LOGIC[30]), .ZN(n638) );
  OAI221_X1 U4309 ( .B1(S_B_LOGIC[30]), .B2(n1399), .C1(n638), .C2(n1402), .A(
        s_A_LOGIC[30]), .ZN(n640) );
  OR3_X1 U4310 ( .A1(n638), .A2(n1436), .A3(s_A_LOGIC[30]), .ZN(n639) );
  NAND4_X1 U4311 ( .A1(n642), .A2(n641), .A3(n640), .A4(n639), .ZN(Y[30]) );
  OAI222_X1 U4312 ( .A1(n677), .A2(n674), .B1(n698), .B2(n705), .C1(n704), 
        .C2(n653), .ZN(n672) );
  NAND2_X1 U4314 ( .A1(S_B_LOGIC[3]), .A2(s_A_LOGIC[3]), .ZN(n656) );
  INV_X1 U4320 ( .A(n662), .ZN(n664) );
  AOI222_X1 U4321 ( .A1(n664), .A2(n687), .B1(n723), .B2(n663), .C1(n721), 
        .C2(n686), .ZN(n685) );
  AOI22_X1 U4322 ( .A1(n666), .A2(n701), .B1(n665), .B2(n688), .ZN(n670) );
  NAND2_X1 U4323 ( .A1(S_B_LOGIC[4]), .A2(s_A_LOGIC[4]), .ZN(n668) );
  OAI221_X1 U4325 ( .B1(n668), .B2(n1402), .C1(S_B_LOGIC[4]), .C2(s_A_LOGIC[4]), .A(n667), .ZN(n669) );
  OAI211_X1 U4326 ( .C1(n1405), .C2(\intadd_1/SUM[2] ), .A(n670), .B(n669), 
        .ZN(n671) );
  AOI21_X1 U4327 ( .B1(n1419), .B2(n672), .A(n671), .ZN(n673) );
  OAI21_X1 U4328 ( .B1(n685), .B2(n1397), .A(n673), .ZN(Y[4]) );
  OAI22_X1 U4329 ( .A1(n674), .A2(n704), .B1(n699), .B2(n696), .ZN(n675) );
  AOI21_X1 U4330 ( .B1(n686), .B2(n701), .A(n675), .ZN(n676) );
  OAI21_X1 U4331 ( .B1(n705), .B2(n677), .A(n676), .ZN(n691) );
  INV_X1 U4332 ( .A(S_B_LOGIC[5]), .ZN(n682) );
  NOR3_X1 U4333 ( .A1(s_A_LOGIC[5]), .A2(n682), .A3(n68), .ZN(n681) );
  OAI22_X1 U4334 ( .A1(n679), .A2(n1423), .B1(n732), .B2(\intadd_1/SUM[3] ), 
        .ZN(n680) );
  AOI211_X1 U4335 ( .C1(n1434), .C2(n691), .A(n681), .B(n680), .ZN(n684) );
  OAI221_X1 U4336 ( .B1(S_B_LOGIC[5]), .B2(n1399), .C1(n682), .C2(n1403), .A(
        s_A_LOGIC[5]), .ZN(n683) );
  OAI211_X1 U4337 ( .C1(n685), .C2(n711), .A(n684), .B(n683), .ZN(Y[5]) );
  AOI222_X1 U4338 ( .A1(n688), .A2(n687), .B1(n721), .B2(n702), .C1(n723), 
        .C2(n686), .ZN(n712) );
  INV_X1 U4339 ( .A(S_B_LOGIC[6]), .ZN(n692) );
  NOR3_X1 U4340 ( .A1(s_A_LOGIC[6]), .A2(n692), .A3(n1436), .ZN(n690) );
  OAI22_X1 U4341 ( .A1(n1406), .A2(\intadd_1/SUM[4] ), .B1(n725), .B2(n728), 
        .ZN(n689) );
  AOI211_X1 U4342 ( .C1(n1418), .C2(n691), .A(n689), .B(n690), .ZN(n694) );
  OAI221_X1 U4343 ( .B1(S_B_LOGIC[6]), .B2(n1428), .C1(n692), .C2(n1402), .A(
        s_A_LOGIC[6]), .ZN(n693) );
  OAI211_X1 U4344 ( .C1(n712), .C2(n1397), .A(n694), .B(n693), .ZN(Y[6]) );
  OAI22_X1 U4345 ( .A1(n699), .A2(n698), .B1(n697), .B2(n696), .ZN(n700) );
  AOI21_X1 U4346 ( .B1(n702), .B2(n701), .A(n700), .ZN(n703) );
  OAI21_X1 U4347 ( .B1(n705), .B2(n704), .A(n703), .ZN(n719) );
  INV_X1 U4348 ( .A(S_B_LOGIC[7]), .ZN(n708) );
  NOR3_X1 U4349 ( .A1(s_A_LOGIC[7]), .A2(n708), .A3(n68), .ZN(n707) );
  OAI22_X1 U4350 ( .A1(n732), .A2(\intadd_1/SUM[5] ), .B1(n725), .B2(n1427), 
        .ZN(n706) );
  AOI211_X1 U4351 ( .C1(n1434), .C2(n719), .A(n707), .B(n706), .ZN(n710) );
  OAI221_X1 U4352 ( .B1(S_B_LOGIC[7]), .B2(n1428), .C1(n708), .C2(n1403), .A(
        s_A_LOGIC[7]), .ZN(n709) );
  OAI211_X1 U4353 ( .C1(n712), .C2(n711), .A(n710), .B(n709), .ZN(Y[7]) );
  AOI22_X1 U4354 ( .A1(n724), .A2(n723), .B1(n722), .B2(n721), .ZN(n742) );
  OAI22_X1 U4355 ( .A1(n728), .A2(n727), .B1(n726), .B2(n725), .ZN(n729) );
  INV_X1 U4356 ( .A(n729), .ZN(n741) );
  INV_X1 U4357 ( .A(s_A_LOGIC[9]), .ZN(n738) );
  NOR3_X1 U4358 ( .A1(S_B_LOGIC[9]), .A2(n738), .A3(n1435), .ZN(n734) );
  OAI22_X1 U4359 ( .A1(n1406), .A2(\intadd_1/SUM[7] ), .B1(n731), .B2(n1427), 
        .ZN(n733) );
  AOI211_X1 U4360 ( .C1(n1434), .C2(n735), .A(n734), .B(n733), .ZN(n740) );
  OAI221_X1 U4361 ( .B1(s_A_LOGIC[9]), .B2(n1399), .C1(n738), .C2(n1402), .A(
        S_B_LOGIC[9]), .ZN(n739) );
  NAND4_X1 U4362 ( .A1(n742), .A2(n741), .A3(n740), .A4(n739), .ZN(Y[9]) );
  XNOR2_X1 U4363 ( .A(S_B_ADDER[24]), .B(n77), .ZN(\intadd_0/B[0] ) );
  XNOR2_X1 U4364 ( .A(S_B_ADDER[25]), .B(n77), .ZN(\intadd_0/B[1] ) );
  XNOR2_X1 U4365 ( .A(S_B_ADDER[26]), .B(n77), .ZN(\intadd_0/B[2] ) );
  XNOR2_X1 U4366 ( .A(S_B_ADDER[27]), .B(n77), .ZN(\intadd_0/B[3] ) );
  XNOR2_X1 U4367 ( .A(S_B_ADDER[28]), .B(n77), .ZN(\intadd_0/B[4] ) );
  XNOR2_X1 U4368 ( .A(S_B_ADDER[29]), .B(n77), .ZN(\intadd_0/B[5] ) );
  XNOR2_X1 U4369 ( .A(S_B_ADDER[30]), .B(n77), .ZN(\intadd_0/B[6] ) );
  XNOR2_X1 U4370 ( .A(S_B_ADDER[31]), .B(n77), .ZN(\intadd_0/B[7] ) );
  AOI22_X1 U4371 ( .A1(n754), .A2(n753), .B1(n744), .B2(n743), .ZN(n756) );
  INV_X1 U4372 ( .A(n745), .ZN(n751) );
  OAI21_X1 U4373 ( .B1(n24), .B2(n747), .A(n746), .ZN(n750) );
  OAI22_X1 U4374 ( .A1(n751), .A2(n750), .B1(n749), .B2(n748), .ZN(n752) );
  OAI21_X1 U4375 ( .B1(n754), .B2(n753), .A(n752), .ZN(n755) );
  AOI22_X1 U4376 ( .A1(n757), .A2(s_A_ADDER[22]), .B1(n756), .B2(n755), .ZN(
        n760) );
  NAND2_X1 U4377 ( .A1(n758), .A2(s_A_ADDER[23]), .ZN(n759) );
  OAI21_X1 U4378 ( .B1(n761), .B2(n760), .A(n759), .ZN(\intadd_0/CI ) );
  AOI21_X1 U4379 ( .B1(n77), .B2(n763), .A(n762), .ZN(n764) );
  AOI222_X1 U4380 ( .A1(s_A_ADDER[1]), .A2(n765), .B1(s_A_ADDER[1]), .B2(n764), 
        .C1(n765), .C2(n764), .ZN(\intadd_1/B[0] ) );
  XNOR2_X1 U4381 ( .A(\ADD_SUB/carry_ST[0] ), .B(S_B_ADDER[3]), .ZN(
        \intadd_1/B[1] ) );
  XNOR2_X1 U4382 ( .A(\ADD_SUB/carry_ST[0] ), .B(S_B_ADDER[4]), .ZN(
        \intadd_1/B[2] ) );
  XNOR2_X1 U4383 ( .A(n76), .B(S_B_ADDER[5]), .ZN(\intadd_1/B[3] ) );
  XNOR2_X1 U4384 ( .A(\ADD_SUB/carry_ST[0] ), .B(S_B_ADDER[6]), .ZN(
        \intadd_1/B[4] ) );
  XNOR2_X1 U4385 ( .A(n76), .B(S_B_ADDER[7]), .ZN(\intadd_1/B[5] ) );
  XNOR2_X1 U4386 ( .A(\ADD_SUB/carry_ST[0] ), .B(S_B_ADDER[8]), .ZN(
        \intadd_1/B[6] ) );
  XNOR2_X1 U4387 ( .A(n76), .B(S_B_ADDER[9]), .ZN(\intadd_1/B[7] ) );
  XNOR2_X1 U4388 ( .A(\ADD_SUB/carry_ST[0] ), .B(S_B_ADDER[2]), .ZN(
        \intadd_1/CI ) );
  NOR2_X1 U4389 ( .A1(n766), .A2(n945), .ZN(n768) );
  INV_X1 U4390 ( .A(n1068), .ZN(n981) );
  OAI22_X1 U4391 ( .A1(n941), .A2(n981), .B1(n936), .B2(n1087), .ZN(n767) );
  AOI211_X1 U4392 ( .C1(n948), .C2(s_A_MULT[8]), .A(n768), .B(n767), .ZN(
        \intadd_10/A[0] ) );
  INV_X1 U4393 ( .A(n1160), .ZN(n1002) );
  NAND3_X1 U4394 ( .A1(S_B_MULT[11]), .A2(n1161), .A3(n816), .ZN(n1252) );
  NAND2_X1 U4395 ( .A1(n1002), .A2(n1252), .ZN(n769) );
  AOI222_X1 U4396 ( .A1(n769), .A2(\MULT/SHIFTERi_0/N19 ), .B1(n1159), .B2(
        n1307), .C1(s_A_MULT[1]), .C2(n1085), .ZN(n778) );
  AOI22_X1 U4397 ( .A1(n1070), .A2(s_A_MULT[3]), .B1(n1073), .B2(s_A_MULT[2]), 
        .ZN(n770) );
  OAI21_X1 U4398 ( .B1(n1041), .B2(n934), .A(n770), .ZN(n771) );
  AOI21_X1 U4399 ( .B1(n908), .B2(n56), .A(n771), .ZN(n777) );
  AOI22_X1 U4400 ( .A1(s_A_MULT[5]), .A2(n1048), .B1(s_A_MULT[4]), .B2(n1076), 
        .ZN(n772) );
  OAI21_X1 U4401 ( .B1(n1046), .B2(n988), .A(n772), .ZN(n773) );
  AOI21_X1 U4402 ( .B1(n959), .B2(n1075), .A(n773), .ZN(n776) );
  OAI21_X1 U4403 ( .B1(n1262), .B2(n1258), .A(\MULT/SHIFTERi_0/N19 ), .ZN(
        n1147) );
  XNOR2_X1 U4404 ( .A(n1148), .B(n1147), .ZN(\intadd_10/A[2] ) );
  AOI22_X1 U4405 ( .A1(s_A_MULT[5]), .A2(n968), .B1(n967), .B2(n1089), .ZN(
        n774) );
  OAI21_X1 U4406 ( .B1(n988), .B2(n1056), .A(n774), .ZN(n775) );
  AOI21_X1 U4407 ( .B1(s_A_MULT[6]), .B2(n966), .A(n775), .ZN(\intadd_10/B[0] ) );
  FA_X1 U4408 ( .A(n778), .B(n777), .CI(n776), .CO(n1148), .S(\intadd_10/B[1] ) );
  AOI21_X1 U4409 ( .B1(s_A_MULT[10]), .B2(n779), .A(n824), .ZN(n1171) );
  AOI222_X1 U4410 ( .A1(s_A_MULT[10]), .A2(n1309), .B1(n1308), .B2(n1171), 
        .C1(n55), .C2(n979), .ZN(\intadd_10/CI ) );
  INV_X1 U4411 ( .A(n1087), .ZN(n920) );
  AOI222_X1 U4412 ( .A1(s_A_MULT[8]), .A2(n1309), .B1(n1308), .B2(n1068), .C1(
        n55), .C2(n920), .ZN(\intadd_11/A[0] ) );
  NOR2_X1 U4413 ( .A1(n1073), .A2(n56), .ZN(n780) );
  INV_X1 U4414 ( .A(n1070), .ZN(n999) );
  OAI222_X1 U4415 ( .A1(n838), .A2(n1041), .B1(n797), .B2(n780), .C1(n999), 
        .C2(n910), .ZN(n783) );
  AOI22_X1 U4416 ( .A1(s_A_MULT[3]), .A2(n1048), .B1(s_A_MULT[2]), .B2(n1076), 
        .ZN(n782) );
  NAND2_X1 U4417 ( .A1(n908), .A2(n1075), .ZN(n781) );
  OAI211_X1 U4418 ( .C1(n934), .C2(n1046), .A(n782), .B(n781), .ZN(n784) );
  NAND2_X1 U4419 ( .A1(n783), .A2(n784), .ZN(\intadd_11/B[2] ) );
  OAI21_X1 U4420 ( .B1(n784), .B2(n783), .A(\intadd_11/B[2] ), .ZN(
        \intadd_11/A[1] ) );
  FA_X1 U4421 ( .A(\intadd_10/SUM[0] ), .B(n786), .CI(n785), .CO(n184), .S(
        \intadd_11/A[2] ) );
  NOR2_X1 U4422 ( .A1(n941), .A2(n922), .ZN(n789) );
  OAI22_X1 U4423 ( .A1(n787), .A2(n945), .B1(n988), .B2(n936), .ZN(n788) );
  AOI211_X1 U4424 ( .C1(n948), .C2(s_A_MULT[6]), .A(n789), .B(n788), .ZN(
        \intadd_11/B[0] ) );
  FA_X1 U4425 ( .A(n792), .B(n791), .CI(n790), .CO(n786), .S(\intadd_11/B[1] )
         );
  AOI22_X1 U4426 ( .A1(s_A_MULT[4]), .A2(n966), .B1(n967), .B2(n959), .ZN(n793) );
  OAI21_X1 U4427 ( .B1(n934), .B2(n1056), .A(n793), .ZN(n794) );
  AOI21_X1 U4428 ( .B1(s_A_MULT[3]), .B2(n968), .A(n794), .ZN(\intadd_11/CI )
         );
  AOI22_X1 U4429 ( .A1(s_A_MULT[3]), .A2(n966), .B1(n967), .B2(n899), .ZN(n795) );
  OAI21_X1 U4430 ( .B1(n902), .B2(n1056), .A(n795), .ZN(n796) );
  AOI21_X1 U4431 ( .B1(s_A_MULT[2]), .B2(n968), .A(n796), .ZN(\intadd_12/A[0] ) );
  AOI21_X1 U4432 ( .B1(n999), .B2(n1041), .A(n797), .ZN(n801) );
  AOI22_X1 U4433 ( .A1(s_A_MULT[1]), .A2(n1076), .B1(s_A_MULT[2]), .B2(n1048), 
        .ZN(n799) );
  NAND2_X1 U4434 ( .A1(n1307), .A2(n1075), .ZN(n798) );
  OAI211_X1 U4435 ( .C1(n902), .C2(n1046), .A(n799), .B(n798), .ZN(n800) );
  NAND2_X1 U4436 ( .A1(n801), .A2(n800), .ZN(\intadd_12/A[2] ) );
  OAI21_X1 U4437 ( .B1(n801), .B2(n800), .A(\intadd_12/A[2] ), .ZN(
        \intadd_12/A[1] ) );
  AOI222_X1 U4438 ( .A1(s_A_MULT[7]), .A2(n1309), .B1(n1308), .B2(n920), .C1(
        n1089), .C2(n55), .ZN(\intadd_12/B[0] ) );
  INV_X1 U4439 ( .A(s_A_MULT[4]), .ZN(n802) );
  NOR2_X1 U4440 ( .A1(n802), .A2(n945), .ZN(n804) );
  OAI22_X1 U4441 ( .A1(n941), .A2(n988), .B1(n833), .B2(n936), .ZN(n803) );
  AOI211_X1 U4442 ( .C1(n948), .C2(s_A_MULT[5]), .A(n804), .B(n803), .ZN(
        \intadd_12/CI ) );
  AOI22_X1 U4443 ( .A1(s_A_MULT[6]), .A2(n968), .B1(n967), .B2(n920), .ZN(n805) );
  OAI21_X1 U4444 ( .B1(n922), .B2(n1056), .A(n805), .ZN(n806) );
  AOI21_X1 U4445 ( .B1(s_A_MULT[7]), .B2(n966), .A(n806), .ZN(\intadd_2/A[0] )
         );
  AOI22_X1 U4446 ( .A1(s_A_MULT[6]), .A2(n1048), .B1(s_A_MULT[5]), .B2(n1076), 
        .ZN(n807) );
  OAI21_X1 U4447 ( .B1(n1046), .B2(n922), .A(n807), .ZN(n808) );
  AOI21_X1 U4448 ( .B1(n831), .B2(n1075), .A(n808), .ZN(n815) );
  AOI22_X1 U4449 ( .A1(n1073), .A2(s_A_MULT[3]), .B1(n1069), .B2(n959), .ZN(
        n809) );
  OAI21_X1 U4450 ( .B1(n934), .B2(n53), .A(n809), .ZN(n810) );
  AOI21_X1 U4451 ( .B1(n1070), .B2(s_A_MULT[4]), .A(n810), .ZN(n814) );
  AOI22_X1 U4452 ( .A1(s_A_MULT[2]), .A2(n1085), .B1(n1159), .B2(n908), .ZN(
        n811) );
  OAI21_X1 U4453 ( .B1(n838), .B2(n1252), .A(n811), .ZN(n812) );
  AOI21_X1 U4454 ( .B1(s_A_MULT[1]), .B2(n1160), .A(n812), .ZN(n813) );
  FA_X1 U4455 ( .A(n815), .B(n814), .CI(n813), .CO(n820), .S(\intadd_2/A[1] )
         );
  INV_X1 U4456 ( .A(n1259), .ZN(n1235) );
  NOR2_X1 U4457 ( .A1(S_B_MULT[11]), .A2(S_B_MULT[12]), .ZN(n817) );
  NAND3_X1 U4458 ( .A1(S_B_MULT[13]), .A2(n817), .A3(n816), .ZN(n1231) );
  NAND2_X1 U4459 ( .A1(n1235), .A2(n1231), .ZN(n818) );
  AOI222_X1 U4460 ( .A1(n818), .A2(\MULT/SHIFTERi_0/N19 ), .B1(n1258), .B2(
        n1307), .C1(s_A_MULT[1]), .C2(n1262), .ZN(n819) );
  OR2_X1 U4461 ( .A1(n820), .A2(n819), .ZN(\intadd_2/B[3] ) );
  XNOR2_X1 U4462 ( .A(n820), .B(n819), .ZN(\intadd_2/A[2] ) );
  NOR2_X1 U4463 ( .A1(n941), .A2(n1083), .ZN(n823) );
  INV_X1 U4464 ( .A(s_A_MULT[8]), .ZN(n821) );
  OAI22_X1 U4465 ( .A1(n821), .A2(n945), .B1(n936), .B2(n981), .ZN(n822) );
  AOI211_X1 U4466 ( .C1(n948), .C2(s_A_MULT[9]), .A(n823), .B(n822), .ZN(
        \intadd_2/B[0] ) );
  OAI21_X1 U4467 ( .B1(n824), .B2(n840), .A(n841), .ZN(n1243) );
  INV_X1 U4468 ( .A(n1243), .ZN(n1036) );
  AOI222_X1 U4469 ( .A1(s_A_MULT[11]), .A2(n1309), .B1(n1308), .B2(n1036), 
        .C1(n55), .C2(n1171), .ZN(\intadd_2/CI ) );
  AOI22_X1 U4470 ( .A1(s_A_MULT[9]), .A2(n968), .B1(n967), .B2(n1171), .ZN(
        n825) );
  OAI21_X1 U4471 ( .B1(n1056), .B2(n1083), .A(n825), .ZN(n826) );
  AOI21_X1 U4472 ( .B1(s_A_MULT[10]), .B2(n966), .A(n826), .ZN(\intadd_3/A[0] ) );
  AOI22_X1 U4473 ( .A1(s_A_MULT[3]), .A2(n1259), .B1(n1258), .B2(n959), .ZN(
        n827) );
  OAI21_X1 U4474 ( .B1(n1231), .B2(n934), .A(n827), .ZN(n828) );
  AOI21_X1 U4475 ( .B1(s_A_MULT[4]), .B2(n1262), .A(n828), .ZN(n849) );
  AOI22_X1 U4476 ( .A1(n1070), .A2(s_A_MULT[7]), .B1(n1089), .B2(n56), .ZN(
        n829) );
  OAI21_X1 U4477 ( .B1(n1041), .B2(n1087), .A(n829), .ZN(n830) );
  AOI21_X1 U4478 ( .B1(n1073), .B2(s_A_MULT[6]), .A(n830), .ZN(n846) );
  AOI22_X1 U4479 ( .A1(s_A_MULT[4]), .A2(n1160), .B1(n1159), .B2(n831), .ZN(
        n832) );
  OAI21_X1 U4480 ( .B1(n833), .B2(n1252), .A(n832), .ZN(n834) );
  AOI21_X1 U4481 ( .B1(s_A_MULT[5]), .B2(n1085), .A(n834), .ZN(n845) );
  AOI22_X1 U4482 ( .A1(s_A_MULT[9]), .A2(n1048), .B1(s_A_MULT[8]), .B2(n1076), 
        .ZN(n835) );
  OAI21_X1 U4483 ( .B1(n1046), .B2(n1083), .A(n835), .ZN(n836) );
  AOI21_X1 U4484 ( .B1(n1075), .B2(n1068), .A(n836), .ZN(n844) );
  AOI22_X1 U4485 ( .A1(s_A_MULT[1]), .A2(n1246), .B1(n1239), .B2(n908), .ZN(
        n837) );
  OAI21_X1 U4486 ( .B1(n1242), .B2(n838), .A(n837), .ZN(n839) );
  AOI21_X1 U4487 ( .B1(s_A_MULT[2]), .B2(n1247), .A(n839), .ZN(n847) );
  NOR2_X1 U4488 ( .A1(n840), .A2(n945), .ZN(n843) );
  AOI21_X1 U4489 ( .B1(s_A_MULT[12]), .B2(n841), .A(n853), .ZN(n1244) );
  INV_X1 U4490 ( .A(n1244), .ZN(n996) );
  OAI22_X1 U4491 ( .A1(n941), .A2(n996), .B1(n936), .B2(n1243), .ZN(n842) );
  AOI211_X1 U4492 ( .C1(n948), .C2(s_A_MULT[12]), .A(n843), .B(n842), .ZN(
        \intadd_3/B[0] ) );
  FA_X1 U4493 ( .A(n846), .B(n845), .CI(n844), .CO(n848), .S(\intadd_3/B[1] )
         );
  FA_X1 U4494 ( .A(n849), .B(n848), .CI(n847), .CO(\intadd_3/B[3] ), .S(
        \intadd_3/A[2] ) );
  AND2_X1 U4495 ( .A1(S_B_MULT[1]), .A2(S_B_MULT[0]), .ZN(n854) );
  OAI21_X1 U4496 ( .B1(n851), .B2(n1079), .A(n850), .ZN(n1232) );
  INV_X1 U4497 ( .A(n1232), .ZN(n1261) );
  OAI21_X1 U4498 ( .B1(n853), .B2(n1236), .A(n852), .ZN(n1250) );
  INV_X1 U4499 ( .A(n1250), .ZN(n1074) );
  AOI222_X1 U4500 ( .A1(s_A_MULT[14]), .A2(n1309), .B1(n854), .B2(n1261), .C1(
        n55), .C2(n1074), .ZN(\intadd_3/CI ) );
  NOR2_X1 U4501 ( .A1(S_B_MULT[0]), .A2(n942), .ZN(n858) );
  OAI22_X1 U4502 ( .A1(n1253), .A2(n856), .B1(n1164), .B2(n855), .ZN(n857) );
  AOI21_X1 U4503 ( .B1(n1261), .B2(n858), .A(n857), .ZN(\intadd_4/A[0] ) );
  AOI22_X1 U4504 ( .A1(n1073), .A2(s_A_MULT[7]), .B1(n1069), .B2(n1068), .ZN(
        n859) );
  OAI21_X1 U4505 ( .B1(n53), .B2(n1087), .A(n859), .ZN(n860) );
  AOI21_X1 U4506 ( .B1(n1070), .B2(s_A_MULT[8]), .A(n860), .ZN(n871) );
  AOI22_X1 U4507 ( .A1(s_A_MULT[5]), .A2(n1160), .B1(n1159), .B2(n1089), .ZN(
        n861) );
  OAI21_X1 U4508 ( .B1(n988), .B2(n1252), .A(n861), .ZN(n862) );
  AOI21_X1 U4509 ( .B1(s_A_MULT[6]), .B2(n1085), .A(n862), .ZN(n870) );
  INV_X1 U4510 ( .A(n1171), .ZN(n1038) );
  AOI22_X1 U4511 ( .A1(s_A_MULT[9]), .A2(n1076), .B1(n1075), .B2(n979), .ZN(
        n863) );
  OAI21_X1 U4512 ( .B1(n1046), .B2(n1038), .A(n863), .ZN(n864) );
  AOI21_X1 U4513 ( .B1(s_A_MULT[10]), .B2(n1048), .A(n864), .ZN(n869) );
  AOI22_X1 U4514 ( .A1(s_A_MULT[2]), .A2(n1246), .B1(n1239), .B2(n899), .ZN(
        n865) );
  OAI21_X1 U4515 ( .B1(n1242), .B2(n902), .A(n865), .ZN(n866) );
  AOI21_X1 U4516 ( .B1(s_A_MULT[3]), .B2(n1247), .A(n866), .ZN(n877) );
  AOI22_X1 U4517 ( .A1(s_A_MULT[5]), .A2(n1262), .B1(s_A_MULT[4]), .B2(n1259), 
        .ZN(n867) );
  OAI21_X1 U4518 ( .B1(n63), .B2(n988), .A(n867), .ZN(n868) );
  AOI21_X1 U4519 ( .B1(n1260), .B2(n959), .A(n868), .ZN(n876) );
  FA_X1 U4520 ( .A(n871), .B(n870), .CI(n869), .CO(n875), .S(\intadd_4/A[1] )
         );
  INV_X1 U4521 ( .A(s_A_MULT[12]), .ZN(n872) );
  NOR2_X1 U4522 ( .A1(n872), .A2(n945), .ZN(n874) );
  OAI22_X1 U4523 ( .A1(n941), .A2(n1250), .B1(n936), .B2(n996), .ZN(n873) );
  AOI211_X1 U4524 ( .C1(n948), .C2(s_A_MULT[13]), .A(n874), .B(n873), .ZN(
        \intadd_4/B[0] ) );
  FA_X1 U4525 ( .A(n877), .B(n876), .CI(n875), .CO(\intadd_4/B[3] ), .S(
        \intadd_4/A[2] ) );
  AOI22_X1 U4526 ( .A1(s_A_MULT[10]), .A2(n968), .B1(n967), .B2(n1036), .ZN(
        n878) );
  OAI21_X1 U4527 ( .B1(n1056), .B2(n1038), .A(n878), .ZN(n879) );
  AOI21_X1 U4528 ( .B1(s_A_MULT[11]), .B2(n966), .A(n879), .ZN(\intadd_4/CI )
         );
  AOI222_X1 U4529 ( .A1(s_A_MULT[13]), .A2(n1309), .B1(n1308), .B2(n1074), 
        .C1(n55), .C2(n1244), .ZN(\intadd_5/A[0] ) );
  AOI22_X1 U4530 ( .A1(s_A_MULT[3]), .A2(n1262), .B1(s_A_MULT[2]), .B2(n1259), 
        .ZN(n880) );
  OAI21_X1 U4531 ( .B1(n63), .B2(n934), .A(n880), .ZN(n881) );
  AOI21_X1 U4532 ( .B1(n1260), .B2(n908), .A(n881), .ZN(n1328) );
  INV_X1 U4533 ( .A(n1242), .ZN(n1245) );
  OR2_X1 U4534 ( .A1(n1245), .A2(n1246), .ZN(n882) );
  AOI222_X1 U4535 ( .A1(n882), .A2(\MULT/SHIFTERi_0/N19 ), .B1(n1239), .B2(
        n1307), .C1(s_A_MULT[1]), .C2(n1247), .ZN(n1327) );
  AOI22_X1 U4536 ( .A1(n1070), .A2(s_A_MULT[6]), .B1(n1073), .B2(s_A_MULT[5]), 
        .ZN(n883) );
  OAI21_X1 U4537 ( .B1(n988), .B2(n53), .A(n883), .ZN(n884) );
  AOI21_X1 U4538 ( .B1(n1069), .B2(n1089), .A(n884), .ZN(n894) );
  AOI22_X1 U4539 ( .A1(s_A_MULT[3]), .A2(n1160), .B1(n1159), .B2(n959), .ZN(
        n885) );
  OAI21_X1 U4540 ( .B1(n934), .B2(n1252), .A(n885), .ZN(n886) );
  AOI21_X1 U4541 ( .B1(s_A_MULT[4]), .B2(n1085), .A(n886), .ZN(n893) );
  AOI22_X1 U4542 ( .A1(s_A_MULT[8]), .A2(n1048), .B1(n1075), .B2(n920), .ZN(
        n887) );
  OAI21_X1 U4543 ( .B1(n1046), .B2(n981), .A(n887), .ZN(n888) );
  AOI21_X1 U4544 ( .B1(s_A_MULT[7]), .B2(n1076), .A(n888), .ZN(n892) );
  INV_X1 U4545 ( .A(s_A_MULT[10]), .ZN(n889) );
  NOR2_X1 U4546 ( .A1(n889), .A2(n945), .ZN(n891) );
  OAI22_X1 U4547 ( .A1(n941), .A2(n1243), .B1(n936), .B2(n1038), .ZN(n890) );
  AOI211_X1 U4548 ( .C1(n948), .C2(s_A_MULT[11]), .A(n891), .B(n890), .ZN(
        \intadd_5/B[0] ) );
  FA_X1 U4549 ( .A(n894), .B(n893), .CI(n892), .CO(n1326), .S(\intadd_5/B[1] )
         );
  AOI22_X1 U4550 ( .A1(s_A_MULT[8]), .A2(n968), .B1(n967), .B2(n979), .ZN(n895) );
  OAI21_X1 U4551 ( .B1(n1056), .B2(n981), .A(n895), .ZN(n896) );
  AOI21_X1 U4552 ( .B1(s_A_MULT[9]), .B2(n966), .A(n896), .ZN(\intadd_5/CI )
         );
  AOI22_X1 U4553 ( .A1(s_A_MULT[8]), .A2(n966), .B1(n967), .B2(n1068), .ZN(
        n897) );
  OAI21_X1 U4554 ( .B1(n1056), .B2(n1087), .A(n897), .ZN(n898) );
  AOI21_X1 U4555 ( .B1(s_A_MULT[7]), .B2(n968), .A(n898), .ZN(\intadd_6/A[0] )
         );
  AOI22_X1 U4556 ( .A1(s_A_MULT[3]), .A2(n1085), .B1(n1159), .B2(n899), .ZN(
        n901) );
  OAI21_X1 U4557 ( .B1(n902), .B2(n1252), .A(n901), .ZN(n903) );
  AOI21_X1 U4558 ( .B1(s_A_MULT[2]), .B2(n1160), .A(n903), .ZN(n914) );
  AOI22_X1 U4559 ( .A1(n1070), .A2(s_A_MULT[5]), .B1(n1073), .B2(s_A_MULT[4]), 
        .ZN(n904) );
  OAI21_X1 U4560 ( .B1(n1041), .B2(n988), .A(n904), .ZN(n905) );
  AOI21_X1 U4561 ( .B1(n959), .B2(n56), .A(n905), .ZN(n913) );
  AOI22_X1 U4562 ( .A1(s_A_MULT[7]), .A2(n1048), .B1(s_A_MULT[6]), .B2(n1076), 
        .ZN(n906) );
  OAI21_X1 U4563 ( .B1(n1046), .B2(n1087), .A(n906), .ZN(n907) );
  AOI21_X1 U4564 ( .B1(n1089), .B2(n1075), .A(n907), .ZN(n912) );
  AOI22_X1 U4565 ( .A1(s_A_MULT[2]), .A2(n1262), .B1(n1258), .B2(n908), .ZN(
        n909) );
  OAI21_X1 U4566 ( .B1(n910), .B2(n1235), .A(n909), .ZN(n911) );
  AOI21_X1 U4567 ( .B1(n1260), .B2(n1307), .A(n911), .ZN(n1132) );
  OAI21_X1 U4568 ( .B1(n1247), .B2(n1239), .A(\MULT/SHIFTERi_0/N19 ), .ZN(
        n1131) );
  FA_X1 U4569 ( .A(n914), .B(n913), .CI(n912), .CO(n1130), .S(\intadd_6/A[1] )
         );
  AOI222_X1 U4570 ( .A1(s_A_MULT[12]), .A2(n1309), .B1(n1308), .B2(n1244), 
        .C1(n55), .C2(n1036), .ZN(\intadd_6/B[0] ) );
  NOR2_X1 U4571 ( .A1(n941), .A2(n1038), .ZN(n917) );
  OAI22_X1 U4572 ( .A1(n915), .A2(n945), .B1(n936), .B2(n1083), .ZN(n916) );
  AOI211_X1 U4573 ( .C1(n948), .C2(s_A_MULT[10]), .A(n917), .B(n916), .ZN(
        \intadd_6/CI ) );
  AOI22_X1 U4574 ( .A1(s_A_MULT[11]), .A2(n968), .B1(n967), .B2(n1244), .ZN(
        n918) );
  OAI21_X1 U4575 ( .B1(n1056), .B2(n1243), .A(n918), .ZN(n919) );
  AOI21_X1 U4576 ( .B1(s_A_MULT[12]), .B2(n966), .A(n919), .ZN(\intadd_7/A[0] ) );
  AOI22_X1 U4577 ( .A1(s_A_MULT[7]), .A2(n1085), .B1(n1159), .B2(n920), .ZN(
        n921) );
  OAI21_X1 U4578 ( .B1(n922), .B2(n1252), .A(n921), .ZN(n923) );
  AOI21_X1 U4579 ( .B1(s_A_MULT[6]), .B2(n1160), .A(n923), .ZN(n932) );
  AOI22_X1 U4580 ( .A1(n1070), .A2(s_A_MULT[9]), .B1(n56), .B2(n1068), .ZN(
        n924) );
  OAI21_X1 U4581 ( .B1(n1041), .B2(n1083), .A(n924), .ZN(n925) );
  AOI21_X1 U4582 ( .B1(n1073), .B2(s_A_MULT[8]), .A(n925), .ZN(n931) );
  AOI22_X1 U4583 ( .A1(s_A_MULT[11]), .A2(n1048), .B1(n1075), .B2(n1171), .ZN(
        n926) );
  OAI21_X1 U4584 ( .B1(n1046), .B2(n1243), .A(n926), .ZN(n927) );
  AOI21_X1 U4585 ( .B1(s_A_MULT[10]), .B2(n1076), .A(n927), .ZN(n930) );
  AOI22_X1 U4586 ( .A1(s_A_MULT[5]), .A2(n1259), .B1(n1258), .B2(n1089), .ZN(
        n928) );
  OAI21_X1 U4587 ( .B1(n988), .B2(n1231), .A(n928), .ZN(n929) );
  AOI21_X1 U4588 ( .B1(s_A_MULT[6]), .B2(n1262), .A(n929), .ZN(n1117) );
  FA_X1 U4589 ( .A(n932), .B(n931), .CI(n930), .CO(n1118), .S(\intadd_7/A[1] )
         );
  AOI22_X1 U4590 ( .A1(s_A_MULT[3]), .A2(n1246), .B1(n1239), .B2(n959), .ZN(
        n933) );
  OAI21_X1 U4591 ( .B1(n1242), .B2(n934), .A(n933), .ZN(n935) );
  AOI21_X1 U4592 ( .B1(s_A_MULT[4]), .B2(n1247), .A(n935), .ZN(n1116) );
  INV_X1 U4593 ( .A(n936), .ZN(n994) );
  AOI22_X1 U4594 ( .A1(s_A_MULT[14]), .A2(n948), .B1(n994), .B2(n1074), .ZN(
        n937) );
  OAI21_X1 U4595 ( .B1(n1236), .B2(n945), .A(n937), .ZN(n938) );
  AOI21_X1 U4596 ( .B1(n939), .B2(n1261), .A(n938), .ZN(\intadd_7/B[0] ) );
  AOI21_X1 U4597 ( .B1(n55), .B2(n1257), .A(n940), .ZN(\intadd_7/CI ) );
  NOR2_X1 U4598 ( .A1(n1253), .A2(n941), .ZN(n947) );
  NAND2_X1 U4599 ( .A1(n943), .A2(n942), .ZN(n944) );
  OAI22_X1 U4600 ( .A1(n1079), .A2(n945), .B1(n1232), .B2(n944), .ZN(n946) );
  AOI211_X1 U4601 ( .C1(n948), .C2(s_A_MULT[15]), .A(n947), .B(n946), .ZN(
        \intadd_8/A[0] ) );
  AOI22_X1 U4602 ( .A1(n1070), .A2(s_A_MULT[10]), .B1(n1069), .B2(n1171), .ZN(
        n949) );
  OAI21_X1 U4603 ( .B1(n53), .B2(n1083), .A(n949), .ZN(n950) );
  AOI21_X1 U4604 ( .B1(n1073), .B2(s_A_MULT[9]), .A(n950), .ZN(n962) );
  AOI22_X1 U4605 ( .A1(s_A_MULT[12]), .A2(n1048), .B1(n1075), .B2(n1036), .ZN(
        n951) );
  OAI21_X1 U4606 ( .B1(n1046), .B2(n996), .A(n951), .ZN(n952) );
  AOI21_X1 U4607 ( .B1(s_A_MULT[11]), .B2(n1076), .A(n952), .ZN(n961) );
  AOI22_X1 U4608 ( .A1(s_A_MULT[8]), .A2(n1085), .B1(n1159), .B2(n1068), .ZN(
        n953) );
  OAI21_X1 U4609 ( .B1(n1252), .B2(n1087), .A(n953), .ZN(n954) );
  AOI21_X1 U4610 ( .B1(s_A_MULT[7]), .B2(n1160), .A(n954), .ZN(n960) );
  AOI22_X1 U4611 ( .A1(s_A_MULT[6]), .A2(n1259), .B1(n1260), .B2(n1089), .ZN(
        n955) );
  OAI21_X1 U4612 ( .B1(n63), .B2(n1087), .A(n955), .ZN(n956) );
  AOI21_X1 U4613 ( .B1(s_A_MULT[7]), .B2(n1262), .A(n956), .ZN(n1112) );
  AOI22_X1 U4614 ( .A1(s_A_MULT[5]), .A2(n1247), .B1(s_A_MULT[4]), .B2(n1246), 
        .ZN(n957) );
  OAI21_X1 U4615 ( .B1(n61), .B2(n988), .A(n957), .ZN(n958) );
  AOI21_X1 U4616 ( .B1(n1245), .B2(n959), .A(n958), .ZN(n1111) );
  FA_X1 U4617 ( .A(n962), .B(n961), .CI(n960), .CO(n1110), .S(\intadd_8/B[1] )
         );
  AOI22_X1 U4618 ( .A1(s_A_MULT[12]), .A2(n968), .B1(n967), .B2(n1074), .ZN(
        n963) );
  OAI21_X1 U4619 ( .B1(n1056), .B2(n996), .A(n963), .ZN(n964) );
  AOI21_X1 U4620 ( .B1(s_A_MULT[13]), .B2(n966), .A(n964), .ZN(\intadd_8/CI )
         );
  INV_X1 U4621 ( .A(n1103), .ZN(n965) );
  NOR2_X1 U4622 ( .A1(n1101), .A2(n965), .ZN(n1100) );
  INV_X1 U4623 ( .A(n966), .ZN(n974) );
  AOI22_X1 U4624 ( .A1(s_A_MULT[14]), .A2(n968), .B1(n967), .B2(n1257), .ZN(
        n971) );
  NAND3_X1 U4625 ( .A1(S_B_MULT[5]), .A2(n969), .A3(n1261), .ZN(n970) );
  OAI211_X1 U4626 ( .C1(n974), .C2(n1164), .A(n971), .B(n970), .ZN(n1102) );
  XNOR2_X1 U4627 ( .A(n1100), .B(n1102), .ZN(\intadd_9/A[1] ) );
  OAI22_X1 U4628 ( .A1(n972), .A2(n1232), .B1(n1056), .B2(n1250), .ZN(n976) );
  OAI22_X1 U4629 ( .A1(n1079), .A2(n974), .B1(n1236), .B2(n973), .ZN(n975) );
  NOR2_X1 U4630 ( .A1(n976), .A2(n975), .ZN(\intadd_9/B[0] ) );
  AOI22_X1 U4631 ( .A1(n1070), .A2(s_A_MULT[11]), .B1(n56), .B2(n1171), .ZN(
        n977) );
  OAI21_X1 U4632 ( .B1(n1041), .B2(n1243), .A(n977), .ZN(n978) );
  AOI21_X1 U4633 ( .B1(n1073), .B2(s_A_MULT[10]), .A(n978), .ZN(n992) );
  AOI22_X1 U4634 ( .A1(s_A_MULT[8]), .A2(n1160), .B1(n1159), .B2(n979), .ZN(
        n980) );
  OAI21_X1 U4635 ( .B1(n1252), .B2(n981), .A(n980), .ZN(n982) );
  AOI21_X1 U4636 ( .B1(s_A_MULT[9]), .B2(n1085), .A(n982), .ZN(n991) );
  AOI22_X1 U4637 ( .A1(s_A_MULT[13]), .A2(n1048), .B1(n1075), .B2(n1244), .ZN(
        n983) );
  OAI21_X1 U4638 ( .B1(n1046), .B2(n1250), .A(n983), .ZN(n984) );
  AOI21_X1 U4639 ( .B1(s_A_MULT[12]), .B2(n1076), .A(n984), .ZN(n990) );
  AOI22_X1 U4640 ( .A1(s_A_MULT[7]), .A2(n1259), .B1(n1068), .B2(n1258), .ZN(
        n985) );
  OAI21_X1 U4641 ( .B1(n1231), .B2(n1087), .A(n985), .ZN(n986) );
  AOI21_X1 U4642 ( .B1(s_A_MULT[8]), .B2(n1262), .A(n986), .ZN(n1144) );
  AOI22_X1 U4643 ( .A1(s_A_MULT[5]), .A2(n1246), .B1(n1239), .B2(n1089), .ZN(
        n987) );
  OAI21_X1 U4644 ( .B1(n1242), .B2(n988), .A(n987), .ZN(n989) );
  AOI21_X1 U4645 ( .B1(s_A_MULT[6]), .B2(n1247), .A(n989), .ZN(n1143) );
  FA_X1 U4646 ( .A(n992), .B(n991), .CI(n990), .CO(n1142), .S(\intadd_9/B[1] )
         );
  AOI21_X1 U4647 ( .B1(n994), .B2(n1257), .A(n993), .ZN(\intadd_9/CI ) );
  AOI22_X1 U4648 ( .A1(s_A_MULT[13]), .A2(n1085), .B1(n1159), .B2(n1074), .ZN(
        n995) );
  OAI21_X1 U4649 ( .B1(n1252), .B2(n996), .A(n995), .ZN(n997) );
  AOI21_X1 U4650 ( .B1(s_A_MULT[12]), .B2(n1160), .A(n997), .ZN(n1007) );
  AOI22_X1 U4651 ( .A1(n1073), .A2(s_A_MULT[14]), .B1(n1069), .B2(n1257), .ZN(
        n998) );
  OAI21_X1 U4652 ( .B1(n1164), .B2(n999), .A(n998), .ZN(n1000) );
  AOI21_X1 U4653 ( .B1(n1261), .B2(n56), .A(n1000), .ZN(n1006) );
  OAI21_X1 U4654 ( .B1(n1269), .B2(n1013), .A(n1267), .ZN(n1183) );
  INV_X1 U4655 ( .A(n1267), .ZN(n1270) );
  NOR2_X1 U4656 ( .A1(n1270), .A2(n1269), .ZN(n1273) );
  OAI22_X1 U4657 ( .A1(n1079), .A2(n1165), .B1(n1252), .B2(n1250), .ZN(n1004)
         );
  OAI22_X1 U4658 ( .A1(n1236), .A2(n1002), .B1(n1001), .B2(n1232), .ZN(n1003)
         );
  NOR2_X1 U4659 ( .A1(n1004), .A2(n1003), .ZN(n1169) );
  AOI21_X1 U4660 ( .B1(n56), .B2(n1257), .A(n1005), .ZN(n1168) );
  XNOR2_X1 U4661 ( .A(n1273), .B(n1166), .ZN(n1182) );
  FA_X1 U4662 ( .A(n1170), .B(n1007), .CI(n1006), .CO(n1179), .S(n1013) );
  AOI22_X1 U4663 ( .A1(s_A_MULT[11]), .A2(n1259), .B1(n1258), .B2(n1244), .ZN(
        n1008) );
  OAI21_X1 U4664 ( .B1(n1231), .B2(n1243), .A(n1008), .ZN(n1009) );
  AOI21_X1 U4665 ( .B1(s_A_MULT[12]), .B2(n1262), .A(n1009), .ZN(n1178) );
  AOI22_X1 U4666 ( .A1(s_A_MULT[9]), .A2(n1246), .B1(n1239), .B2(n1171), .ZN(
        n1010) );
  OAI21_X1 U4667 ( .B1(n1242), .B2(n1083), .A(n1010), .ZN(n1011) );
  AOI21_X1 U4668 ( .B1(s_A_MULT[10]), .B2(n1247), .A(n1011), .ZN(n1177) );
  INV_X1 U4669 ( .A(n1012), .ZN(n1181) );
  XNOR2_X1 U4670 ( .A(n1273), .B(n1013), .ZN(n1035) );
  AOI21_X1 U4671 ( .B1(n1075), .B2(n1257), .A(n1014), .ZN(n1025) );
  AOI22_X1 U4672 ( .A1(n1070), .A2(s_A_MULT[14]), .B1(n1069), .B2(n1261), .ZN(
        n1015) );
  OAI21_X1 U4673 ( .B1(n53), .B2(n1250), .A(n1015), .ZN(n1016) );
  AOI21_X1 U4674 ( .B1(n1073), .B2(s_A_MULT[13]), .A(n1016), .ZN(n1024) );
  AOI22_X1 U4675 ( .A1(s_A_MULT[11]), .A2(n1160), .B1(n1159), .B2(n1244), .ZN(
        n1017) );
  OAI21_X1 U4676 ( .B1(n1252), .B2(n1243), .A(n1017), .ZN(n1018) );
  AOI21_X1 U4677 ( .B1(s_A_MULT[12]), .B2(n1085), .A(n1018), .ZN(n1023) );
  OAI21_X1 U4678 ( .B1(n1269), .B2(n1053), .A(n1267), .ZN(n1034) );
  AOI22_X1 U4679 ( .A1(s_A_MULT[10]), .A2(n1259), .B1(n1260), .B2(n1171), .ZN(
        n1019) );
  OAI21_X1 U4680 ( .B1(n63), .B2(n1243), .A(n1019), .ZN(n1020) );
  AOI21_X1 U4681 ( .B1(s_A_MULT[11]), .B2(n1262), .A(n1020), .ZN(n1029) );
  AOI22_X1 U4682 ( .A1(s_A_MULT[9]), .A2(n1247), .B1(s_A_MULT[8]), .B2(n1246), 
        .ZN(n1021) );
  OAI21_X1 U4683 ( .B1(n61), .B2(n1083), .A(n1021), .ZN(n1022) );
  AOI21_X1 U4684 ( .B1(n1245), .B2(n1068), .A(n1022), .ZN(n1028) );
  FA_X1 U4685 ( .A(n1025), .B(n1024), .CI(n1023), .CO(n1027), .S(n1053) );
  INV_X1 U4686 ( .A(n1026), .ZN(n1033) );
  FA_X1 U4687 ( .A(n1029), .B(n1028), .CI(n1027), .CO(n1030), .S(n1026) );
  INV_X1 U4688 ( .A(n1030), .ZN(n1337) );
  AOI22_X1 U4689 ( .A1(n72), .A2(n1031), .B1(A[24]), .B2(n1374), .ZN(n1032) );
  INV_X1 U4690 ( .A(n1032), .ZN(n105) );
  INV_X1 U4691 ( .A(A[23]), .ZN(n1065) );
  FA_X1 U4692 ( .A(n1035), .B(n1034), .CI(n1033), .CO(n1338), .S(n1355) );
  AOI22_X1 U4693 ( .A1(s_A_MULT[11]), .A2(n1085), .B1(n1159), .B2(n1036), .ZN(
        n1037) );
  OAI21_X1 U4694 ( .B1(n1252), .B2(n1038), .A(n1037), .ZN(n1039) );
  AOI21_X1 U4695 ( .B1(s_A_MULT[10]), .B2(n1160), .A(n1039), .ZN(n1059) );
  AOI22_X1 U4696 ( .A1(n1070), .A2(s_A_MULT[13]), .B1(n56), .B2(n1244), .ZN(
        n1040) );
  OAI21_X1 U4697 ( .B1(n1041), .B2(n1250), .A(n1040), .ZN(n1042) );
  AOI21_X1 U4698 ( .B1(n1073), .B2(s_A_MULT[12]), .A(n1042), .ZN(n1058) );
  NOR3_X1 U4699 ( .A1(S_B_MULT[6]), .A2(S_B_MULT[5]), .A3(n1043), .ZN(n1044)
         );
  AOI22_X1 U4700 ( .A1(s_A_MULT[14]), .A2(n1076), .B1(n1261), .B2(n1044), .ZN(
        n1045) );
  OAI21_X1 U4701 ( .B1(n1253), .B2(n1046), .A(n1045), .ZN(n1047) );
  AOI21_X1 U4702 ( .B1(s_A_MULT[15]), .B2(n1048), .A(n1047), .ZN(n1057) );
  AOI22_X1 U4703 ( .A1(s_A_MULT[7]), .A2(n1246), .B1(n1239), .B2(n1068), .ZN(
        n1049) );
  OAI21_X1 U4704 ( .B1(n1242), .B2(n1087), .A(n1049), .ZN(n1050) );
  AOI21_X1 U4705 ( .B1(s_A_MULT[8]), .B2(n1247), .A(n1050), .ZN(n1061) );
  AOI22_X1 U4706 ( .A1(s_A_MULT[9]), .A2(n1259), .B1(n1258), .B2(n1171), .ZN(
        n1051) );
  OAI21_X1 U4707 ( .B1(n1231), .B2(n1083), .A(n1051), .ZN(n1052) );
  AOI21_X1 U4708 ( .B1(s_A_MULT[10]), .B2(n1262), .A(n1052), .ZN(n1060) );
  XOR2_X1 U4709 ( .A(n1273), .B(n1053), .Z(n1092) );
  XNOR2_X1 U4710 ( .A(n1100), .B(n1054), .ZN(n1095) );
  OAI21_X1 U4711 ( .B1(n1253), .B2(n1056), .A(n1055), .ZN(n1099) );
  AOI21_X1 U4712 ( .B1(n1103), .B2(n1099), .A(n1101), .ZN(n1094) );
  FA_X1 U4713 ( .A(n1059), .B(n1058), .CI(n1057), .CO(n1062), .S(n1093) );
  FA_X1 U4714 ( .A(n1062), .B(n1061), .CI(n1060), .CO(n1351), .S(n1090) );
  NOR2_X1 U4715 ( .A1(n1352), .A2(n1351), .ZN(n1353) );
  AOI21_X1 U4716 ( .B1(n1351), .B2(n1352), .A(n1353), .ZN(n1063) );
  XNOR2_X1 U4717 ( .A(n1355), .B(n1063), .ZN(n1064) );
  OAI22_X1 U4718 ( .A1(n1396), .A2(n1065), .B1(n73), .B2(n1064), .ZN(n107) );
  INV_X1 U4719 ( .A(A[22]), .ZN(n1109) );
  AOI22_X1 U4720 ( .A1(s_A_MULT[9]), .A2(n1262), .B1(s_A_MULT[8]), .B2(n1259), 
        .ZN(n1066) );
  OAI21_X1 U4721 ( .B1(n63), .B2(n1083), .A(n1066), .ZN(n1067) );
  AOI21_X1 U4722 ( .B1(n1260), .B2(n1068), .A(n1067), .ZN(n1098) );
  AOI22_X1 U4723 ( .A1(n1070), .A2(s_A_MULT[12]), .B1(n1069), .B2(n1244), .ZN(
        n1071) );
  OAI21_X1 U4724 ( .B1(n53), .B2(n1243), .A(n1071), .ZN(n1072) );
  AOI21_X1 U4725 ( .B1(n1073), .B2(s_A_MULT[11]), .A(n1072), .ZN(n1106) );
  AOI22_X1 U4726 ( .A1(s_A_MULT[13]), .A2(n1076), .B1(n1075), .B2(n1074), .ZN(
        n1077) );
  OAI21_X1 U4727 ( .B1(n1079), .B2(n1078), .A(n1077), .ZN(n1080) );
  AOI21_X1 U4728 ( .B1(n1081), .B2(n1261), .A(n1080), .ZN(n1105) );
  AOI22_X1 U4729 ( .A1(s_A_MULT[9]), .A2(n1160), .B1(n1159), .B2(n1171), .ZN(
        n1082) );
  OAI21_X1 U4730 ( .B1(n1252), .B2(n1083), .A(n1082), .ZN(n1084) );
  AOI21_X1 U4731 ( .B1(s_A_MULT[10]), .B2(n1085), .A(n1084), .ZN(n1104) );
  AOI22_X1 U4732 ( .A1(s_A_MULT[7]), .A2(n1247), .B1(s_A_MULT[6]), .B2(n1246), 
        .ZN(n1086) );
  OAI21_X1 U4733 ( .B1(n61), .B2(n1087), .A(n1086), .ZN(n1088) );
  AOI21_X1 U4734 ( .B1(n1245), .B2(n1089), .A(n1088), .ZN(n1096) );
  FA_X1 U4735 ( .A(n1092), .B(n1091), .CI(n1090), .CO(n1352), .S(n1347) );
  XNOR2_X1 U4736 ( .A(n1348), .B(n1347), .ZN(n1107) );
  FA_X1 U4737 ( .A(n1095), .B(n1094), .CI(n1093), .CO(n1091), .S(n1141) );
  FA_X1 U4738 ( .A(n1098), .B(n1097), .CI(n1096), .CO(n1348), .S(n1140) );
  XNOR2_X1 U4739 ( .A(n1100), .B(n1099), .ZN(n1306) );
  AOI21_X1 U4740 ( .B1(n1103), .B2(n1102), .A(n1101), .ZN(n1305) );
  FA_X1 U4741 ( .A(n1106), .B(n1105), .CI(n1104), .CO(n1097), .S(n1304) );
  XNOR2_X1 U4742 ( .A(n1107), .B(n1346), .ZN(n1108) );
  OAI22_X1 U4743 ( .A1(n1396), .A2(n1109), .B1(n1108), .B2(n74), .ZN(n110) );
  FA_X1 U4744 ( .A(n1112), .B(n1111), .CI(n1110), .CO(n1334), .S(
        \intadd_8/B[2] ) );
  NOR2_X1 U4745 ( .A1(n1113), .A2(n74), .ZN(n1114) );
  AOI21_X1 U4746 ( .B1(A[20]), .B2(n1374), .A(n1114), .ZN(n1119) );
  FA_X1 U4747 ( .A(n1117), .B(n1118), .CI(n1116), .CO(n1122), .S(
        \intadd_7/A[2] ) );
  AND2_X1 U4748 ( .A1(n1118), .A2(n1117), .ZN(n1115) );
  OAI221_X1 U4749 ( .B1(n1118), .B2(n1117), .C1(n1116), .C2(n1115), .A(
        \intadd_7/n1 ), .ZN(n1124) );
  OAI21_X1 U4750 ( .B1(\intadd_7/n1 ), .B2(n1122), .A(n1124), .ZN(n1120) );
  XOR2_X1 U4751 ( .A(\intadd_8/SUM[2] ), .B(n1120), .Z(n1121) );
  AOI22_X1 U4752 ( .A1(n72), .A2(n1121), .B1(A[19]), .B2(n1374), .ZN(n1155) );
  INV_X1 U4753 ( .A(B[20]), .ZN(n1127) );
  INV_X1 U4754 ( .A(\intadd_8/SUM[2] ), .ZN(n1125) );
  NOR2_X1 U4755 ( .A1(\intadd_7/n1 ), .A2(n1122), .ZN(n1123) );
  AOI21_X1 U4756 ( .B1(n1125), .B2(n1124), .A(n1123), .ZN(n1126) );
  OAI22_X1 U4757 ( .A1(n1396), .A2(n1127), .B1(n1126), .B2(n74), .ZN(n118) );
  INV_X1 U4758 ( .A(A[18]), .ZN(n1128) );
  OAI22_X1 U4759 ( .A1(n1396), .A2(n1128), .B1(\intadd_4/SUM[3] ), .B2(n74), 
        .ZN(n119) );
  INV_X1 U4760 ( .A(A[17]), .ZN(n1129) );
  OAI22_X1 U4761 ( .A1(n1396), .A2(n1129), .B1(\intadd_3/SUM[3] ), .B2(n73), 
        .ZN(n122) );
  INV_X1 U4762 ( .A(A[15]), .ZN(n1134) );
  FA_X1 U4763 ( .A(n1132), .B(n1131), .CI(n1130), .CO(n1323), .S(
        \intadd_6/A[2] ) );
  OAI22_X1 U4764 ( .A1(n70), .A2(n1134), .B1(n1133), .B2(n74), .ZN(n127) );
  NOR3_X1 U4765 ( .A1(n1452), .A2(n1451), .A3(n1135), .ZN(n1619) );
  INV_X1 U4766 ( .A(B[19]), .ZN(n1137) );
  OAI22_X1 U4767 ( .A1(n1396), .A2(n1137), .B1(\intadd_4/n1 ), .B2(n73), .ZN(
        n3308) );
  INV_X1 U4768 ( .A(B[18]), .ZN(n1138) );
  OAI22_X1 U4769 ( .A1(n70), .A2(n1138), .B1(\intadd_3/n1 ), .B2(n74), .ZN(
        n3309) );
  INV_X1 U4770 ( .A(A[21]), .ZN(n1146) );
  FA_X1 U4771 ( .A(n1141), .B(n1140), .CI(n1139), .CO(n1346), .S(n1343) );
  FA_X1 U4772 ( .A(n1144), .B(n1143), .CI(n1142), .CO(n1342), .S(
        \intadd_9/B[2] ) );
  OAI22_X1 U4773 ( .A1(n1396), .A2(n1146), .B1(n1145), .B2(n74), .ZN(n3314) );
  INV_X1 U4774 ( .A(A[13]), .ZN(n1150) );
  OR2_X1 U4775 ( .A1(n1148), .A2(n1147), .ZN(n1320) );
  OAI22_X1 U4776 ( .A1(n1396), .A2(n1150), .B1(n1149), .B2(n73), .ZN(n3331) );
  INV_X1 U4777 ( .A(B[15]), .ZN(n1151) );
  OAI22_X1 U4778 ( .A1(n70), .A2(n1151), .B1(\intadd_2/n1 ), .B2(n74), .ZN(
        n3332) );
  INV_X1 U4779 ( .A(A[14]), .ZN(n1152) );
  OAI22_X1 U4780 ( .A1(n1396), .A2(n1152), .B1(\intadd_2/SUM[3] ), .B2(n74), 
        .ZN(n3333) );
  NAND2_X1 U4781 ( .A1(n1154), .A2(n1432), .ZN(n1158) );
  OAI21_X1 U4782 ( .B1(n1158), .B2(n1526), .A(n1156), .ZN(n3432) );
  AOI22_X1 U4783 ( .A1(s_A_MULT[14]), .A2(n1160), .B1(n1159), .B2(n1257), .ZN(
        n1163) );
  NAND3_X1 U4784 ( .A1(S_B_MULT[11]), .A2(n1161), .A3(n1261), .ZN(n1162) );
  OAI211_X1 U4785 ( .C1(n1165), .C2(n1164), .A(n1163), .B(n1162), .ZN(n1237)
         );
  XOR2_X1 U4786 ( .A(n1266), .B(n1237), .Z(n1271) );
  XNOR2_X1 U4787 ( .A(n1273), .B(n1271), .ZN(n1287) );
  OAI21_X1 U4788 ( .B1(n1269), .B2(n1166), .A(n1267), .ZN(n1167) );
  INV_X1 U4789 ( .A(n1167), .ZN(n1286) );
  FA_X1 U4790 ( .A(n1170), .B(n1169), .CI(n1168), .CO(n1290), .S(n1166) );
  AOI22_X1 U4791 ( .A1(s_A_MULT[10]), .A2(n1246), .B1(n1245), .B2(n1171), .ZN(
        n1172) );
  OAI21_X1 U4792 ( .B1(n61), .B2(n1243), .A(n1172), .ZN(n1173) );
  AOI21_X1 U4793 ( .B1(s_A_MULT[11]), .B2(n1247), .A(n1173), .ZN(n1289) );
  AOI22_X1 U4794 ( .A1(s_A_MULT[12]), .A2(n1259), .B1(n1260), .B2(n1244), .ZN(
        n1174) );
  OAI21_X1 U4795 ( .B1(n63), .B2(n1250), .A(n1174), .ZN(n1175) );
  AOI21_X1 U4796 ( .B1(s_A_MULT[13]), .B2(n1262), .A(n1175), .ZN(n1288) );
  INV_X1 U4797 ( .A(n1176), .ZN(n1360) );
  FA_X1 U4798 ( .A(n1179), .B(n1178), .CI(n1177), .CO(n1180), .S(n1012) );
  INV_X1 U4799 ( .A(n1180), .ZN(n1359) );
  FA_X1 U4800 ( .A(n1183), .B(n1182), .CI(n1181), .CO(n1358), .S(n1339) );
  AOI22_X1 U4801 ( .A1(n72), .A2(n1184), .B1(A[25]), .B2(n1374), .ZN(n1185) );
  INV_X1 U4802 ( .A(n1185), .ZN(n4840) );
  INV_X1 U4803 ( .A(A[4]), .ZN(n1191) );
  NAND2_X1 U4804 ( .A1(n1187), .A2(n1186), .ZN(n1188) );
  XOR2_X1 U4805 ( .A(n1189), .B(n1188), .Z(n1190) );
  OAI22_X1 U4806 ( .A1(n70), .A2(n1191), .B1(n73), .B2(n1190), .ZN(n4841) );
  AOI211_X1 U4807 ( .C1(n1194), .C2(n1193), .A(n1192), .B(n73), .ZN(n1195) );
  AOI21_X1 U4808 ( .B1(A[2]), .B2(n1374), .A(n1195), .ZN(n1196) );
  INV_X1 U4809 ( .A(n1196), .ZN(n4842) );
  INV_X1 U4810 ( .A(A[30]), .ZN(n1207) );
  INV_X1 U4811 ( .A(n1221), .ZN(n1197) );
  NAND2_X1 U4812 ( .A1(n1197), .A2(n1223), .ZN(n1297) );
  XNOR2_X1 U4813 ( .A(n1198), .B(n1297), .ZN(n1210) );
  AOI22_X1 U4814 ( .A1(s_A_MULT[15]), .A2(n1247), .B1(n1239), .B2(n1257), .ZN(
        n1199) );
  OAI21_X1 U4815 ( .B1(n1242), .B2(n1232), .A(n1199), .ZN(n1200) );
  AOI21_X1 U4816 ( .B1(s_A_MULT[14]), .B2(n1246), .A(n1200), .ZN(n1202) );
  XNOR2_X1 U4817 ( .A(n1201), .B(n1202), .ZN(n1213) );
  AOI21_X1 U4818 ( .B1(n1223), .B2(n1213), .A(n1221), .ZN(n1209) );
  INV_X1 U4819 ( .A(n1202), .ZN(n1204) );
  AOI21_X1 U4820 ( .B1(n1205), .B2(n1204), .A(n1203), .ZN(n1208) );
  OAI22_X1 U4821 ( .A1(n1396), .A2(n1207), .B1(n1206), .B2(n73), .ZN(n87) );
  FA_X1 U4822 ( .A(n1210), .B(n1209), .CI(n1208), .CO(n1211), .S(n1206) );
  OAI22_X1 U4823 ( .A1(n70), .A2(n1212), .B1(n1211), .B2(n73), .ZN(n88) );
  INV_X1 U4824 ( .A(B[30]), .ZN(n1225) );
  XOR2_X1 U4825 ( .A(n1213), .B(n1297), .Z(n1228) );
  AOI22_X1 U4826 ( .A1(s_A_MULT[14]), .A2(n1247), .B1(n1239), .B2(n1261), .ZN(
        n1214) );
  OAI21_X1 U4827 ( .B1(n1242), .B2(n1250), .A(n1214), .ZN(n1215) );
  AOI21_X1 U4828 ( .B1(s_A_MULT[13]), .B2(n1246), .A(n1215), .ZN(n1219) );
  INV_X1 U4829 ( .A(n1216), .ZN(n1217) );
  AOI21_X1 U4830 ( .B1(n1260), .B2(n1257), .A(n1217), .ZN(n1218) );
  FA_X1 U4831 ( .A(n1220), .B(n1219), .CI(n1218), .CO(n1227), .S(n1298) );
  INV_X1 U4832 ( .A(n1298), .ZN(n1222) );
  AOI21_X1 U4833 ( .B1(n1223), .B2(n1222), .A(n1221), .ZN(n1226) );
  OAI22_X1 U4834 ( .A1(n1396), .A2(n1225), .B1(n1224), .B2(n74), .ZN(n89) );
  FA_X1 U4835 ( .A(n1228), .B(n1227), .CI(n1226), .CO(n1224), .S(n1229) );
  NOR2_X1 U4836 ( .A1(n1229), .A2(n73), .ZN(n1230) );
  AOI21_X1 U4837 ( .B1(A[29]), .B2(n1374), .A(n1230), .ZN(n900) );
  INV_X1 U4838 ( .A(A[27]), .ZN(n1281) );
  OAI22_X1 U4839 ( .A1(n63), .A2(n1232), .B1(n1231), .B2(n1250), .ZN(n1233) );
  AOI21_X1 U4840 ( .B1(s_A_MULT[14]), .B2(n1262), .A(n1233), .ZN(n1234) );
  OAI21_X1 U4841 ( .B1(n1236), .B2(n1235), .A(n1234), .ZN(n1277) );
  OAI21_X1 U4842 ( .B1(n1237), .B2(n1255), .A(n1254), .ZN(n1238) );
  INV_X1 U4843 ( .A(n1238), .ZN(n1276) );
  AOI22_X1 U4844 ( .A1(s_A_MULT[11]), .A2(n1246), .B1(n1239), .B2(n1244), .ZN(
        n1241) );
  NAND2_X1 U4845 ( .A1(s_A_MULT[12]), .A2(n1247), .ZN(n1240) );
  OAI211_X1 U4846 ( .C1(n1243), .C2(n1242), .A(n1241), .B(n1240), .ZN(n1275)
         );
  AOI22_X1 U4847 ( .A1(s_A_MULT[12]), .A2(n1246), .B1(n1245), .B2(n1244), .ZN(
        n1249) );
  NAND2_X1 U4848 ( .A1(s_A_MULT[13]), .A2(n1247), .ZN(n1248) );
  OAI211_X1 U4849 ( .C1(n1250), .C2(n61), .A(n1249), .B(n1248), .ZN(n1301) );
  OAI21_X1 U4850 ( .B1(n1253), .B2(n1252), .A(n1251), .ZN(n1265) );
  OAI21_X1 U4851 ( .B1(n1265), .B2(n1255), .A(n1254), .ZN(n1256) );
  INV_X1 U4852 ( .A(n1256), .ZN(n1300) );
  AOI22_X1 U4853 ( .A1(s_A_MULT[14]), .A2(n1259), .B1(n1258), .B2(n1257), .ZN(
        n1264) );
  AOI22_X1 U4854 ( .A1(s_A_MULT[15]), .A2(n1262), .B1(n1261), .B2(n1260), .ZN(
        n1263) );
  NAND2_X1 U4855 ( .A1(n1264), .A2(n1263), .ZN(n1299) );
  XNOR2_X1 U4856 ( .A(n1266), .B(n1265), .ZN(n1274) );
  OAI21_X1 U4857 ( .B1(n1269), .B2(n1274), .A(n1267), .ZN(n1295) );
  XNOR2_X1 U4858 ( .A(n1268), .B(n1273), .ZN(n1294) );
  XNOR2_X1 U4859 ( .A(n1380), .B(n1379), .ZN(n1279) );
  INV_X1 U4860 ( .A(n1269), .ZN(n1272) );
  AOI21_X1 U4861 ( .B1(n1272), .B2(n1271), .A(n1270), .ZN(n1284) );
  XOR2_X1 U4862 ( .A(n1274), .B(n1273), .Z(n1283) );
  FA_X1 U4863 ( .A(n1277), .B(n1276), .CI(n1275), .CO(n1380), .S(n1278) );
  INV_X1 U4864 ( .A(n1278), .ZN(n1282) );
  XNOR2_X1 U4865 ( .A(n1279), .B(n1377), .ZN(n1280) );
  OAI22_X1 U4866 ( .A1(n70), .A2(n1281), .B1(n1280), .B2(n74), .ZN(n93) );
  INV_X1 U4867 ( .A(A[26]), .ZN(n1293) );
  FA_X1 U4868 ( .A(n1284), .B(n1283), .CI(n1282), .CO(n1377), .S(n1363) );
  FA_X1 U4869 ( .A(n1287), .B(n1286), .CI(n1285), .CO(n1365), .S(n1176) );
  FA_X1 U4870 ( .A(n1290), .B(n1289), .CI(n1288), .CO(n1364), .S(n1285) );
  NAND2_X1 U4871 ( .A1(n1365), .A2(n1364), .ZN(n1367) );
  OAI21_X1 U4872 ( .B1(n1365), .B2(n1364), .A(n1367), .ZN(n1291) );
  XNOR2_X1 U4873 ( .A(n1363), .B(n1291), .ZN(n1292) );
  OAI22_X1 U4874 ( .A1(n1396), .A2(n1293), .B1(n73), .B2(n1292), .ZN(n96) );
  FA_X1 U4875 ( .A(n1296), .B(n1295), .CI(n1294), .CO(n1373), .S(n1379) );
  XOR2_X1 U4876 ( .A(n1298), .B(n1297), .Z(n1372) );
  FA_X1 U4877 ( .A(n1301), .B(n1300), .CI(n1299), .CO(n1371), .S(n1296) );
  AOI22_X1 U4878 ( .A1(n72), .A2(n1302), .B1(A[28]), .B2(n1374), .ZN(n1303) );
  INV_X1 U4879 ( .A(n1303), .ZN(n7620) );
  FA_X1 U4880 ( .A(n1306), .B(n1305), .CI(n1304), .CO(n1139), .S(n7619) );
  INV_X1 U4881 ( .A(n1), .ZN(n6433) );
  INV_X1 U4882 ( .A(s_A_ADDER[2]), .ZN(n6432) );
  INV_X1 U4883 ( .A(s_A_ADDER[3]), .ZN(n6431) );
  INV_X1 U4884 ( .A(s_A_ADDER[4]), .ZN(n6430) );
  INV_X1 U4885 ( .A(s_A_ADDER[5]), .ZN(n6429) );
  INV_X1 U4886 ( .A(s_A_ADDER[6]), .ZN(n6428) );
  INV_X1 U4887 ( .A(s_A_ADDER[7]), .ZN(n6427) );
  INV_X1 U4888 ( .A(s_A_ADDER[8]), .ZN(n6426) );
  INV_X1 U4889 ( .A(s_A_ADDER[9]), .ZN(n6425) );
  INV_X1 U4890 ( .A(A[1]), .ZN(n1311) );
  AOI222_X1 U4891 ( .A1(s_A_MULT[1]), .A2(n1309), .B1(\MULT/SHIFTERi_0/N19 ), 
        .B2(n55), .C1(n1308), .C2(n1307), .ZN(n1310) );
  OAI22_X1 U4892 ( .A1(n70), .A2(n1311), .B1(n1310), .B2(n73), .ZN(n6346) );
  INV_X1 U4893 ( .A(B[10]), .ZN(n1315) );
  INV_X1 U4894 ( .A(\intadd_12/SUM[2] ), .ZN(n1312) );
  NAND2_X1 U4895 ( .A1(n1313), .A2(n1312), .ZN(n1314) );
  OAI22_X1 U4896 ( .A1(n1396), .A2(n1315), .B1(n74), .B2(n1314), .ZN(n6339) );
  INV_X1 U4897 ( .A(B[11]), .ZN(n1316) );
  OR2_X1 U4898 ( .A1(\intadd_11/SUM[2] ), .A2(\intadd_12/n1 ), .ZN(n1317) );
  OAI22_X1 U4899 ( .A1(n1396), .A2(n1316), .B1(n73), .B2(n1317), .ZN(n6337) );
  AOI21_X1 U4900 ( .B1(\intadd_11/SUM[2] ), .B2(\intadd_12/n1 ), .A(n74), .ZN(
        n1318) );
  AOI22_X1 U4901 ( .A1(n1318), .A2(n1317), .B1(A[10]), .B2(n1374), .ZN(n1319)
         );
  INV_X1 U4902 ( .A(n1319), .ZN(n6336) );
  INV_X1 U4903 ( .A(B[14]), .ZN(n1322) );
  FA_X1 U4904 ( .A(\intadd_10/n1 ), .B(\intadd_2/SUM[2] ), .CI(n1320), .CO(
        n1321), .S(n1149) );
  OAI22_X1 U4905 ( .A1(n70), .A2(n1322), .B1(n1321), .B2(n74), .ZN(n6334) );
  INV_X1 U4906 ( .A(B[16]), .ZN(n1325) );
  FA_X1 U4907 ( .A(\intadd_6/n1 ), .B(\intadd_5/SUM[2] ), .CI(n1323), .CO(
        n1324), .S(n1133) );
  OAI22_X1 U4908 ( .A1(n70), .A2(n1325), .B1(n1324), .B2(n74), .ZN(n6333) );
  INV_X1 U4909 ( .A(A[16]), .ZN(n1330) );
  FA_X1 U4910 ( .A(n1328), .B(n1327), .CI(n1326), .CO(n1331), .S(
        \intadd_5/A[2] ) );
  OAI22_X1 U4911 ( .A1(n1396), .A2(n1330), .B1(n1329), .B2(n74), .ZN(n6331) );
  INV_X1 U4912 ( .A(B[17]), .ZN(n1333) );
  FA_X1 U4913 ( .A(\intadd_5/n1 ), .B(\intadd_3/SUM[2] ), .CI(n1331), .CO(
        n1332), .S(n1329) );
  OAI22_X1 U4914 ( .A1(n70), .A2(n1333), .B1(n1332), .B2(n74), .ZN(n6330) );
  INV_X1 U4915 ( .A(B[21]), .ZN(n1336) );
  FA_X1 U4916 ( .A(\intadd_9/SUM[2] ), .B(\intadd_8/n1 ), .CI(n1334), .CO(
        n1335), .S(n1113) );
  OAI22_X1 U4917 ( .A1(n1396), .A2(n1336), .B1(n1335), .B2(n74), .ZN(n6329) );
  FA_X1 U4918 ( .A(n1339), .B(n1338), .CI(n1337), .CO(n1340), .S(n1031) );
  AOI22_X1 U4919 ( .A1(n1617), .A2(n1340), .B1(B[25]), .B2(n1374), .ZN(n1341)
         );
  INV_X1 U4920 ( .A(n1341), .ZN(n6327) );
  INV_X1 U4921 ( .A(B[22]), .ZN(n1345) );
  FA_X1 U4922 ( .A(\intadd_9/n1 ), .B(n1343), .CI(n1342), .CO(n1344), .S(n1145) );
  OAI22_X1 U4923 ( .A1(n1396), .A2(n1345), .B1(n1344), .B2(n74), .ZN(n6326) );
  AOI222_X1 U4924 ( .A1(n1348), .A2(n1347), .B1(n1348), .B2(n1346), .C1(n1347), 
        .C2(n1346), .ZN(n1349) );
  AOI22_X1 U4925 ( .A1(n72), .A2(n1349), .B1(B[23]), .B2(n1374), .ZN(n1350) );
  INV_X1 U4926 ( .A(n1350), .ZN(n6325) );
  INV_X1 U4927 ( .A(B[24]), .ZN(n1357) );
  NAND2_X1 U4928 ( .A1(n1352), .A2(n1351), .ZN(n1354) );
  AOI21_X1 U4929 ( .B1(n1355), .B2(n1354), .A(n1353), .ZN(n1356) );
  OAI22_X1 U4930 ( .A1(n70), .A2(n1357), .B1(n1356), .B2(n74), .ZN(n6324) );
  FA_X1 U4931 ( .A(n1360), .B(n1359), .CI(n1358), .CO(n1361), .S(n1184) );
  AOI22_X1 U4932 ( .A1(n72), .A2(n1361), .B1(B[26]), .B2(n1374), .ZN(n1362) );
  INV_X1 U4933 ( .A(n1362), .ZN(n6323) );
  INV_X1 U4934 ( .A(B[27]), .ZN(n1370) );
  INV_X1 U4935 ( .A(n1363), .ZN(n1368) );
  NOR2_X1 U4936 ( .A1(n1365), .A2(n1364), .ZN(n1366) );
  AOI21_X1 U4937 ( .B1(n1368), .B2(n1367), .A(n1366), .ZN(n1369) );
  OAI22_X1 U4938 ( .A1(n70), .A2(n1370), .B1(n1369), .B2(n74), .ZN(n6322) );
  FA_X1 U4939 ( .A(n1373), .B(n1372), .CI(n1371), .CO(n1375), .S(n1302) );
  AOI22_X1 U4940 ( .A1(n1617), .A2(n1375), .B1(B[29]), .B2(n1416), .ZN(n1376)
         );
  INV_X1 U4941 ( .A(n1376), .ZN(n6321) );
  INV_X1 U4942 ( .A(B[28]), .ZN(n1382) );
  INV_X1 U4943 ( .A(n1377), .ZN(n1378) );
  AOI222_X1 U4944 ( .A1(n1380), .A2(n1379), .B1(n1380), .B2(n1378), .C1(n1379), 
        .C2(n1378), .ZN(n1381) );
  OAI22_X1 U4945 ( .A1(n1396), .A2(n1382), .B1(n1381), .B2(n74), .ZN(n6320) );
  INV_X1 U4946 ( .A(B[7]), .ZN(n1387) );
  NAND3_X1 U4947 ( .A1(n1385), .A2(n1384), .A3(n1383), .ZN(n1386) );
  OAI22_X1 U4948 ( .A1(n70), .A2(n1387), .B1(n74), .B2(n1386), .ZN(N61) );
  INV_X1 U4949 ( .A(B[9]), .ZN(n1391) );
  NAND2_X1 U4950 ( .A1(n1389), .A2(n1388), .ZN(n1390) );
  OAI22_X1 U4951 ( .A1(n1396), .A2(n1391), .B1(n73), .B2(n1390), .ZN(N63) );
  INV_X1 U4952 ( .A(B[12]), .ZN(n1395) );
  INV_X1 U4953 ( .A(\intadd_11/n1 ), .ZN(n1392) );
  NAND2_X1 U4954 ( .A1(n1393), .A2(n1392), .ZN(n1394) );
  OAI22_X1 U4955 ( .A1(n1396), .A2(n1395), .B1(n74), .B2(n1394), .ZN(N66) );
  BUF_X1 U3448 ( .A(n1429), .Z(n1398) );
  CLKBUF_X1 U3452 ( .A(n695), .Z(n1397) );
  CLKBUF_X3 U3455 ( .A(n1429), .Z(n1399) );
  AND2_X1 U3459 ( .A1(N87), .A2(s_LOGIC[1]), .ZN(n1429) );
  NAND2_X2 U3460 ( .A1(n687), .A2(n736), .ZN(n538) );
  INV_X1 U3461 ( .A(n1441), .ZN(n1400) );
  CLKBUF_X1 U3464 ( .A(n328), .Z(n1441) );
  INV_X1 U3466 ( .A(n1432), .ZN(n1401) );
  BUF_X4 U3468 ( .A(n1616), .Z(n75) );
  AOI222_X1 U3484 ( .A1(n1418), .A2(n652), .B1(n718), .B2(n651), .C1(n650), 
        .C2(n665), .ZN(n5) );
  AND2_X1 U3494 ( .A1(n718), .A2(n517), .ZN(n1440) );
  OR2_X1 U3495 ( .A1(n1428), .A2(n1492), .ZN(n388) );
  OR2_X1 U3499 ( .A1(n1399), .A2(n1490), .ZN(n400) );
  OAI21_X1 U3529 ( .B1(n1428), .B2(n1501), .A(n1500), .ZN(n1499) );
  AND2_X1 U3535 ( .A1(n1398), .A2(n1487), .ZN(n11) );
  NAND2_X2 U3538 ( .A1(n702), .A2(n736), .ZN(n714) );
  NOR2_X1 U3555 ( .A1(n1428), .A2(n1503), .ZN(n1502) );
  AND2_X1 U3556 ( .A1(n1428), .A2(n1488), .ZN(n19) );
  OR2_X1 U3558 ( .A1(n1428), .A2(n1489), .ZN(n377) );
  OR2_X1 U3561 ( .A1(n1399), .A2(n1491), .ZN(n365) );
  OR2_X1 U3562 ( .A1(n1399), .A2(n1493), .ZN(n8) );
  NAND2_X2 U3563 ( .A1(n1466), .A2(n1469), .ZN(n1402) );
  NAND2_X1 U3564 ( .A1(n1466), .A2(n1469), .ZN(n1403) );
  NAND2_X1 U3565 ( .A1(n1466), .A2(n1469), .ZN(n737) );
  CLKBUF_X1 U3566 ( .A(n6451), .Z(n1404) );
  INV_X1 U3568 ( .A(n335), .ZN(n6451) );
  CLKBUF_X1 U3570 ( .A(n1404), .Z(n71) );
  NAND2_X1 U3572 ( .A1(n1467), .A2(n1465), .ZN(n1466) );
  INV_X1 U3596 ( .A(n649), .ZN(n1405) );
  INV_X1 U3598 ( .A(n649), .ZN(n1406) );
  INV_X1 U3604 ( .A(n649), .ZN(n732) );
  NOR2_X1 U3605 ( .A1(n515), .A2(n1439), .ZN(n518) );
  OR2_X1 U3853 ( .A1(n1399), .A2(n1486), .ZN(n655) );
  OR2_X1 U3861 ( .A1(n58), .A2(n1484), .ZN(n667) );
  OR2_X1 U3862 ( .A1(n58), .A2(n1485), .ZN(n607) );
  NAND2_X1 U3954 ( .A1(n1474), .A2(n1473), .ZN(n720) );
  OAI22_X1 U3980 ( .A1(n728), .A2(n556), .B1(n695), .B2(n488), .ZN(n1458) );
  NOR2_X1 U3983 ( .A1(n1458), .A2(n1517), .ZN(n1457) );
  NAND4_X1 U3989 ( .A1(n1413), .A2(n1410), .A3(n1408), .A4(n1407), .ZN(Y[3])
         );
  NAND2_X1 U4003 ( .A1(n716), .A2(n701), .ZN(n1407) );
  INV_X1 U4031 ( .A(n1409), .ZN(n1408) );
  NOR2_X1 U4037 ( .A1(n711), .A2(n661), .ZN(n1409) );
  AOI211_X1 U4039 ( .C1(n654), .C2(n688), .A(n1412), .B(n1411), .ZN(n1410) );
  AND2_X1 U4048 ( .A1(n1434), .A2(n672), .ZN(n1411) );
  NOR2_X1 U4050 ( .A1(n1406), .A2(\intadd_1/SUM[1] ), .ZN(n1412) );
  NAND2_X1 U4055 ( .A1(n655), .A2(n1414), .ZN(n1413) );
  INV_X1 U4064 ( .A(n1415), .ZN(n1414) );
  OAI22_X1 U4067 ( .A1(n1403), .A2(n656), .B1(S_B_LOGIC[3]), .B2(s_A_LOGIC[3]), 
        .ZN(n1415) );
  INV_X1 U4080 ( .A(n1396), .ZN(n1416) );
  NOR2_X1 U4086 ( .A1(n1516), .A2(n1618), .ZN(n335) );
  NAND3_X2 U4096 ( .A1(n1153), .A2(n1154), .A3(OP[3]), .ZN(n424) );
  INV_X1 U4114 ( .A(n1454), .ZN(n1417) );
  CLKBUF_X1 U4115 ( .A(n330), .Z(n1454) );
  INV_X1 U4116 ( .A(n1524), .ZN(n423) );
  NAND2_X1 U4117 ( .A1(n1520), .A2(n1524), .ZN(n1157) );
  NAND2_X1 U4130 ( .A1(n1474), .A2(n1473), .ZN(n1418) );
  NAND2_X1 U4131 ( .A1(n1474), .A2(n1473), .ZN(n1419) );
  AOI211_X4 U4134 ( .C1(n1419), .C2(n407), .A(n406), .B(n405), .ZN(n408) );
  OAI21_X1 U4135 ( .B1(n1452), .B2(n1405), .A(n1156), .ZN(n1374) );
  OR2_X1 U4138 ( .A1(n1405), .A2(n434), .ZN(n1446) );
  INV_X1 U4143 ( .A(n726), .ZN(n654) );
  NOR2_X1 U4147 ( .A1(n35), .A2(n1449), .ZN(n36) );
  OR2_X1 U4165 ( .A1(n33), .A2(n1450), .ZN(n1449) );
  INV_X1 U4180 ( .A(n737), .ZN(n1420) );
  INV_X1 U4192 ( .A(n1499), .ZN(n470) );
  NAND2_X1 U4196 ( .A1(n687), .A2(n720), .ZN(n1421) );
  NAND2_X1 U4284 ( .A1(n687), .A2(n1419), .ZN(n614) );
  OR2_X1 U4313 ( .A1(n711), .A2(n454), .ZN(n1422) );
  NAND2_X1 U4315 ( .A1(n702), .A2(n720), .ZN(n1423) );
  NOR2_X1 U4316 ( .A1(n382), .A2(n383), .ZN(n1424) );
  NOR3_X1 U4317 ( .A1(n381), .A2(n384), .A3(n1425), .ZN(n385) );
  INV_X1 U4318 ( .A(n1424), .ZN(n1425) );
  NAND2_X1 U4319 ( .A1(n702), .A2(n720), .ZN(n678) );
  AND2_X1 U4324 ( .A1(n466), .A2(n1433), .ZN(n1426) );
  NOR2_X1 U4956 ( .A1(n1426), .A2(n1462), .ZN(n1461) );
  INV_X2 U4957 ( .A(n666), .ZN(n1427) );
  INV_X1 U4958 ( .A(n666), .ZN(n730) );
  INV_X1 U4959 ( .A(n1508), .ZN(n1453) );
  CLKBUF_X1 U4960 ( .A(OP[3]), .Z(n1452) );
  NAND2_X1 U4961 ( .A1(OP[3]), .A2(n1512), .ZN(n1511) );
  AND2_X1 U4962 ( .A1(n246), .A2(n247), .ZN(n1516) );
  INV_X1 U4963 ( .A(OP[3]), .ZN(n1520) );
  AND2_X1 U4964 ( .A1(n246), .A2(s_LOGIC[3]), .ZN(n1465) );
  INV_X1 U4965 ( .A(n737), .ZN(n544) );
  AND2_X2 U4966 ( .A1(N87), .A2(s_LOGIC[1]), .ZN(n1428) );
  AND2_X1 U4967 ( .A1(N87), .A2(s_LOGIC[1]), .ZN(n58) );
  NOR2_X1 U4968 ( .A1(n325), .A2(n424), .ZN(n1618) );
  CLKBUF_X1 U4969 ( .A(OP[4]), .Z(n1430) );
  NAND2_X1 U4970 ( .A1(n328), .A2(n330), .ZN(n325) );
  INV_X1 U4971 ( .A(OP[1]), .ZN(n1437) );
  CLKBUF_X2 U4972 ( .A(n1136), .Z(n1451) );
  INV_X1 U4973 ( .A(n1136), .ZN(n1519) );
  NAND2_X1 U4974 ( .A1(n1524), .A2(n1521), .ZN(n1431) );
  INV_X1 U4975 ( .A(OP[2]), .ZN(n330) );
  OR2_X1 U4976 ( .A1(n58), .A2(n1483), .ZN(n510) );
  NOR2_X2 U4977 ( .A1(n424), .A2(n423), .ZN(n1616) );
  INV_X1 U4978 ( .A(OP[0]), .ZN(n1432) );
  INV_X1 U4979 ( .A(n728), .ZN(n1433) );
  BUF_X1 U4980 ( .A(n736), .Z(n1434) );
  INV_X1 U4981 ( .A(OP[0]), .ZN(n1153) );
  OAI21_X2 U4982 ( .B1(n1510), .B2(n1511), .A(n1513), .ZN(n736) );
  AOI21_X1 U4983 ( .B1(n1420), .B2(n1532), .A(n1531), .ZN(n1530) );
  NAND2_X1 U4984 ( .A1(n544), .A2(S_B_LOGIC[1]), .ZN(n1500) );
  NAND2_X1 U4985 ( .A1(n1479), .A2(n1478), .ZN(n1474) );
  NOR2_X1 U4986 ( .A1(n424), .A2(n1529), .ZN(n1479) );
  AND2_X1 U4987 ( .A1(n75), .A2(S_B_LHI[3]), .ZN(n1533) );
  INV_X1 U4988 ( .A(n58), .ZN(n1435) );
  INV_X1 U4989 ( .A(n1398), .ZN(n1436) );
  INV_X1 U4990 ( .A(n1494), .ZN(n492) );
  NOR2_X2 U4991 ( .A1(n1437), .A2(OP[2]), .ZN(n1524) );
  NAND3_X1 U4992 ( .A1(n1466), .A2(n1431), .A3(S_B_LOGIC[21]), .ZN(n1438) );
  OAI21_X1 U4993 ( .B1(n1428), .B2(n1498), .A(n1438), .ZN(n1497) );
  OR2_X2 U4994 ( .A1(n516), .A2(n1440), .ZN(n1439) );
  NAND4_X2 U4995 ( .A1(n1442), .A2(n1446), .A3(n1443), .A4(n438), .ZN(Y[16])
         );
  AND2_X2 U4996 ( .A1(n1447), .A2(n1444), .ZN(n1442) );
  AOI21_X1 U4997 ( .B1(n716), .B2(n517), .A(n1445), .ZN(n1444) );
  NOR2_X1 U4998 ( .A1(n711), .A2(n439), .ZN(n1445) );
  BUF_X2 U4999 ( .A(n1455), .Z(n1443) );
  NAND2_X1 U5000 ( .A1(n1530), .A2(n1448), .ZN(n1447) );
  OR2_X1 U5001 ( .A1(n1428), .A2(S_B_LOGIC[16]), .ZN(n1448) );
  AND2_X2 U5002 ( .A1(n649), .A2(n30), .ZN(n1450) );
  NAND3_X1 U5003 ( .A1(n1453), .A2(n1461), .A3(n452), .ZN(n1460) );
  NAND2_X1 U5004 ( .A1(n544), .A2(S_B_LOGIC[20]), .ZN(n1495) );
  OAI21_X1 U5005 ( .B1(n1428), .B2(n1496), .A(n1495), .ZN(n1494) );
  NAND2_X2 U5006 ( .A1(n736), .A2(n663), .ZN(n728) );
  INV_X2 U5007 ( .A(n436), .ZN(n1455) );
  OR4_X2 U5008 ( .A1(n14), .A2(n1456), .A3(n1533), .A4(n15), .ZN(Y[19]) );
  NAND3_X1 U5009 ( .A1(n1459), .A2(n1457), .A3(n17), .ZN(n1456) );
  INV_X2 U5010 ( .A(n11), .ZN(n1459) );
  OR2_X1 U5011 ( .A1(n1460), .A2(n1504), .ZN(Y[18]) );
  NAND2_X1 U5012 ( .A1(n458), .A2(n1463), .ZN(n1462) );
  INV_X1 U5013 ( .A(n1464), .ZN(n1463) );
  NOR2_X1 U5014 ( .A1(n730), .A2(n460), .ZN(n1464) );
  NAND2_X1 U5015 ( .A1(n1467), .A2(n246), .ZN(n242) );
  INV_X1 U5016 ( .A(n1468), .ZN(n1467) );
  NAND2_X1 U5017 ( .A1(n328), .A2(OP[2]), .ZN(n1468) );
  NAND2_X1 U5018 ( .A1(n1521), .A2(n1524), .ZN(n1469) );
  NAND2_X1 U5019 ( .A1(n1516), .A2(n1480), .ZN(n1473) );
  NAND2_X1 U5020 ( .A1(n1478), .A2(n1470), .ZN(n1477) );
  NOR2_X1 U5021 ( .A1(n424), .A2(n1471), .ZN(n1470) );
  NAND2_X1 U5022 ( .A1(n1528), .A2(n1472), .ZN(n1471) );
  INV_X1 U5023 ( .A(n1529), .ZN(n1472) );
  INV_X1 U5024 ( .A(n325), .ZN(n1478) );
  NAND2_X1 U5025 ( .A1(n1516), .A2(n1476), .ZN(n1475) );
  NAND2_X2 U5026 ( .A1(n1477), .A2(n1475), .ZN(n666) );
  AND2_X2 U5027 ( .A1(n1480), .A2(n1528), .ZN(n1476) );
  INV_X2 U5028 ( .A(n1529), .ZN(n1480) );
  OR2_X2 U5029 ( .A1(n335), .A2(n1481), .ZN(n726) );
  NAND2_X2 U5030 ( .A1(n686), .A2(n1482), .ZN(n1481) );
  INV_X2 U5031 ( .A(n1529), .ZN(n1482) );
  INV_X2 U5032 ( .A(n511), .ZN(n1483) );
  INV_X2 U5033 ( .A(n668), .ZN(n1484) );
  INV_X2 U5034 ( .A(n608), .ZN(n1485) );
  INV_X2 U5035 ( .A(n656), .ZN(n1486) );
  NOR2_X2 U5036 ( .A1(s_A_LOGIC[19]), .A2(n10), .ZN(n1487) );
  NOR2_X2 U5037 ( .A1(s_A_LOGIC[17]), .A2(n18), .ZN(n1488) );
  INV_X2 U5038 ( .A(n378), .ZN(n1489) );
  INV_X2 U5039 ( .A(n401), .ZN(n1490) );
  INV_X2 U5040 ( .A(n366), .ZN(n1491) );
  INV_X2 U5041 ( .A(n389), .ZN(n1492) );
  INV_X2 U5042 ( .A(n7), .ZN(n1493) );
  INV_X2 U5043 ( .A(n487), .ZN(n1496) );
  INV_X2 U5044 ( .A(n1497), .ZN(n505) );
  INV_X2 U5045 ( .A(n501), .ZN(n1498) );
  INV_X2 U5046 ( .A(n468), .ZN(n1501) );
  NOR2_X2 U5047 ( .A1(n49), .A2(n1502), .ZN(n50) );
  INV_X2 U5048 ( .A(n48), .ZN(n1503) );
  OAI21_X1 U5049 ( .B1(n1435), .B2(n1506), .A(n1505), .ZN(n1504) );
  NAND2_X1 U5050 ( .A1(n75), .A2(S_B_LHI[2]), .ZN(n1505) );
  NAND2_X1 U5051 ( .A1(S_B_LOGIC[18]), .A2(n1507), .ZN(n1506) );
  INV_X1 U5052 ( .A(s_A_LOGIC[18]), .ZN(n1507) );
  NAND2_X1 U5053 ( .A1(n1509), .A2(n1422), .ZN(n1508) );
  INV_X1 U5054 ( .A(n456), .ZN(n1509) );
  NAND3_X1 U5055 ( .A1(n246), .A2(n247), .A3(n1514), .ZN(n1513) );
  NAND4_X1 U5056 ( .A1(n328), .A2(n1153), .A3(n1154), .A4(n330), .ZN(n1510) );
  INV_X2 U5057 ( .A(n334), .ZN(n1512) );
  INV_X2 U5058 ( .A(n334), .ZN(n1514) );
  CLKBUF_X1 U5059 ( .A(n325), .Z(n1515) );
  AND2_X2 U5060 ( .A1(n666), .A2(n466), .ZN(n1517) );
  OAI21_X1 U5061 ( .B1(n1518), .B2(n423), .A(n242), .ZN(N87) );
  NAND2_X2 U5062 ( .A1(n1519), .A2(n1520), .ZN(n1518) );
  NOR2_X1 U5063 ( .A1(n1136), .A2(n1522), .ZN(n1521) );
  OR2_X1 U5064 ( .A1(OP[3]), .A2(n1523), .ZN(n1522) );
  INV_X1 U5065 ( .A(s_LOGIC[3]), .ZN(n1523) );
  CLKBUF_X1 U5066 ( .A(N87), .Z(n1525) );
  CLKBUF_X1 U5067 ( .A(n1157), .Z(n1526) );
  CLKBUF_X1 U5068 ( .A(n1525), .Z(n1527) );
  INV_X2 U5069 ( .A(n720), .ZN(n711) );
  INV_X2 U5070 ( .A(n1534), .ZN(n1528) );
  INV_X2 U5071 ( .A(n334), .ZN(n1529) );
  INV_X2 U5072 ( .A(s_A_LOGIC[16]), .ZN(n1531) );
  INV_X2 U5073 ( .A(n432), .ZN(n1532) );
  INV_X2 U5074 ( .A(n663), .ZN(n1534) );
  CLKBUF_X1 U5075 ( .A(n1527), .Z(n1535) );
  NOR2_X2 U5076 ( .A1(n966), .A2(n968), .ZN(n1536) );
  INV_X2 U5077 ( .A(n967), .ZN(n1537) );
  MUX2_X1 U5078 ( .A(n1536), .B(n1537), .S(n1164), .Z(n1055) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_0 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_31 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_30 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_29 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_28 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_27 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_26 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_25 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_24 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_23 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_22 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_21 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_20 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_19 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_18 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_17 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_16 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_15 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_14 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_13 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_12 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_11 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_10 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_9 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_8 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_7 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_6 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_5 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_4 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_3 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_2 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_1 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7088, net7090, net7092, net7093, net7096, net7099;
  assign net7088 = EN;
  assign net7090 = CLK;
  assign ENCLK = net7092;
  assign net7099 = TE;

  DLL_X1 latch ( .D(net7093), .GN(net7090), .Q(net7096) );
  OR2_X1 test_or ( .A1(net7088), .A2(net7099), .ZN(net7093) );
  AND2_X1 main_gate ( .A1(net7096), .A2(net7090), .ZN(net7092) );
endmodule


module REGISTER_FILE_WIDTH32_LENGTH5 ( CLK, RST, EN, RD1, RD2, WR, DATAIN, 
        OUT1, OUT2, ADD_WR, ADD_RD1, ADD_RD2 );
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input CLK, RST, EN, RD1, RD2, WR;
  wire   \REGISTERS[0][31] , \REGISTERS[0][30] , \REGISTERS[0][29] ,
         \REGISTERS[0][28] , \REGISTERS[0][27] , \REGISTERS[0][26] ,
         \REGISTERS[0][25] , \REGISTERS[0][24] , \REGISTERS[0][23] ,
         \REGISTERS[0][22] , \REGISTERS[0][21] , \REGISTERS[0][20] ,
         \REGISTERS[0][19] , \REGISTERS[0][18] , \REGISTERS[0][17] ,
         \REGISTERS[0][16] , \REGISTERS[0][15] , \REGISTERS[0][14] ,
         \REGISTERS[0][13] , \REGISTERS[0][12] , \REGISTERS[0][11] ,
         \REGISTERS[0][10] , \REGISTERS[0][9] , \REGISTERS[0][8] ,
         \REGISTERS[0][7] , \REGISTERS[0][6] , \REGISTERS[0][5] ,
         \REGISTERS[0][4] , \REGISTERS[0][3] , \REGISTERS[0][2] ,
         \REGISTERS[0][1] , \REGISTERS[0][0] , \REGISTERS[1][31] ,
         \REGISTERS[1][30] , \REGISTERS[1][29] , \REGISTERS[1][28] ,
         \REGISTERS[1][27] , \REGISTERS[1][26] , \REGISTERS[1][25] ,
         \REGISTERS[1][24] , \REGISTERS[1][23] , \REGISTERS[1][22] ,
         \REGISTERS[1][21] , \REGISTERS[1][20] , \REGISTERS[1][19] ,
         \REGISTERS[1][18] , \REGISTERS[1][17] , \REGISTERS[1][16] ,
         \REGISTERS[1][15] , \REGISTERS[1][14] , \REGISTERS[1][13] ,
         \REGISTERS[1][12] , \REGISTERS[1][11] , \REGISTERS[1][10] ,
         \REGISTERS[1][9] , \REGISTERS[1][8] , \REGISTERS[1][7] ,
         \REGISTERS[1][6] , \REGISTERS[1][5] , \REGISTERS[1][4] ,
         \REGISTERS[1][3] , \REGISTERS[1][2] , \REGISTERS[1][1] ,
         \REGISTERS[1][0] , \REGISTERS[2][31] , \REGISTERS[2][30] ,
         \REGISTERS[2][29] , \REGISTERS[2][28] , \REGISTERS[2][27] ,
         \REGISTERS[2][26] , \REGISTERS[2][25] , \REGISTERS[2][24] ,
         \REGISTERS[2][23] , \REGISTERS[2][22] , \REGISTERS[2][21] ,
         \REGISTERS[2][20] , \REGISTERS[2][19] , \REGISTERS[2][18] ,
         \REGISTERS[2][17] , \REGISTERS[2][16] , \REGISTERS[2][15] ,
         \REGISTERS[2][14] , \REGISTERS[2][13] , \REGISTERS[2][12] ,
         \REGISTERS[2][11] , \REGISTERS[2][10] , \REGISTERS[2][9] ,
         \REGISTERS[2][8] , \REGISTERS[2][7] , \REGISTERS[2][6] ,
         \REGISTERS[2][5] , \REGISTERS[2][4] , \REGISTERS[2][3] ,
         \REGISTERS[2][2] , \REGISTERS[2][1] , \REGISTERS[2][0] ,
         \REGISTERS[3][31] , \REGISTERS[3][30] , \REGISTERS[3][29] ,
         \REGISTERS[3][28] , \REGISTERS[3][27] , \REGISTERS[3][26] ,
         \REGISTERS[3][25] , \REGISTERS[3][24] , \REGISTERS[3][23] ,
         \REGISTERS[3][22] , \REGISTERS[3][21] , \REGISTERS[3][20] ,
         \REGISTERS[3][19] , \REGISTERS[3][18] , \REGISTERS[3][17] ,
         \REGISTERS[3][16] , \REGISTERS[3][15] , \REGISTERS[3][14] ,
         \REGISTERS[3][13] , \REGISTERS[3][12] , \REGISTERS[3][11] ,
         \REGISTERS[3][10] , \REGISTERS[3][9] , \REGISTERS[3][8] ,
         \REGISTERS[3][7] , \REGISTERS[3][6] , \REGISTERS[3][5] ,
         \REGISTERS[3][4] , \REGISTERS[3][3] , \REGISTERS[3][2] ,
         \REGISTERS[3][1] , \REGISTERS[3][0] , \REGISTERS[4][31] ,
         \REGISTERS[4][30] , \REGISTERS[4][29] , \REGISTERS[4][28] ,
         \REGISTERS[4][27] , \REGISTERS[4][26] , \REGISTERS[4][25] ,
         \REGISTERS[4][24] , \REGISTERS[4][23] , \REGISTERS[4][22] ,
         \REGISTERS[4][21] , \REGISTERS[4][20] , \REGISTERS[4][19] ,
         \REGISTERS[4][18] , \REGISTERS[4][17] , \REGISTERS[4][16] ,
         \REGISTERS[4][15] , \REGISTERS[4][14] , \REGISTERS[4][13] ,
         \REGISTERS[4][12] , \REGISTERS[4][11] , \REGISTERS[4][10] ,
         \REGISTERS[4][9] , \REGISTERS[4][8] , \REGISTERS[4][7] ,
         \REGISTERS[4][6] , \REGISTERS[4][5] , \REGISTERS[4][4] ,
         \REGISTERS[4][3] , \REGISTERS[4][2] , \REGISTERS[4][1] ,
         \REGISTERS[4][0] , \REGISTERS[5][31] , \REGISTERS[5][30] ,
         \REGISTERS[5][29] , \REGISTERS[5][28] , \REGISTERS[5][27] ,
         \REGISTERS[5][26] , \REGISTERS[5][25] , \REGISTERS[5][24] ,
         \REGISTERS[5][23] , \REGISTERS[5][22] , \REGISTERS[5][21] ,
         \REGISTERS[5][20] , \REGISTERS[5][19] , \REGISTERS[5][18] ,
         \REGISTERS[5][17] , \REGISTERS[5][16] , \REGISTERS[5][15] ,
         \REGISTERS[5][14] , \REGISTERS[5][13] , \REGISTERS[5][12] ,
         \REGISTERS[5][11] , \REGISTERS[5][10] , \REGISTERS[5][9] ,
         \REGISTERS[5][8] , \REGISTERS[5][7] , \REGISTERS[5][6] ,
         \REGISTERS[5][5] , \REGISTERS[5][4] , \REGISTERS[5][3] ,
         \REGISTERS[5][2] , \REGISTERS[5][1] , \REGISTERS[5][0] ,
         \REGISTERS[6][31] , \REGISTERS[6][30] , \REGISTERS[6][29] ,
         \REGISTERS[6][28] , \REGISTERS[6][27] , \REGISTERS[6][26] ,
         \REGISTERS[6][25] , \REGISTERS[6][24] , \REGISTERS[6][23] ,
         \REGISTERS[6][22] , \REGISTERS[6][21] , \REGISTERS[6][20] ,
         \REGISTERS[6][19] , \REGISTERS[6][18] , \REGISTERS[6][17] ,
         \REGISTERS[6][16] , \REGISTERS[6][15] , \REGISTERS[6][14] ,
         \REGISTERS[6][13] , \REGISTERS[6][12] , \REGISTERS[6][11] ,
         \REGISTERS[6][10] , \REGISTERS[6][9] , \REGISTERS[6][8] ,
         \REGISTERS[6][7] , \REGISTERS[6][6] , \REGISTERS[6][5] ,
         \REGISTERS[6][4] , \REGISTERS[6][3] , \REGISTERS[6][2] ,
         \REGISTERS[6][1] , \REGISTERS[6][0] , \REGISTERS[7][31] ,
         \REGISTERS[7][30] , \REGISTERS[7][29] , \REGISTERS[7][28] ,
         \REGISTERS[7][27] , \REGISTERS[7][26] , \REGISTERS[7][25] ,
         \REGISTERS[7][24] , \REGISTERS[7][23] , \REGISTERS[7][22] ,
         \REGISTERS[7][21] , \REGISTERS[7][20] , \REGISTERS[7][19] ,
         \REGISTERS[7][18] , \REGISTERS[7][17] , \REGISTERS[7][16] ,
         \REGISTERS[7][15] , \REGISTERS[7][14] , \REGISTERS[7][13] ,
         \REGISTERS[7][12] , \REGISTERS[7][11] , \REGISTERS[7][10] ,
         \REGISTERS[7][9] , \REGISTERS[7][8] , \REGISTERS[7][7] ,
         \REGISTERS[7][6] , \REGISTERS[7][5] , \REGISTERS[7][4] ,
         \REGISTERS[7][3] , \REGISTERS[7][2] , \REGISTERS[7][1] ,
         \REGISTERS[7][0] , \REGISTERS[8][31] , \REGISTERS[8][30] ,
         \REGISTERS[8][29] , \REGISTERS[8][28] , \REGISTERS[8][27] ,
         \REGISTERS[8][26] , \REGISTERS[8][25] , \REGISTERS[8][24] ,
         \REGISTERS[8][23] , \REGISTERS[8][22] , \REGISTERS[8][21] ,
         \REGISTERS[8][20] , \REGISTERS[8][19] , \REGISTERS[8][18] ,
         \REGISTERS[8][17] , \REGISTERS[8][16] , \REGISTERS[8][15] ,
         \REGISTERS[8][14] , \REGISTERS[8][13] , \REGISTERS[8][12] ,
         \REGISTERS[8][11] , \REGISTERS[8][10] , \REGISTERS[8][9] ,
         \REGISTERS[8][8] , \REGISTERS[8][7] , \REGISTERS[8][6] ,
         \REGISTERS[8][5] , \REGISTERS[8][4] , \REGISTERS[8][3] ,
         \REGISTERS[8][2] , \REGISTERS[8][1] , \REGISTERS[8][0] ,
         \REGISTERS[9][31] , \REGISTERS[9][30] , \REGISTERS[9][29] ,
         \REGISTERS[9][28] , \REGISTERS[9][27] , \REGISTERS[9][26] ,
         \REGISTERS[9][25] , \REGISTERS[9][24] , \REGISTERS[9][23] ,
         \REGISTERS[9][22] , \REGISTERS[9][21] , \REGISTERS[9][20] ,
         \REGISTERS[9][19] , \REGISTERS[9][18] , \REGISTERS[9][17] ,
         \REGISTERS[9][16] , \REGISTERS[9][15] , \REGISTERS[9][14] ,
         \REGISTERS[9][13] , \REGISTERS[9][12] , \REGISTERS[9][11] ,
         \REGISTERS[9][10] , \REGISTERS[9][9] , \REGISTERS[9][8] ,
         \REGISTERS[9][7] , \REGISTERS[9][6] , \REGISTERS[9][5] ,
         \REGISTERS[9][4] , \REGISTERS[9][3] , \REGISTERS[9][2] ,
         \REGISTERS[9][1] , \REGISTERS[9][0] , \REGISTERS[10][31] ,
         \REGISTERS[10][30] , \REGISTERS[10][29] , \REGISTERS[10][28] ,
         \REGISTERS[10][27] , \REGISTERS[10][26] , \REGISTERS[10][25] ,
         \REGISTERS[10][24] , \REGISTERS[10][23] , \REGISTERS[10][22] ,
         \REGISTERS[10][21] , \REGISTERS[10][20] , \REGISTERS[10][19] ,
         \REGISTERS[10][18] , \REGISTERS[10][17] , \REGISTERS[10][16] ,
         \REGISTERS[10][15] , \REGISTERS[10][14] , \REGISTERS[10][13] ,
         \REGISTERS[10][12] , \REGISTERS[10][11] , \REGISTERS[10][10] ,
         \REGISTERS[10][9] , \REGISTERS[10][8] , \REGISTERS[10][7] ,
         \REGISTERS[10][6] , \REGISTERS[10][5] , \REGISTERS[10][4] ,
         \REGISTERS[10][3] , \REGISTERS[10][2] , \REGISTERS[10][1] ,
         \REGISTERS[10][0] , \REGISTERS[11][31] , \REGISTERS[11][30] ,
         \REGISTERS[11][29] , \REGISTERS[11][28] , \REGISTERS[11][27] ,
         \REGISTERS[11][26] , \REGISTERS[11][25] , \REGISTERS[11][24] ,
         \REGISTERS[11][23] , \REGISTERS[11][22] , \REGISTERS[11][21] ,
         \REGISTERS[11][20] , \REGISTERS[11][19] , \REGISTERS[11][18] ,
         \REGISTERS[11][17] , \REGISTERS[11][16] , \REGISTERS[11][15] ,
         \REGISTERS[11][14] , \REGISTERS[11][13] , \REGISTERS[11][12] ,
         \REGISTERS[11][11] , \REGISTERS[11][10] , \REGISTERS[11][9] ,
         \REGISTERS[11][8] , \REGISTERS[11][7] , \REGISTERS[11][6] ,
         \REGISTERS[11][5] , \REGISTERS[11][4] , \REGISTERS[11][3] ,
         \REGISTERS[11][2] , \REGISTERS[11][1] , \REGISTERS[11][0] ,
         \REGISTERS[12][31] , \REGISTERS[12][30] , \REGISTERS[12][29] ,
         \REGISTERS[12][28] , \REGISTERS[12][27] , \REGISTERS[12][26] ,
         \REGISTERS[12][25] , \REGISTERS[12][24] , \REGISTERS[12][23] ,
         \REGISTERS[12][22] , \REGISTERS[12][21] , \REGISTERS[12][20] ,
         \REGISTERS[12][19] , \REGISTERS[12][18] , \REGISTERS[12][17] ,
         \REGISTERS[12][16] , \REGISTERS[12][15] , \REGISTERS[12][14] ,
         \REGISTERS[12][13] , \REGISTERS[12][12] , \REGISTERS[12][11] ,
         \REGISTERS[12][10] , \REGISTERS[12][9] , \REGISTERS[12][8] ,
         \REGISTERS[12][7] , \REGISTERS[12][6] , \REGISTERS[12][5] ,
         \REGISTERS[12][4] , \REGISTERS[12][3] , \REGISTERS[12][2] ,
         \REGISTERS[12][1] , \REGISTERS[12][0] , \REGISTERS[13][31] ,
         \REGISTERS[13][30] , \REGISTERS[13][29] , \REGISTERS[13][28] ,
         \REGISTERS[13][27] , \REGISTERS[13][26] , \REGISTERS[13][25] ,
         \REGISTERS[13][24] , \REGISTERS[13][23] , \REGISTERS[13][22] ,
         \REGISTERS[13][21] , \REGISTERS[13][20] , \REGISTERS[13][19] ,
         \REGISTERS[13][18] , \REGISTERS[13][17] , \REGISTERS[13][16] ,
         \REGISTERS[13][15] , \REGISTERS[13][14] , \REGISTERS[13][13] ,
         \REGISTERS[13][12] , \REGISTERS[13][11] , \REGISTERS[13][10] ,
         \REGISTERS[13][9] , \REGISTERS[13][8] , \REGISTERS[13][7] ,
         \REGISTERS[13][6] , \REGISTERS[13][5] , \REGISTERS[13][4] ,
         \REGISTERS[13][3] , \REGISTERS[13][2] , \REGISTERS[13][1] ,
         \REGISTERS[13][0] , \REGISTERS[14][31] , \REGISTERS[14][30] ,
         \REGISTERS[14][29] , \REGISTERS[14][28] , \REGISTERS[14][27] ,
         \REGISTERS[14][26] , \REGISTERS[14][25] , \REGISTERS[14][24] ,
         \REGISTERS[14][23] , \REGISTERS[14][22] , \REGISTERS[14][21] ,
         \REGISTERS[14][20] , \REGISTERS[14][19] , \REGISTERS[14][18] ,
         \REGISTERS[14][17] , \REGISTERS[14][16] , \REGISTERS[14][15] ,
         \REGISTERS[14][14] , \REGISTERS[14][13] , \REGISTERS[14][12] ,
         \REGISTERS[14][11] , \REGISTERS[14][10] , \REGISTERS[14][9] ,
         \REGISTERS[14][8] , \REGISTERS[14][7] , \REGISTERS[14][6] ,
         \REGISTERS[14][5] , \REGISTERS[14][4] , \REGISTERS[14][3] ,
         \REGISTERS[14][2] , \REGISTERS[14][1] , \REGISTERS[14][0] ,
         \REGISTERS[15][31] , \REGISTERS[15][30] , \REGISTERS[15][29] ,
         \REGISTERS[15][28] , \REGISTERS[15][27] , \REGISTERS[15][26] ,
         \REGISTERS[15][25] , \REGISTERS[15][24] , \REGISTERS[15][23] ,
         \REGISTERS[15][22] , \REGISTERS[15][21] , \REGISTERS[15][20] ,
         \REGISTERS[15][19] , \REGISTERS[15][18] , \REGISTERS[15][17] ,
         \REGISTERS[15][16] , \REGISTERS[15][15] , \REGISTERS[15][14] ,
         \REGISTERS[15][13] , \REGISTERS[15][12] , \REGISTERS[15][11] ,
         \REGISTERS[15][10] , \REGISTERS[15][9] , \REGISTERS[15][8] ,
         \REGISTERS[15][7] , \REGISTERS[15][6] , \REGISTERS[15][5] ,
         \REGISTERS[15][4] , \REGISTERS[15][3] , \REGISTERS[15][2] ,
         \REGISTERS[15][1] , \REGISTERS[15][0] , \REGISTERS[16][31] ,
         \REGISTERS[16][30] , \REGISTERS[16][29] , \REGISTERS[16][28] ,
         \REGISTERS[16][27] , \REGISTERS[16][26] , \REGISTERS[16][25] ,
         \REGISTERS[16][24] , \REGISTERS[16][23] , \REGISTERS[16][22] ,
         \REGISTERS[16][21] , \REGISTERS[16][20] , \REGISTERS[16][19] ,
         \REGISTERS[16][18] , \REGISTERS[16][17] , \REGISTERS[16][16] ,
         \REGISTERS[16][15] , \REGISTERS[16][14] , \REGISTERS[16][13] ,
         \REGISTERS[16][12] , \REGISTERS[16][11] , \REGISTERS[16][10] ,
         \REGISTERS[16][9] , \REGISTERS[16][8] , \REGISTERS[16][7] ,
         \REGISTERS[16][6] , \REGISTERS[16][5] , \REGISTERS[16][4] ,
         \REGISTERS[16][3] , \REGISTERS[16][2] , \REGISTERS[16][1] ,
         \REGISTERS[16][0] , \REGISTERS[17][31] , \REGISTERS[17][30] ,
         \REGISTERS[17][29] , \REGISTERS[17][28] , \REGISTERS[17][27] ,
         \REGISTERS[17][26] , \REGISTERS[17][25] , \REGISTERS[17][24] ,
         \REGISTERS[17][23] , \REGISTERS[17][22] , \REGISTERS[17][21] ,
         \REGISTERS[17][20] , \REGISTERS[17][19] , \REGISTERS[17][18] ,
         \REGISTERS[17][17] , \REGISTERS[17][16] , \REGISTERS[17][15] ,
         \REGISTERS[17][14] , \REGISTERS[17][13] , \REGISTERS[17][12] ,
         \REGISTERS[17][11] , \REGISTERS[17][10] , \REGISTERS[17][9] ,
         \REGISTERS[17][8] , \REGISTERS[17][7] , \REGISTERS[17][6] ,
         \REGISTERS[17][5] , \REGISTERS[17][4] , \REGISTERS[17][3] ,
         \REGISTERS[17][2] , \REGISTERS[17][1] , \REGISTERS[17][0] ,
         \REGISTERS[18][31] , \REGISTERS[18][30] , \REGISTERS[18][29] ,
         \REGISTERS[18][28] , \REGISTERS[18][27] , \REGISTERS[18][26] ,
         \REGISTERS[18][25] , \REGISTERS[18][24] , \REGISTERS[18][23] ,
         \REGISTERS[18][22] , \REGISTERS[18][21] , \REGISTERS[18][20] ,
         \REGISTERS[18][19] , \REGISTERS[18][18] , \REGISTERS[18][17] ,
         \REGISTERS[18][16] , \REGISTERS[18][15] , \REGISTERS[18][14] ,
         \REGISTERS[18][13] , \REGISTERS[18][12] , \REGISTERS[18][11] ,
         \REGISTERS[18][10] , \REGISTERS[18][9] , \REGISTERS[18][8] ,
         \REGISTERS[18][7] , \REGISTERS[18][6] , \REGISTERS[18][5] ,
         \REGISTERS[18][4] , \REGISTERS[18][3] , \REGISTERS[18][2] ,
         \REGISTERS[18][1] , \REGISTERS[18][0] , \REGISTERS[19][31] ,
         \REGISTERS[19][30] , \REGISTERS[19][29] , \REGISTERS[19][28] ,
         \REGISTERS[19][27] , \REGISTERS[19][26] , \REGISTERS[19][25] ,
         \REGISTERS[19][24] , \REGISTERS[19][23] , \REGISTERS[19][22] ,
         \REGISTERS[19][21] , \REGISTERS[19][20] , \REGISTERS[19][19] ,
         \REGISTERS[19][18] , \REGISTERS[19][17] , \REGISTERS[19][16] ,
         \REGISTERS[19][15] , \REGISTERS[19][14] , \REGISTERS[19][13] ,
         \REGISTERS[19][12] , \REGISTERS[19][11] , \REGISTERS[19][10] ,
         \REGISTERS[19][9] , \REGISTERS[19][8] , \REGISTERS[19][7] ,
         \REGISTERS[19][6] , \REGISTERS[19][5] , \REGISTERS[19][4] ,
         \REGISTERS[19][3] , \REGISTERS[19][2] , \REGISTERS[19][1] ,
         \REGISTERS[19][0] , \REGISTERS[20][31] , \REGISTERS[20][30] ,
         \REGISTERS[20][29] , \REGISTERS[20][28] , \REGISTERS[20][27] ,
         \REGISTERS[20][26] , \REGISTERS[20][25] , \REGISTERS[20][24] ,
         \REGISTERS[20][23] , \REGISTERS[20][22] , \REGISTERS[20][21] ,
         \REGISTERS[20][20] , \REGISTERS[20][19] , \REGISTERS[20][18] ,
         \REGISTERS[20][17] , \REGISTERS[20][16] , \REGISTERS[20][15] ,
         \REGISTERS[20][14] , \REGISTERS[20][13] , \REGISTERS[20][12] ,
         \REGISTERS[20][11] , \REGISTERS[20][10] , \REGISTERS[20][9] ,
         \REGISTERS[20][8] , \REGISTERS[20][7] , \REGISTERS[20][6] ,
         \REGISTERS[20][5] , \REGISTERS[20][4] , \REGISTERS[20][3] ,
         \REGISTERS[20][2] , \REGISTERS[20][1] , \REGISTERS[20][0] ,
         \REGISTERS[21][31] , \REGISTERS[21][30] , \REGISTERS[21][29] ,
         \REGISTERS[21][28] , \REGISTERS[21][27] , \REGISTERS[21][26] ,
         \REGISTERS[21][25] , \REGISTERS[21][24] , \REGISTERS[21][23] ,
         \REGISTERS[21][22] , \REGISTERS[21][21] , \REGISTERS[21][20] ,
         \REGISTERS[21][19] , \REGISTERS[21][18] , \REGISTERS[21][17] ,
         \REGISTERS[21][16] , \REGISTERS[21][15] , \REGISTERS[21][14] ,
         \REGISTERS[21][13] , \REGISTERS[21][12] , \REGISTERS[21][11] ,
         \REGISTERS[21][10] , \REGISTERS[21][9] , \REGISTERS[21][8] ,
         \REGISTERS[21][7] , \REGISTERS[21][6] , \REGISTERS[21][5] ,
         \REGISTERS[21][4] , \REGISTERS[21][3] , \REGISTERS[21][2] ,
         \REGISTERS[21][1] , \REGISTERS[21][0] , \REGISTERS[22][31] ,
         \REGISTERS[22][30] , \REGISTERS[22][29] , \REGISTERS[22][28] ,
         \REGISTERS[22][27] , \REGISTERS[22][26] , \REGISTERS[22][25] ,
         \REGISTERS[22][24] , \REGISTERS[22][23] , \REGISTERS[22][22] ,
         \REGISTERS[22][21] , \REGISTERS[22][20] , \REGISTERS[22][19] ,
         \REGISTERS[22][18] , \REGISTERS[22][17] , \REGISTERS[22][16] ,
         \REGISTERS[22][15] , \REGISTERS[22][14] , \REGISTERS[22][13] ,
         \REGISTERS[22][12] , \REGISTERS[22][11] , \REGISTERS[22][10] ,
         \REGISTERS[22][9] , \REGISTERS[22][8] , \REGISTERS[22][7] ,
         \REGISTERS[22][6] , \REGISTERS[22][5] , \REGISTERS[22][4] ,
         \REGISTERS[22][3] , \REGISTERS[22][2] , \REGISTERS[22][1] ,
         \REGISTERS[22][0] , \REGISTERS[23][31] , \REGISTERS[23][30] ,
         \REGISTERS[23][29] , \REGISTERS[23][28] , \REGISTERS[23][27] ,
         \REGISTERS[23][26] , \REGISTERS[23][25] , \REGISTERS[23][24] ,
         \REGISTERS[23][23] , \REGISTERS[23][22] , \REGISTERS[23][21] ,
         \REGISTERS[23][20] , \REGISTERS[23][19] , \REGISTERS[23][18] ,
         \REGISTERS[23][17] , \REGISTERS[23][16] , \REGISTERS[23][15] ,
         \REGISTERS[23][14] , \REGISTERS[23][13] , \REGISTERS[23][12] ,
         \REGISTERS[23][11] , \REGISTERS[23][10] , \REGISTERS[23][9] ,
         \REGISTERS[23][8] , \REGISTERS[23][7] , \REGISTERS[23][6] ,
         \REGISTERS[23][5] , \REGISTERS[23][4] , \REGISTERS[23][3] ,
         \REGISTERS[23][2] , \REGISTERS[23][1] , \REGISTERS[23][0] ,
         \REGISTERS[24][31] , \REGISTERS[24][30] , \REGISTERS[24][29] ,
         \REGISTERS[24][28] , \REGISTERS[24][27] , \REGISTERS[24][26] ,
         \REGISTERS[24][25] , \REGISTERS[24][24] , \REGISTERS[24][23] ,
         \REGISTERS[24][22] , \REGISTERS[24][21] , \REGISTERS[24][20] ,
         \REGISTERS[24][19] , \REGISTERS[24][18] , \REGISTERS[24][17] ,
         \REGISTERS[24][16] , \REGISTERS[24][15] , \REGISTERS[24][14] ,
         \REGISTERS[24][13] , \REGISTERS[24][12] , \REGISTERS[24][11] ,
         \REGISTERS[24][10] , \REGISTERS[24][9] , \REGISTERS[24][8] ,
         \REGISTERS[24][7] , \REGISTERS[24][6] , \REGISTERS[24][5] ,
         \REGISTERS[24][4] , \REGISTERS[24][3] , \REGISTERS[24][2] ,
         \REGISTERS[24][1] , \REGISTERS[24][0] , \REGISTERS[25][31] ,
         \REGISTERS[25][30] , \REGISTERS[25][29] , \REGISTERS[25][28] ,
         \REGISTERS[25][27] , \REGISTERS[25][26] , \REGISTERS[25][25] ,
         \REGISTERS[25][24] , \REGISTERS[25][23] , \REGISTERS[25][22] ,
         \REGISTERS[25][21] , \REGISTERS[25][20] , \REGISTERS[25][19] ,
         \REGISTERS[25][18] , \REGISTERS[25][17] , \REGISTERS[25][16] ,
         \REGISTERS[25][15] , \REGISTERS[25][14] , \REGISTERS[25][13] ,
         \REGISTERS[25][12] , \REGISTERS[25][11] , \REGISTERS[25][10] ,
         \REGISTERS[25][9] , \REGISTERS[25][8] , \REGISTERS[25][7] ,
         \REGISTERS[25][6] , \REGISTERS[25][5] , \REGISTERS[25][4] ,
         \REGISTERS[25][3] , \REGISTERS[25][2] , \REGISTERS[25][1] ,
         \REGISTERS[25][0] , \REGISTERS[26][31] , \REGISTERS[26][30] ,
         \REGISTERS[26][29] , \REGISTERS[26][28] , \REGISTERS[26][27] ,
         \REGISTERS[26][26] , \REGISTERS[26][25] , \REGISTERS[26][24] ,
         \REGISTERS[26][23] , \REGISTERS[26][22] , \REGISTERS[26][21] ,
         \REGISTERS[26][20] , \REGISTERS[26][19] , \REGISTERS[26][18] ,
         \REGISTERS[26][17] , \REGISTERS[26][16] , \REGISTERS[26][15] ,
         \REGISTERS[26][14] , \REGISTERS[26][13] , \REGISTERS[26][12] ,
         \REGISTERS[26][11] , \REGISTERS[26][10] , \REGISTERS[26][9] ,
         \REGISTERS[26][8] , \REGISTERS[26][7] , \REGISTERS[26][6] ,
         \REGISTERS[26][5] , \REGISTERS[26][4] , \REGISTERS[26][3] ,
         \REGISTERS[26][2] , \REGISTERS[26][1] , \REGISTERS[26][0] ,
         \REGISTERS[27][31] , \REGISTERS[27][30] , \REGISTERS[27][29] ,
         \REGISTERS[27][28] , \REGISTERS[27][27] , \REGISTERS[27][26] ,
         \REGISTERS[27][25] , \REGISTERS[27][24] , \REGISTERS[27][23] ,
         \REGISTERS[27][22] , \REGISTERS[27][21] , \REGISTERS[27][20] ,
         \REGISTERS[27][19] , \REGISTERS[27][18] , \REGISTERS[27][17] ,
         \REGISTERS[27][16] , \REGISTERS[27][15] , \REGISTERS[27][14] ,
         \REGISTERS[27][13] , \REGISTERS[27][12] , \REGISTERS[27][11] ,
         \REGISTERS[27][10] , \REGISTERS[27][9] , \REGISTERS[27][8] ,
         \REGISTERS[27][7] , \REGISTERS[27][6] , \REGISTERS[27][5] ,
         \REGISTERS[27][4] , \REGISTERS[27][3] , \REGISTERS[27][2] ,
         \REGISTERS[27][1] , \REGISTERS[27][0] , \REGISTERS[28][31] ,
         \REGISTERS[28][30] , \REGISTERS[28][29] , \REGISTERS[28][28] ,
         \REGISTERS[28][27] , \REGISTERS[28][26] , \REGISTERS[28][25] ,
         \REGISTERS[28][24] , \REGISTERS[28][23] , \REGISTERS[28][22] ,
         \REGISTERS[28][21] , \REGISTERS[28][20] , \REGISTERS[28][19] ,
         \REGISTERS[28][18] , \REGISTERS[28][17] , \REGISTERS[28][16] ,
         \REGISTERS[28][15] , \REGISTERS[28][14] , \REGISTERS[28][13] ,
         \REGISTERS[28][12] , \REGISTERS[28][11] , \REGISTERS[28][10] ,
         \REGISTERS[28][9] , \REGISTERS[28][8] , \REGISTERS[28][7] ,
         \REGISTERS[28][6] , \REGISTERS[28][5] , \REGISTERS[28][4] ,
         \REGISTERS[28][3] , \REGISTERS[28][2] , \REGISTERS[28][1] ,
         \REGISTERS[28][0] , \REGISTERS[29][31] , \REGISTERS[29][30] ,
         \REGISTERS[29][29] , \REGISTERS[29][28] , \REGISTERS[29][27] ,
         \REGISTERS[29][26] , \REGISTERS[29][25] , \REGISTERS[29][24] ,
         \REGISTERS[29][23] , \REGISTERS[29][22] , \REGISTERS[29][21] ,
         \REGISTERS[29][20] , \REGISTERS[29][19] , \REGISTERS[29][18] ,
         \REGISTERS[29][17] , \REGISTERS[29][16] , \REGISTERS[29][15] ,
         \REGISTERS[29][14] , \REGISTERS[29][13] , \REGISTERS[29][12] ,
         \REGISTERS[29][11] , \REGISTERS[29][10] , \REGISTERS[29][9] ,
         \REGISTERS[29][8] , \REGISTERS[29][7] , \REGISTERS[29][6] ,
         \REGISTERS[29][5] , \REGISTERS[29][4] , \REGISTERS[29][3] ,
         \REGISTERS[29][2] , \REGISTERS[29][1] , \REGISTERS[29][0] ,
         \REGISTERS[30][31] , \REGISTERS[30][30] , \REGISTERS[30][29] ,
         \REGISTERS[30][28] , \REGISTERS[30][27] , \REGISTERS[30][26] ,
         \REGISTERS[30][25] , \REGISTERS[30][24] , \REGISTERS[30][23] ,
         \REGISTERS[30][22] , \REGISTERS[30][21] , \REGISTERS[30][20] ,
         \REGISTERS[30][19] , \REGISTERS[30][18] , \REGISTERS[30][17] ,
         \REGISTERS[30][16] , \REGISTERS[30][15] , \REGISTERS[30][14] ,
         \REGISTERS[30][13] , \REGISTERS[30][12] , \REGISTERS[30][11] ,
         \REGISTERS[30][10] , \REGISTERS[30][9] , \REGISTERS[30][8] ,
         \REGISTERS[30][7] , \REGISTERS[30][6] , \REGISTERS[30][5] ,
         \REGISTERS[30][4] , \REGISTERS[30][3] , \REGISTERS[30][2] ,
         \REGISTERS[30][1] , \REGISTERS[30][0] , \REGISTERS[31][31] ,
         \REGISTERS[31][30] , \REGISTERS[31][29] , \REGISTERS[31][28] ,
         \REGISTERS[31][27] , \REGISTERS[31][26] , \REGISTERS[31][25] ,
         \REGISTERS[31][24] , \REGISTERS[31][23] , \REGISTERS[31][22] ,
         \REGISTERS[31][21] , \REGISTERS[31][20] , \REGISTERS[31][19] ,
         \REGISTERS[31][18] , \REGISTERS[31][17] , \REGISTERS[31][16] ,
         \REGISTERS[31][15] , \REGISTERS[31][14] , \REGISTERS[31][13] ,
         \REGISTERS[31][12] , \REGISTERS[31][11] , \REGISTERS[31][10] ,
         \REGISTERS[31][9] , \REGISTERS[31][8] , \REGISTERS[31][7] ,
         \REGISTERS[31][6] , \REGISTERS[31][5] , \REGISTERS[31][4] ,
         \REGISTERS[31][3] , \REGISTERS[31][2] , \REGISTERS[31][1] ,
         \REGISTERS[31][0] , N81, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, net7104, net7110, net7115, net7120, net7125, net7130,
         net7135, net7140, net7145, net7150, net7155, net7160, net7165,
         net7170, net7175, net7180, net7185, net7190, net7195, net7200,
         net7205, net7210, net7215, net7220, net7225, net7230, net7235,
         net7240, net7245, net7250, net7255, net7260, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77,
         n78, n80, n81, n82, n83, n84, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n116, n117, n118,
         n119, n120, n121, n122, n124, n125, n126, n127, n128, n129, n130,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1810, n1811, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695;

  DLH_X1 \OUT1_reg[31]  ( .G(N411), .D(N278), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(N411), .D(N277), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(N411), .D(N276), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(N411), .D(N275), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(N411), .D(N274), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(N411), .D(N273), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(N411), .D(N272), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(N411), .D(N271), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(N411), .D(N270), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(N411), .D(N269), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(N411), .D(N268), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(N411), .D(N267), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(N411), .D(N266), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(N411), .D(N265), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(N411), .D(N264), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(N411), .D(N263), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(N411), .D(N262), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(N411), .D(N261), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(N411), .D(N260), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(N411), .D(N259), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(N411), .D(N258), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(N411), .D(N257), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(N411), .D(N256), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(N411), .D(N255), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(N411), .D(N254), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(N411), .D(N253), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(N411), .D(N252), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(N411), .D(N251), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(N411), .D(N250), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(N411), .D(N249), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(N411), .D(N248), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(N411), .D(N247), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(N412), .D(N410), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(N412), .D(N409), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(N412), .D(N408), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(N412), .D(N407), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(N412), .D(N406), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(N412), .D(N405), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(N412), .D(N404), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(N412), .D(N403), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(N412), .D(N402), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(N412), .D(N401), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(N412), .D(N400), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(N412), .D(N399), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(N412), .D(N398), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(N412), .D(N397), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(N412), .D(N396), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(N412), .D(N395), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(N412), .D(N394), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(N412), .D(N393), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(N412), .D(N392), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(N412), .D(N391), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(N412), .D(N390), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(N412), .D(N389), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(N412), .D(N388), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(N412), .D(N387), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(N412), .D(N386), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(N412), .D(N385), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(N412), .D(N384), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(N412), .D(N383), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(N412), .D(N382), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(N412), .D(N381), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(N412), .D(N380), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(N412), .D(N379), .Q(OUT2[0]) );
  INV_X1 U40 ( .A(n120), .ZN(n119) );
  INV_X1 U42 ( .A(n122), .ZN(n121) );
  AND2_X1 U54 ( .A1(n1806), .A2(RD1), .ZN(N411) );
  AND2_X1 U55 ( .A1(n1806), .A2(RD2), .ZN(N412) );
  INV_X1 U56 ( .A(DATAIN[6]), .ZN(n124) );
  INV_X1 U57 ( .A(DATAIN[14]), .ZN(n108) );
  INV_X1 U58 ( .A(DATAIN[26]), .ZN(n84) );
  INV_X1 U59 ( .A(DATAIN[18]), .ZN(n100) );
  INV_X1 U60 ( .A(DATAIN[22]), .ZN(n92) );
  INV_X1 U61 ( .A(n71), .ZN(n69) );
  BUF_X1 U62 ( .A(n1575), .Z(n38) );
  BUF_X1 U63 ( .A(n1599), .Z(n54) );
  BUF_X1 U64 ( .A(n1577), .Z(n40) );
  BUF_X1 U65 ( .A(n1613), .Z(n64) );
  BUF_X1 U66 ( .A(n1579), .Z(n42) );
  BUF_X1 U67 ( .A(n1589), .Z(n48) );
  BUF_X1 U68 ( .A(n1601), .Z(n56) );
  BUF_X1 U69 ( .A(n1581), .Z(n44) );
  BUF_X1 U70 ( .A(n1617), .Z(n68) );
  BUF_X1 U71 ( .A(n1605), .Z(n60) );
  BUF_X1 U72 ( .A(n1615), .Z(n66) );
  BUF_X1 U73 ( .A(n72), .Z(n71) );
  BUF_X1 U74 ( .A(n1616), .Z(n67) );
  BUF_X1 U75 ( .A(n1614), .Z(n65) );
  BUF_X1 U76 ( .A(n1612), .Z(n63) );
  BUF_X1 U77 ( .A(n1610), .Z(n61) );
  BUF_X1 U78 ( .A(n1611), .Z(n62) );
  BUF_X1 U79 ( .A(n1604), .Z(n59) );
  BUF_X1 U80 ( .A(n1602), .Z(n57) );
  BUF_X1 U81 ( .A(n1603), .Z(n58) );
  BUF_X1 U82 ( .A(n1600), .Z(n55) );
  BUF_X1 U83 ( .A(n1598), .Z(n53) );
  BUF_X1 U84 ( .A(n1592), .Z(n51) );
  BUF_X1 U85 ( .A(n1593), .Z(n52) );
  BUF_X1 U86 ( .A(n1590), .Z(n49) );
  BUF_X1 U87 ( .A(n1591), .Z(n50) );
  BUF_X1 U88 ( .A(n1588), .Z(n47) );
  BUF_X1 U89 ( .A(n1586), .Z(n45) );
  BUF_X1 U90 ( .A(n1587), .Z(n46) );
  BUF_X1 U91 ( .A(n1580), .Z(n43) );
  BUF_X1 U92 ( .A(n1578), .Z(n41) );
  BUF_X1 U93 ( .A(n1576), .Z(n39) );
  BUF_X1 U94 ( .A(n1574), .Z(n37) );
  INV_X1 U95 ( .A(n72), .ZN(n70) );
  INV_X1 U96 ( .A(n1627), .ZN(n72) );
  NOR3_X1 U97 ( .A1(n903), .A2(n902), .A3(n901), .ZN(n1627) );
  INV_X1 U98 ( .A(ADD_RD2[4]), .ZN(n912) );
  INV_X1 U99 ( .A(DATAIN[2]), .ZN(n132) );
  INV_X1 U100 ( .A(n35), .ZN(n33) );
  BUF_X1 U101 ( .A(n843), .Z(n4) );
  BUF_X1 U102 ( .A(n878), .Z(n27) );
  BUF_X1 U103 ( .A(n845), .Z(n6) );
  BUF_X1 U104 ( .A(n866), .Z(n19) );
  BUF_X1 U105 ( .A(n880), .Z(n29) );
  BUF_X1 U106 ( .A(n868), .Z(n21) );
  BUF_X1 U107 ( .A(n865), .Z(n18) );
  INV_X1 U108 ( .A(DATAIN[9]), .ZN(n118) );
  BUF_X1 U109 ( .A(n36), .Z(n35) );
  BUF_X1 U110 ( .A(n856), .Z(n13) );
  BUF_X1 U111 ( .A(n846), .Z(n7) );
  BUF_X1 U112 ( .A(n842), .Z(n3) );
  BUF_X1 U113 ( .A(n844), .Z(n5) );
  BUF_X1 U114 ( .A(n867), .Z(n20) );
  BUF_X1 U115 ( .A(n858), .Z(n15) );
  BUF_X1 U116 ( .A(n877), .Z(n26) );
  BUF_X1 U117 ( .A(n876), .Z(n25) );
  BUF_X1 U118 ( .A(n883), .Z(n32) );
  BUF_X1 U119 ( .A(n847), .Z(n8) );
  BUF_X1 U120 ( .A(n859), .Z(n16) );
  BUF_X1 U121 ( .A(n871), .Z(n24) );
  BUF_X1 U122 ( .A(n882), .Z(n31) );
  BUF_X1 U123 ( .A(n869), .Z(n22) );
  BUF_X1 U124 ( .A(n870), .Z(n23) );
  BUF_X1 U125 ( .A(n853), .Z(n10) );
  BUF_X1 U126 ( .A(n879), .Z(n28) );
  BUF_X1 U127 ( .A(n855), .Z(n12) );
  BUF_X1 U128 ( .A(n881), .Z(n30) );
  BUF_X1 U129 ( .A(n841), .Z(n2) );
  BUF_X1 U130 ( .A(n852), .Z(n9) );
  BUF_X1 U131 ( .A(n864), .Z(n17) );
  BUF_X1 U132 ( .A(n840), .Z(n1) );
  BUF_X1 U133 ( .A(n854), .Z(n11) );
  BUF_X1 U134 ( .A(n857), .Z(n14) );
  INV_X1 U135 ( .A(n36), .ZN(n34) );
  INV_X1 U136 ( .A(n893), .ZN(n36) );
  NOR3_X1 U137 ( .A1(n170), .A2(n169), .A3(n168), .ZN(n893) );
  INV_X1 U138 ( .A(ADD_WR[0]), .ZN(n899) );
  INV_X1 U139 ( .A(ADD_WR[3]), .ZN(n897) );
  INV_X1 U140 ( .A(ADD_WR[4]), .ZN(n894) );
  INV_X1 U141 ( .A(ADD_WR[2]), .ZN(n900) );
  INV_X1 U142 ( .A(ADD_WR[1]), .ZN(n896) );
  INV_X1 U143 ( .A(n1639), .ZN(n134) );
  INV_X1 U144 ( .A(DATAIN[0]), .ZN(n136) );
  INV_X1 U145 ( .A(DATAIN[3]), .ZN(n130) );
  INV_X1 U146 ( .A(DATAIN[4]), .ZN(n128) );
  INV_X1 U147 ( .A(DATAIN[5]), .ZN(n126) );
  INV_X1 U148 ( .A(DATAIN[8]), .ZN(n120) );
  INV_X1 U149 ( .A(DATAIN[7]), .ZN(n122) );
  INV_X1 U150 ( .A(DATAIN[10]), .ZN(n116) );
  INV_X1 U151 ( .A(DATAIN[11]), .ZN(n114) );
  INV_X1 U152 ( .A(DATAIN[12]), .ZN(n112) );
  INV_X1 U153 ( .A(DATAIN[13]), .ZN(n110) );
  INV_X1 U154 ( .A(DATAIN[16]), .ZN(n104) );
  INV_X1 U155 ( .A(DATAIN[17]), .ZN(n102) );
  INV_X1 U156 ( .A(DATAIN[19]), .ZN(n98) );
  INV_X1 U157 ( .A(DATAIN[20]), .ZN(n96) );
  INV_X1 U158 ( .A(DATAIN[21]), .ZN(n94) );
  INV_X1 U159 ( .A(DATAIN[23]), .ZN(n90) );
  INV_X1 U160 ( .A(DATAIN[24]), .ZN(n88) );
  INV_X1 U161 ( .A(DATAIN[25]), .ZN(n86) );
  INV_X1 U162 ( .A(DATAIN[27]), .ZN(n82) );
  INV_X1 U163 ( .A(DATAIN[28]), .ZN(n80) );
  INV_X1 U164 ( .A(n1637), .ZN(n78) );
  INV_X1 U165 ( .A(DATAIN[30]), .ZN(n76) );
  INV_X1 U166 ( .A(DATAIN[31]), .ZN(n74) );
  INV_X1 U167 ( .A(DATAIN[15]), .ZN(n106) );
  NAND3_X1 U169 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n899), .ZN(n158) );
  OAI21_X1 U170 ( .B1(n1629), .B2(n158), .A(RST), .ZN(N114) );
  NAND3_X1 U171 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n896), .ZN(n159) );
  OAI21_X1 U172 ( .B1(n1629), .B2(n159), .A(RST), .ZN(N115) );
  NAND3_X1 U173 ( .A1(ADD_WR[2]), .A2(n899), .A3(n896), .ZN(n160) );
  OAI21_X1 U174 ( .B1(n1629), .B2(n160), .A(RST), .ZN(N116) );
  NAND3_X1 U175 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(n900), .ZN(n161) );
  OAI21_X1 U176 ( .B1(n1629), .B2(n161), .A(RST), .ZN(N117) );
  NAND3_X1 U177 ( .A1(ADD_WR[1]), .A2(n899), .A3(n900), .ZN(n162) );
  OAI21_X1 U178 ( .B1(n1629), .B2(n162), .A(RST), .ZN(N118) );
  NAND3_X1 U179 ( .A1(ADD_WR[0]), .A2(n896), .A3(n900), .ZN(n163) );
  OAI21_X1 U180 ( .B1(n1629), .B2(n163), .A(RST), .ZN(N119) );
  NAND3_X1 U181 ( .A1(n899), .A2(n896), .A3(n900), .ZN(n165) );
  OAI21_X1 U182 ( .B1(n1629), .B2(n165), .A(RST), .ZN(N120) );
  NAND3_X1 U183 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(ADD_WR[2]), .ZN(n1628)
         );
  OAI21_X1 U185 ( .B1(n1628), .B2(n156), .A(RST), .ZN(N121) );
  OAI21_X1 U186 ( .B1(n158), .B2(n156), .A(RST), .ZN(N122) );
  OAI21_X1 U187 ( .B1(n159), .B2(n156), .A(RST), .ZN(N123) );
  OAI21_X1 U188 ( .B1(n160), .B2(n156), .A(n145), .ZN(N124) );
  OAI21_X1 U189 ( .B1(n161), .B2(n156), .A(n155), .ZN(N125) );
  OAI21_X1 U190 ( .B1(n162), .B2(n156), .A(n141), .ZN(N126) );
  OAI21_X1 U191 ( .B1(n163), .B2(n156), .A(n138), .ZN(N127) );
  OAI21_X1 U192 ( .B1(n165), .B2(n156), .A(n140), .ZN(N128) );
  OAI21_X1 U194 ( .B1(n1628), .B2(n157), .A(n137), .ZN(N129) );
  OAI21_X1 U195 ( .B1(n158), .B2(n157), .A(n142), .ZN(N130) );
  OAI21_X1 U196 ( .B1(n159), .B2(n157), .A(n152), .ZN(N131) );
  OAI21_X1 U197 ( .B1(n160), .B2(n157), .A(n148), .ZN(N132) );
  OAI21_X1 U198 ( .B1(n161), .B2(n157), .A(n143), .ZN(N133) );
  OAI21_X1 U199 ( .B1(n162), .B2(n157), .A(n154), .ZN(N134) );
  OAI21_X1 U200 ( .B1(n163), .B2(n157), .A(n151), .ZN(N135) );
  OAI21_X1 U201 ( .B1(n165), .B2(n157), .A(RST), .ZN(N136) );
  OAI21_X1 U203 ( .B1(n1628), .B2(n164), .A(RST), .ZN(N137) );
  OAI21_X1 U204 ( .B1(n158), .B2(n164), .A(n145), .ZN(N138) );
  OAI21_X1 U205 ( .B1(n159), .B2(n164), .A(n155), .ZN(N139) );
  OAI21_X1 U206 ( .B1(n160), .B2(n164), .A(n147), .ZN(N140) );
  OAI21_X1 U207 ( .B1(n161), .B2(n164), .A(RST), .ZN(N141) );
  OAI21_X1 U208 ( .B1(n162), .B2(n164), .A(RST), .ZN(N142) );
  OAI21_X1 U209 ( .B1(n163), .B2(n164), .A(RST), .ZN(N143) );
  OAI21_X1 U210 ( .B1(n165), .B2(n164), .A(RST), .ZN(N144) );
  INV_X1 U211 ( .A(ADD_RD1[1]), .ZN(n172) );
  OAI221_X1 U212 ( .B1(ADD_WR[1]), .B2(n172), .C1(n896), .C2(ADD_RD1[1]), .A(
        WR), .ZN(n170) );
  AOI22_X1 U213 ( .A1(n900), .A2(ADD_RD1[2]), .B1(ADD_RD1[4]), .B2(n894), .ZN(
        n166) );
  OAI221_X1 U214 ( .B1(n900), .B2(ADD_RD1[2]), .C1(n894), .C2(ADD_RD1[4]), .A(
        n166), .ZN(n169) );
  AOI22_X1 U215 ( .A1(n897), .A2(ADD_RD1[3]), .B1(ADD_RD1[0]), .B2(n899), .ZN(
        n167) );
  OAI221_X1 U216 ( .B1(n897), .B2(ADD_RD1[3]), .C1(n899), .C2(ADD_RD1[0]), .A(
        n167), .ZN(n168) );
  NAND2_X1 U217 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n200) );
  INV_X1 U218 ( .A(ADD_RD1[3]), .ZN(n173) );
  INV_X1 U219 ( .A(ADD_RD1[4]), .ZN(n178) );
  NAND3_X1 U220 ( .A1(ADD_RD1[0]), .A2(n173), .A3(n178), .ZN(n193) );
  NOR2_X1 U221 ( .A1(n200), .A2(n193), .ZN(n877) );
  INV_X1 U222 ( .A(ADD_RD1[0]), .ZN(n179) );
  NAND3_X1 U223 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n179), .ZN(n185) );
  NOR2_X1 U224 ( .A1(n200), .A2(n185), .ZN(n879) );
  AOI22_X1 U225 ( .A1(\REGISTERS[7][0] ), .A2(n877), .B1(\REGISTERS[30][0] ), 
        .B2(n28), .ZN(n177) );
  INV_X1 U226 ( .A(ADD_RD1[2]), .ZN(n171) );
  NAND2_X1 U227 ( .A1(ADD_RD1[1]), .A2(n171), .ZN(n195) );
  NOR2_X1 U228 ( .A1(n185), .A2(n195), .ZN(n878) );
  NAND3_X1 U229 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n178), .ZN(n198) );
  NAND2_X1 U230 ( .A1(ADD_RD1[2]), .A2(n172), .ZN(n192) );
  NOR2_X1 U231 ( .A1(n198), .A2(n192), .ZN(n883) );
  AOI22_X1 U232 ( .A1(\REGISTERS[26][0] ), .A2(n878), .B1(\REGISTERS[13][0] ), 
        .B2(n32), .ZN(n176) );
  NAND2_X1 U233 ( .A1(n172), .A2(n171), .ZN(n197) );
  NAND3_X1 U234 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[0]), .A3(ADD_RD1[4]), .ZN(n199)
         );
  NOR2_X1 U235 ( .A1(n197), .A2(n199), .ZN(n881) );
  NOR2_X1 U236 ( .A1(n185), .A2(n192), .ZN(n855) );
  AOI22_X1 U237 ( .A1(\REGISTERS[25][0] ), .A2(n881), .B1(\REGISTERS[28][0] ), 
        .B2(n12), .ZN(n175) );
  NAND3_X1 U238 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n173), .ZN(n186) );
  NOR2_X1 U239 ( .A1(n197), .A2(n186), .ZN(n853) );
  NOR2_X1 U240 ( .A1(n192), .A2(n186), .ZN(n869) );
  AOI22_X1 U241 ( .A1(\REGISTERS[17][0] ), .A2(n853), .B1(\REGISTERS[21][0] ), 
        .B2(n22), .ZN(n174) );
  NAND4_X1 U242 ( .A1(n177), .A2(n176), .A3(n175), .A4(n174), .ZN(n208) );
  NOR2_X1 U243 ( .A1(n192), .A2(n199), .ZN(n857) );
  NOR2_X1 U244 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[0]), .ZN(n184) );
  NAND2_X1 U245 ( .A1(n184), .A2(n178), .ZN(n194) );
  NOR2_X1 U246 ( .A1(n200), .A2(n194), .ZN(n859) );
  AOI22_X1 U247 ( .A1(\REGISTERS[29][0] ), .A2(n857), .B1(\REGISTERS[6][0] ), 
        .B2(n16), .ZN(n183) );
  NAND3_X1 U248 ( .A1(ADD_RD1[3]), .A2(n179), .A3(n178), .ZN(n191) );
  NOR2_X1 U249 ( .A1(n195), .A2(n191), .ZN(n882) );
  NOR2_X1 U250 ( .A1(n197), .A2(n191), .ZN(n867) );
  AOI22_X1 U251 ( .A1(\REGISTERS[10][0] ), .A2(n882), .B1(\REGISTERS[8][0] ), 
        .B2(n20), .ZN(n182) );
  NOR2_X1 U252 ( .A1(n200), .A2(n198), .ZN(n876) );
  NOR2_X1 U253 ( .A1(n200), .A2(n191), .ZN(n865) );
  AOI22_X1 U254 ( .A1(\REGISTERS[15][0] ), .A2(n876), .B1(\REGISTERS[14][0] ), 
        .B2(n18), .ZN(n181) );
  NOR2_X1 U255 ( .A1(n200), .A2(n186), .ZN(n841) );
  NOR2_X1 U256 ( .A1(n197), .A2(n194), .ZN(n840) );
  AOI22_X1 U257 ( .A1(\REGISTERS[23][0] ), .A2(n841), .B1(\REGISTERS[0][0] ), 
        .B2(n1), .ZN(n180) );
  NAND4_X1 U258 ( .A1(n183), .A2(n182), .A3(n181), .A4(n180), .ZN(n207) );
  NOR2_X1 U259 ( .A1(n193), .A2(n197), .ZN(n847) );
  NAND2_X1 U260 ( .A1(ADD_RD1[4]), .A2(n184), .ZN(n196) );
  NOR2_X1 U261 ( .A1(n195), .A2(n196), .ZN(n868) );
  AOI22_X1 U262 ( .A1(\REGISTERS[1][0] ), .A2(n847), .B1(\REGISTERS[18][0] ), 
        .B2(n21), .ZN(n190) );
  NOR2_X1 U263 ( .A1(n195), .A2(n199), .ZN(n843) );
  NOR2_X1 U264 ( .A1(n192), .A2(n196), .ZN(n864) );
  AOI22_X1 U265 ( .A1(\REGISTERS[27][0] ), .A2(n843), .B1(\REGISTERS[20][0] ), 
        .B2(n864), .ZN(n189) );
  NOR2_X1 U266 ( .A1(n185), .A2(n197), .ZN(n845) );
  NOR2_X1 U267 ( .A1(n193), .A2(n195), .ZN(n854) );
  AOI22_X1 U268 ( .A1(\REGISTERS[24][0] ), .A2(n845), .B1(\REGISTERS[3][0] ), 
        .B2(n11), .ZN(n188) );
  NOR2_X1 U269 ( .A1(n195), .A2(n186), .ZN(n846) );
  NOR2_X1 U270 ( .A1(n192), .A2(n194), .ZN(n866) );
  AOI22_X1 U271 ( .A1(\REGISTERS[19][0] ), .A2(n846), .B1(\REGISTERS[4][0] ), 
        .B2(n866), .ZN(n187) );
  NAND4_X1 U272 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(n206) );
  NOR2_X1 U273 ( .A1(n192), .A2(n191), .ZN(n856) );
  NOR2_X1 U274 ( .A1(n193), .A2(n192), .ZN(n871) );
  AOI22_X1 U275 ( .A1(\REGISTERS[12][0] ), .A2(n856), .B1(\REGISTERS[5][0] ), 
        .B2(n24), .ZN(n204) );
  NOR2_X1 U276 ( .A1(n195), .A2(n194), .ZN(n842) );
  NOR2_X1 U277 ( .A1(n195), .A2(n198), .ZN(n880) );
  AOI22_X1 U278 ( .A1(\REGISTERS[2][0] ), .A2(n842), .B1(\REGISTERS[11][0] ), 
        .B2(n29), .ZN(n203) );
  NOR2_X1 U279 ( .A1(n200), .A2(n196), .ZN(n858) );
  NOR2_X1 U280 ( .A1(n197), .A2(n196), .ZN(n870) );
  AOI22_X1 U281 ( .A1(\REGISTERS[22][0] ), .A2(n858), .B1(\REGISTERS[16][0] ), 
        .B2(n870), .ZN(n202) );
  NOR2_X1 U282 ( .A1(n198), .A2(n197), .ZN(n852) );
  NOR2_X1 U283 ( .A1(n200), .A2(n199), .ZN(n844) );
  AOI22_X1 U284 ( .A1(\REGISTERS[9][0] ), .A2(n852), .B1(\REGISTERS[31][0] ), 
        .B2(n844), .ZN(n201) );
  NAND4_X1 U285 ( .A1(n204), .A2(n203), .A3(n202), .A4(n201), .ZN(n205) );
  NOR4_X1 U286 ( .A1(n208), .A2(n207), .A3(n206), .A4(n205), .ZN(n209) );
  AOI22_X1 U287 ( .A1(n33), .A2(n136), .B1(n209), .B2(n36), .ZN(N247) );
  AOI22_X1 U288 ( .A1(n841), .A2(\REGISTERS[23][1] ), .B1(n8), .B2(
        \REGISTERS[1][1] ), .ZN(n213) );
  AOI22_X1 U289 ( .A1(n27), .A2(\REGISTERS[26][1] ), .B1(n21), .B2(
        \REGISTERS[18][1] ), .ZN(n212) );
  AOI22_X1 U290 ( .A1(n854), .A2(\REGISTERS[3][1] ), .B1(n856), .B2(
        \REGISTERS[12][1] ), .ZN(n211) );
  AOI22_X1 U291 ( .A1(n867), .A2(\REGISTERS[8][1] ), .B1(n871), .B2(
        \REGISTERS[5][1] ), .ZN(n210) );
  NAND4_X1 U292 ( .A1(n213), .A2(n212), .A3(n211), .A4(n210), .ZN(n229) );
  AOI22_X1 U293 ( .A1(n882), .A2(\REGISTERS[10][1] ), .B1(n18), .B2(
        \REGISTERS[14][1] ), .ZN(n217) );
  AOI22_X1 U294 ( .A1(n12), .A2(\REGISTERS[28][1] ), .B1(n846), .B2(
        \REGISTERS[19][1] ), .ZN(n216) );
  AOI22_X1 U295 ( .A1(n859), .A2(\REGISTERS[6][1] ), .B1(n864), .B2(
        \REGISTERS[20][1] ), .ZN(n215) );
  AOI22_X1 U296 ( .A1(n866), .A2(\REGISTERS[4][1] ), .B1(n9), .B2(
        \REGISTERS[9][1] ), .ZN(n214) );
  NAND4_X1 U297 ( .A1(n217), .A2(n216), .A3(n215), .A4(n214), .ZN(n228) );
  AOI22_X1 U298 ( .A1(n30), .A2(\REGISTERS[25][1] ), .B1(n15), .B2(
        \REGISTERS[22][1] ), .ZN(n221) );
  AOI22_X1 U299 ( .A1(n869), .A2(\REGISTERS[21][1] ), .B1(n880), .B2(
        \REGISTERS[11][1] ), .ZN(n220) );
  AOI22_X1 U300 ( .A1(n3), .A2(\REGISTERS[2][1] ), .B1(n5), .B2(
        \REGISTERS[31][1] ), .ZN(n219) );
  AOI22_X1 U301 ( .A1(n26), .A2(\REGISTERS[7][1] ), .B1(n4), .B2(
        \REGISTERS[27][1] ), .ZN(n218) );
  NAND4_X1 U302 ( .A1(n221), .A2(n220), .A3(n219), .A4(n218), .ZN(n227) );
  AOI22_X1 U303 ( .A1(n840), .A2(\REGISTERS[0][1] ), .B1(n23), .B2(
        \REGISTERS[16][1] ), .ZN(n225) );
  AOI22_X1 U304 ( .A1(n32), .A2(\REGISTERS[13][1] ), .B1(n6), .B2(
        \REGISTERS[24][1] ), .ZN(n224) );
  AOI22_X1 U305 ( .A1(n28), .A2(\REGISTERS[30][1] ), .B1(n10), .B2(
        \REGISTERS[17][1] ), .ZN(n223) );
  AOI22_X1 U306 ( .A1(n14), .A2(\REGISTERS[29][1] ), .B1(n25), .B2(
        \REGISTERS[15][1] ), .ZN(n222) );
  NAND4_X1 U307 ( .A1(n225), .A2(n224), .A3(n223), .A4(n222), .ZN(n226) );
  NOR4_X1 U308 ( .A1(n229), .A2(n228), .A3(n227), .A4(n226), .ZN(n230) );
  AOI22_X1 U309 ( .A1(n34), .A2(n1778), .B1(n230), .B2(n35), .ZN(N248) );
  AOI22_X1 U310 ( .A1(n7), .A2(\REGISTERS[19][2] ), .B1(n13), .B2(
        \REGISTERS[12][2] ), .ZN(n234) );
  AOI22_X1 U311 ( .A1(n10), .A2(\REGISTERS[17][2] ), .B1(n852), .B2(
        \REGISTERS[9][2] ), .ZN(n233) );
  AOI22_X1 U312 ( .A1(n12), .A2(\REGISTERS[28][2] ), .B1(n15), .B2(
        \REGISTERS[22][2] ), .ZN(n232) );
  AOI22_X1 U313 ( .A1(n16), .A2(\REGISTERS[6][2] ), .B1(n23), .B2(
        \REGISTERS[16][2] ), .ZN(n231) );
  NAND4_X1 U314 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(n250) );
  AOI22_X1 U315 ( .A1(n30), .A2(\REGISTERS[25][2] ), .B1(n24), .B2(
        \REGISTERS[5][2] ), .ZN(n238) );
  AOI22_X1 U316 ( .A1(n22), .A2(\REGISTERS[21][2] ), .B1(n21), .B2(
        \REGISTERS[18][2] ), .ZN(n237) );
  AOI22_X1 U317 ( .A1(n847), .A2(\REGISTERS[1][2] ), .B1(n17), .B2(
        \REGISTERS[20][2] ), .ZN(n236) );
  AOI22_X1 U318 ( .A1(n20), .A2(\REGISTERS[8][2] ), .B1(n18), .B2(
        \REGISTERS[14][2] ), .ZN(n235) );
  NAND4_X1 U319 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(n249) );
  AOI22_X1 U320 ( .A1(n27), .A2(\REGISTERS[26][2] ), .B1(n6), .B2(
        \REGISTERS[24][2] ), .ZN(n242) );
  AOI22_X1 U321 ( .A1(n877), .A2(\REGISTERS[7][2] ), .B1(n19), .B2(
        \REGISTERS[4][2] ), .ZN(n241) );
  AOI22_X1 U322 ( .A1(n1), .A2(\REGISTERS[0][2] ), .B1(n4), .B2(
        \REGISTERS[27][2] ), .ZN(n240) );
  AOI22_X1 U323 ( .A1(n842), .A2(\REGISTERS[2][2] ), .B1(n29), .B2(
        \REGISTERS[11][2] ), .ZN(n239) );
  NAND4_X1 U324 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(n248) );
  AOI22_X1 U325 ( .A1(n31), .A2(\REGISTERS[10][2] ), .B1(n2), .B2(
        \REGISTERS[23][2] ), .ZN(n246) );
  AOI22_X1 U326 ( .A1(n28), .A2(\REGISTERS[30][2] ), .B1(n844), .B2(
        \REGISTERS[31][2] ), .ZN(n245) );
  AOI22_X1 U327 ( .A1(n876), .A2(\REGISTERS[15][2] ), .B1(n854), .B2(
        \REGISTERS[3][2] ), .ZN(n244) );
  AOI22_X1 U328 ( .A1(n32), .A2(\REGISTERS[13][2] ), .B1(n14), .B2(
        \REGISTERS[29][2] ), .ZN(n243) );
  NAND4_X1 U329 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(n247) );
  NOR4_X1 U330 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(n251) );
  AOI22_X1 U331 ( .A1(n34), .A2(n132), .B1(n251), .B2(n36), .ZN(N249) );
  AOI22_X1 U332 ( .A1(n840), .A2(\REGISTERS[0][3] ), .B1(n9), .B2(
        \REGISTERS[9][3] ), .ZN(n255) );
  AOI22_X1 U333 ( .A1(n28), .A2(\REGISTERS[30][3] ), .B1(n22), .B2(
        \REGISTERS[21][3] ), .ZN(n254) );
  AOI22_X1 U334 ( .A1(n16), .A2(\REGISTERS[6][3] ), .B1(n29), .B2(
        \REGISTERS[11][3] ), .ZN(n253) );
  AOI22_X1 U335 ( .A1(n19), .A2(\REGISTERS[4][3] ), .B1(n23), .B2(
        \REGISTERS[16][3] ), .ZN(n252) );
  NAND4_X1 U336 ( .A1(n255), .A2(n254), .A3(n253), .A4(n252), .ZN(n271) );
  AOI22_X1 U337 ( .A1(n21), .A2(\REGISTERS[18][3] ), .B1(n11), .B2(
        \REGISTERS[3][3] ), .ZN(n259) );
  AOI22_X1 U338 ( .A1(n26), .A2(\REGISTERS[7][3] ), .B1(n4), .B2(
        \REGISTERS[27][3] ), .ZN(n258) );
  AOI22_X1 U339 ( .A1(n853), .A2(\REGISTERS[17][3] ), .B1(n5), .B2(
        \REGISTERS[31][3] ), .ZN(n257) );
  AOI22_X1 U340 ( .A1(n30), .A2(\REGISTERS[25][3] ), .B1(n12), .B2(
        \REGISTERS[28][3] ), .ZN(n256) );
  NAND4_X1 U341 ( .A1(n259), .A2(n258), .A3(n257), .A4(n256), .ZN(n270) );
  AOI22_X1 U342 ( .A1(n867), .A2(\REGISTERS[8][3] ), .B1(n25), .B2(
        \REGISTERS[15][3] ), .ZN(n263) );
  AOI22_X1 U343 ( .A1(n871), .A2(\REGISTERS[5][3] ), .B1(n3), .B2(
        \REGISTERS[2][3] ), .ZN(n262) );
  AOI22_X1 U344 ( .A1(n882), .A2(\REGISTERS[10][3] ), .B1(n17), .B2(
        \REGISTERS[20][3] ), .ZN(n261) );
  AOI22_X1 U345 ( .A1(n865), .A2(\REGISTERS[14][3] ), .B1(n8), .B2(
        \REGISTERS[1][3] ), .ZN(n260) );
  NAND4_X1 U346 ( .A1(n263), .A2(n262), .A3(n261), .A4(n260), .ZN(n269) );
  AOI22_X1 U347 ( .A1(n14), .A2(\REGISTERS[29][3] ), .B1(n13), .B2(
        \REGISTERS[12][3] ), .ZN(n267) );
  AOI22_X1 U348 ( .A1(n883), .A2(\REGISTERS[13][3] ), .B1(n15), .B2(
        \REGISTERS[22][3] ), .ZN(n266) );
  AOI22_X1 U349 ( .A1(n841), .A2(\REGISTERS[23][3] ), .B1(n6), .B2(
        \REGISTERS[24][3] ), .ZN(n265) );
  AOI22_X1 U350 ( .A1(n27), .A2(\REGISTERS[26][3] ), .B1(n7), .B2(
        \REGISTERS[19][3] ), .ZN(n264) );
  NAND4_X1 U351 ( .A1(n267), .A2(n266), .A3(n265), .A4(n264), .ZN(n268) );
  NOR4_X1 U352 ( .A1(n271), .A2(n270), .A3(n269), .A4(n268), .ZN(n272) );
  AOI22_X1 U353 ( .A1(n34), .A2(n130), .B1(n272), .B2(n35), .ZN(N250) );
  AOI22_X1 U354 ( .A1(n27), .A2(\REGISTERS[26][4] ), .B1(n19), .B2(
        \REGISTERS[4][4] ), .ZN(n276) );
  AOI22_X1 U355 ( .A1(n868), .A2(\REGISTERS[18][4] ), .B1(n11), .B2(
        \REGISTERS[3][4] ), .ZN(n275) );
  AOI22_X1 U356 ( .A1(n855), .A2(\REGISTERS[28][4] ), .B1(n22), .B2(
        \REGISTERS[21][4] ), .ZN(n274) );
  AOI22_X1 U357 ( .A1(n18), .A2(\REGISTERS[14][4] ), .B1(n852), .B2(
        \REGISTERS[9][4] ), .ZN(n273) );
  NAND4_X1 U358 ( .A1(n276), .A2(n275), .A3(n274), .A4(n273), .ZN(n292) );
  AOI22_X1 U359 ( .A1(n25), .A2(\REGISTERS[15][4] ), .B1(n29), .B2(
        \REGISTERS[11][4] ), .ZN(n280) );
  AOI22_X1 U360 ( .A1(n877), .A2(\REGISTERS[7][4] ), .B1(n1), .B2(
        \REGISTERS[0][4] ), .ZN(n279) );
  AOI22_X1 U361 ( .A1(n864), .A2(\REGISTERS[20][4] ), .B1(n13), .B2(
        \REGISTERS[12][4] ), .ZN(n278) );
  AOI22_X1 U362 ( .A1(n14), .A2(\REGISTERS[29][4] ), .B1(n23), .B2(
        \REGISTERS[16][4] ), .ZN(n277) );
  NAND4_X1 U363 ( .A1(n280), .A2(n279), .A3(n278), .A4(n277), .ZN(n291) );
  AOI22_X1 U364 ( .A1(n2), .A2(\REGISTERS[23][4] ), .B1(n24), .B2(
        \REGISTERS[5][4] ), .ZN(n284) );
  AOI22_X1 U365 ( .A1(n4), .A2(\REGISTERS[27][4] ), .B1(n6), .B2(
        \REGISTERS[24][4] ), .ZN(n283) );
  AOI22_X1 U366 ( .A1(n10), .A2(\REGISTERS[17][4] ), .B1(n7), .B2(
        \REGISTERS[19][4] ), .ZN(n282) );
  AOI22_X1 U367 ( .A1(n32), .A2(\REGISTERS[13][4] ), .B1(n30), .B2(
        \REGISTERS[25][4] ), .ZN(n281) );
  NAND4_X1 U368 ( .A1(n284), .A2(n283), .A3(n282), .A4(n281), .ZN(n290) );
  AOI22_X1 U369 ( .A1(n28), .A2(\REGISTERS[30][4] ), .B1(n15), .B2(
        \REGISTERS[22][4] ), .ZN(n288) );
  AOI22_X1 U370 ( .A1(n20), .A2(\REGISTERS[8][4] ), .B1(n8), .B2(
        \REGISTERS[1][4] ), .ZN(n287) );
  AOI22_X1 U371 ( .A1(n31), .A2(\REGISTERS[10][4] ), .B1(n844), .B2(
        \REGISTERS[31][4] ), .ZN(n286) );
  AOI22_X1 U372 ( .A1(n859), .A2(\REGISTERS[6][4] ), .B1(n3), .B2(
        \REGISTERS[2][4] ), .ZN(n285) );
  NAND4_X1 U373 ( .A1(n288), .A2(n287), .A3(n286), .A4(n285), .ZN(n289) );
  NOR4_X1 U374 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .ZN(n293) );
  AOI22_X1 U375 ( .A1(n34), .A2(n128), .B1(n293), .B2(n36), .ZN(N251) );
  AOI22_X1 U376 ( .A1(n14), .A2(\REGISTERS[29][5] ), .B1(n11), .B2(
        \REGISTERS[3][5] ), .ZN(n297) );
  AOI22_X1 U377 ( .A1(n1), .A2(\REGISTERS[0][5] ), .B1(n17), .B2(
        \REGISTERS[20][5] ), .ZN(n296) );
  AOI22_X1 U378 ( .A1(n845), .A2(\REGISTERS[24][5] ), .B1(n9), .B2(
        \REGISTERS[9][5] ), .ZN(n295) );
  AOI22_X1 U379 ( .A1(n878), .A2(\REGISTERS[26][5] ), .B1(n2), .B2(
        \REGISTERS[23][5] ), .ZN(n294) );
  NAND4_X1 U380 ( .A1(n297), .A2(n296), .A3(n295), .A4(n294), .ZN(n313) );
  AOI22_X1 U381 ( .A1(n30), .A2(\REGISTERS[25][5] ), .B1(n12), .B2(
        \REGISTERS[28][5] ), .ZN(n301) );
  AOI22_X1 U382 ( .A1(n28), .A2(\REGISTERS[30][5] ), .B1(n10), .B2(
        \REGISTERS[17][5] ), .ZN(n300) );
  AOI22_X1 U383 ( .A1(n880), .A2(\REGISTERS[11][5] ), .B1(n23), .B2(
        \REGISTERS[16][5] ), .ZN(n299) );
  AOI22_X1 U384 ( .A1(n22), .A2(\REGISTERS[21][5] ), .B1(n31), .B2(
        \REGISTERS[10][5] ), .ZN(n298) );
  NAND4_X1 U385 ( .A1(n301), .A2(n300), .A3(n299), .A4(n298), .ZN(n312) );
  AOI22_X1 U386 ( .A1(n843), .A2(\REGISTERS[27][5] ), .B1(n24), .B2(
        \REGISTERS[5][5] ), .ZN(n305) );
  AOI22_X1 U387 ( .A1(n16), .A2(\REGISTERS[6][5] ), .B1(n8), .B2(
        \REGISTERS[1][5] ), .ZN(n304) );
  AOI22_X1 U388 ( .A1(n32), .A2(\REGISTERS[13][5] ), .B1(n25), .B2(
        \REGISTERS[15][5] ), .ZN(n303) );
  AOI22_X1 U389 ( .A1(n26), .A2(\REGISTERS[7][5] ), .B1(n15), .B2(
        \REGISTERS[22][5] ), .ZN(n302) );
  NAND4_X1 U390 ( .A1(n305), .A2(n304), .A3(n303), .A4(n302), .ZN(n311) );
  AOI22_X1 U391 ( .A1(n20), .A2(\REGISTERS[8][5] ), .B1(n5), .B2(
        \REGISTERS[31][5] ), .ZN(n309) );
  AOI22_X1 U392 ( .A1(n865), .A2(\REGISTERS[14][5] ), .B1(n3), .B2(
        \REGISTERS[2][5] ), .ZN(n308) );
  AOI22_X1 U393 ( .A1(n868), .A2(\REGISTERS[18][5] ), .B1(n7), .B2(
        \REGISTERS[19][5] ), .ZN(n307) );
  AOI22_X1 U394 ( .A1(n866), .A2(\REGISTERS[4][5] ), .B1(n13), .B2(
        \REGISTERS[12][5] ), .ZN(n306) );
  NAND4_X1 U395 ( .A1(n309), .A2(n308), .A3(n307), .A4(n306), .ZN(n310) );
  NOR4_X1 U396 ( .A1(n313), .A2(n312), .A3(n311), .A4(n310), .ZN(n314) );
  AOI22_X1 U397 ( .A1(n34), .A2(n126), .B1(n314), .B2(n35), .ZN(N252) );
  AOI22_X1 U398 ( .A1(n840), .A2(\REGISTERS[0][6] ), .B1(n21), .B2(
        \REGISTERS[18][6] ), .ZN(n318) );
  AOI22_X1 U399 ( .A1(n22), .A2(\REGISTERS[21][6] ), .B1(n844), .B2(
        \REGISTERS[31][6] ), .ZN(n317) );
  AOI22_X1 U400 ( .A1(n880), .A2(\REGISTERS[11][6] ), .B1(n23), .B2(
        \REGISTERS[16][6] ), .ZN(n316) );
  AOI22_X1 U401 ( .A1(n30), .A2(\REGISTERS[25][6] ), .B1(n7), .B2(
        \REGISTERS[19][6] ), .ZN(n315) );
  NAND4_X1 U402 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(n334) );
  AOI22_X1 U403 ( .A1(n877), .A2(\REGISTERS[7][6] ), .B1(n25), .B2(
        \REGISTERS[15][6] ), .ZN(n322) );
  AOI22_X1 U404 ( .A1(n853), .A2(\REGISTERS[17][6] ), .B1(n8), .B2(
        \REGISTERS[1][6] ), .ZN(n321) );
  AOI22_X1 U405 ( .A1(n11), .A2(\REGISTERS[3][6] ), .B1(n24), .B2(
        \REGISTERS[5][6] ), .ZN(n320) );
  AOI22_X1 U406 ( .A1(n855), .A2(\REGISTERS[28][6] ), .B1(n16), .B2(
        \REGISTERS[6][6] ), .ZN(n319) );
  NAND4_X1 U407 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(n333) );
  AOI22_X1 U408 ( .A1(n18), .A2(\REGISTERS[14][6] ), .B1(n2), .B2(
        \REGISTERS[23][6] ), .ZN(n326) );
  AOI22_X1 U409 ( .A1(n32), .A2(\REGISTERS[13][6] ), .B1(n4), .B2(
        \REGISTERS[27][6] ), .ZN(n325) );
  AOI22_X1 U410 ( .A1(n28), .A2(\REGISTERS[30][6] ), .B1(n20), .B2(
        \REGISTERS[8][6] ), .ZN(n324) );
  AOI22_X1 U411 ( .A1(n864), .A2(\REGISTERS[20][6] ), .B1(n19), .B2(
        \REGISTERS[4][6] ), .ZN(n323) );
  NAND4_X1 U412 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(n332) );
  AOI22_X1 U413 ( .A1(n27), .A2(\REGISTERS[26][6] ), .B1(n6), .B2(
        \REGISTERS[24][6] ), .ZN(n330) );
  AOI22_X1 U414 ( .A1(n3), .A2(\REGISTERS[2][6] ), .B1(n852), .B2(
        \REGISTERS[9][6] ), .ZN(n329) );
  AOI22_X1 U415 ( .A1(n14), .A2(\REGISTERS[29][6] ), .B1(n13), .B2(
        \REGISTERS[12][6] ), .ZN(n328) );
  AOI22_X1 U416 ( .A1(n882), .A2(\REGISTERS[10][6] ), .B1(n15), .B2(
        \REGISTERS[22][6] ), .ZN(n327) );
  NAND4_X1 U417 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(n331) );
  NOR4_X1 U418 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(n335) );
  AOI22_X1 U419 ( .A1(n893), .A2(n124), .B1(n335), .B2(n35), .ZN(N253) );
  AOI22_X1 U420 ( .A1(n12), .A2(\REGISTERS[28][7] ), .B1(n852), .B2(
        \REGISTERS[9][7] ), .ZN(n339) );
  AOI22_X1 U421 ( .A1(n16), .A2(\REGISTERS[6][7] ), .B1(n2), .B2(
        \REGISTERS[23][7] ), .ZN(n338) );
  AOI22_X1 U422 ( .A1(n14), .A2(\REGISTERS[29][7] ), .B1(n23), .B2(
        \REGISTERS[16][7] ), .ZN(n337) );
  AOI22_X1 U423 ( .A1(n6), .A2(\REGISTERS[24][7] ), .B1(n7), .B2(
        \REGISTERS[19][7] ), .ZN(n336) );
  NAND4_X1 U424 ( .A1(n339), .A2(n338), .A3(n337), .A4(n336), .ZN(n355) );
  AOI22_X1 U425 ( .A1(n868), .A2(\REGISTERS[18][7] ), .B1(n24), .B2(
        \REGISTERS[5][7] ), .ZN(n343) );
  AOI22_X1 U426 ( .A1(n28), .A2(\REGISTERS[30][7] ), .B1(n3), .B2(
        \REGISTERS[2][7] ), .ZN(n342) );
  AOI22_X1 U427 ( .A1(n883), .A2(\REGISTERS[13][7] ), .B1(n17), .B2(
        \REGISTERS[20][7] ), .ZN(n341) );
  AOI22_X1 U428 ( .A1(n10), .A2(\REGISTERS[17][7] ), .B1(n13), .B2(
        \REGISTERS[12][7] ), .ZN(n340) );
  NAND4_X1 U429 ( .A1(n343), .A2(n342), .A3(n341), .A4(n340), .ZN(n354) );
  AOI22_X1 U430 ( .A1(n20), .A2(\REGISTERS[8][7] ), .B1(n4), .B2(
        \REGISTERS[27][7] ), .ZN(n347) );
  AOI22_X1 U431 ( .A1(n881), .A2(\REGISTERS[25][7] ), .B1(n22), .B2(
        \REGISTERS[21][7] ), .ZN(n346) );
  AOI22_X1 U432 ( .A1(n31), .A2(\REGISTERS[10][7] ), .B1(n8), .B2(
        \REGISTERS[1][7] ), .ZN(n345) );
  AOI22_X1 U433 ( .A1(n27), .A2(\REGISTERS[26][7] ), .B1(n1), .B2(
        \REGISTERS[0][7] ), .ZN(n344) );
  NAND4_X1 U434 ( .A1(n347), .A2(n346), .A3(n345), .A4(n344), .ZN(n353) );
  AOI22_X1 U435 ( .A1(n876), .A2(\REGISTERS[15][7] ), .B1(n29), .B2(
        \REGISTERS[11][7] ), .ZN(n351) );
  AOI22_X1 U436 ( .A1(n877), .A2(\REGISTERS[7][7] ), .B1(n15), .B2(
        \REGISTERS[22][7] ), .ZN(n350) );
  AOI22_X1 U437 ( .A1(n19), .A2(\REGISTERS[4][7] ), .B1(n844), .B2(
        \REGISTERS[31][7] ), .ZN(n349) );
  AOI22_X1 U438 ( .A1(n18), .A2(\REGISTERS[14][7] ), .B1(n11), .B2(
        \REGISTERS[3][7] ), .ZN(n348) );
  NAND4_X1 U439 ( .A1(n351), .A2(n350), .A3(n349), .A4(n348), .ZN(n352) );
  NOR4_X1 U440 ( .A1(n355), .A2(n354), .A3(n353), .A4(n352), .ZN(n356) );
  AOI22_X1 U441 ( .A1(n893), .A2(n122), .B1(n356), .B2(n36), .ZN(N254) );
  AOI22_X1 U442 ( .A1(n877), .A2(\REGISTERS[7][8] ), .B1(n18), .B2(
        \REGISTERS[14][8] ), .ZN(n360) );
  AOI22_X1 U443 ( .A1(n879), .A2(\REGISTERS[30][8] ), .B1(n32), .B2(
        \REGISTERS[13][8] ), .ZN(n359) );
  AOI22_X1 U444 ( .A1(n27), .A2(\REGISTERS[26][8] ), .B1(n30), .B2(
        \REGISTERS[25][8] ), .ZN(n358) );
  AOI22_X1 U445 ( .A1(n12), .A2(\REGISTERS[28][8] ), .B1(n1), .B2(
        \REGISTERS[0][8] ), .ZN(n357) );
  NAND4_X1 U446 ( .A1(n360), .A2(n359), .A3(n358), .A4(n357), .ZN(n376) );
  AOI22_X1 U447 ( .A1(n20), .A2(\REGISTERS[8][8] ), .B1(n19), .B2(
        \REGISTERS[4][8] ), .ZN(n364) );
  AOI22_X1 U448 ( .A1(n857), .A2(\REGISTERS[29][8] ), .B1(n7), .B2(
        \REGISTERS[19][8] ), .ZN(n363) );
  AOI22_X1 U449 ( .A1(n8), .A2(\REGISTERS[1][8] ), .B1(n844), .B2(
        \REGISTERS[31][8] ), .ZN(n362) );
  AOI22_X1 U450 ( .A1(n843), .A2(\REGISTERS[27][8] ), .B1(n11), .B2(
        \REGISTERS[3][8] ), .ZN(n361) );
  NAND4_X1 U451 ( .A1(n364), .A2(n363), .A3(n362), .A4(n361), .ZN(n375) );
  AOI22_X1 U452 ( .A1(n869), .A2(\REGISTERS[21][8] ), .B1(n3), .B2(
        \REGISTERS[2][8] ), .ZN(n368) );
  AOI22_X1 U453 ( .A1(n6), .A2(\REGISTERS[24][8] ), .B1(n13), .B2(
        \REGISTERS[12][8] ), .ZN(n367) );
  AOI22_X1 U454 ( .A1(n16), .A2(\REGISTERS[6][8] ), .B1(n23), .B2(
        \REGISTERS[16][8] ), .ZN(n366) );
  AOI22_X1 U455 ( .A1(n10), .A2(\REGISTERS[17][8] ), .B1(n24), .B2(
        \REGISTERS[5][8] ), .ZN(n365) );
  NAND4_X1 U456 ( .A1(n368), .A2(n367), .A3(n366), .A4(n365), .ZN(n374) );
  AOI22_X1 U457 ( .A1(n868), .A2(\REGISTERS[18][8] ), .B1(n852), .B2(
        \REGISTERS[9][8] ), .ZN(n372) );
  AOI22_X1 U458 ( .A1(n25), .A2(\REGISTERS[15][8] ), .B1(n17), .B2(
        \REGISTERS[20][8] ), .ZN(n371) );
  AOI22_X1 U459 ( .A1(n841), .A2(\REGISTERS[23][8] ), .B1(n15), .B2(
        \REGISTERS[22][8] ), .ZN(n370) );
  AOI22_X1 U460 ( .A1(n31), .A2(\REGISTERS[10][8] ), .B1(n29), .B2(
        \REGISTERS[11][8] ), .ZN(n369) );
  NAND4_X1 U461 ( .A1(n372), .A2(n371), .A3(n370), .A4(n369), .ZN(n373) );
  NOR4_X1 U462 ( .A1(n376), .A2(n375), .A3(n374), .A4(n373), .ZN(n377) );
  AOI22_X1 U463 ( .A1(n893), .A2(n120), .B1(n377), .B2(n36), .ZN(N255) );
  AOI22_X1 U464 ( .A1(n20), .A2(\REGISTERS[8][9] ), .B1(n18), .B2(
        \REGISTERS[14][9] ), .ZN(n381) );
  AOI22_X1 U465 ( .A1(n864), .A2(\REGISTERS[20][9] ), .B1(n15), .B2(
        \REGISTERS[22][9] ), .ZN(n380) );
  AOI22_X1 U466 ( .A1(n22), .A2(\REGISTERS[21][9] ), .B1(n21), .B2(
        \REGISTERS[18][9] ), .ZN(n379) );
  AOI22_X1 U467 ( .A1(n31), .A2(\REGISTERS[10][9] ), .B1(n25), .B2(
        \REGISTERS[15][9] ), .ZN(n378) );
  NAND4_X1 U468 ( .A1(n381), .A2(n380), .A3(n379), .A4(n378), .ZN(n397) );
  AOI22_X1 U469 ( .A1(n857), .A2(\REGISTERS[29][9] ), .B1(n16), .B2(
        \REGISTERS[6][9] ), .ZN(n385) );
  AOI22_X1 U470 ( .A1(n871), .A2(\REGISTERS[5][9] ), .B1(n844), .B2(
        \REGISTERS[31][9] ), .ZN(n384) );
  AOI22_X1 U471 ( .A1(n854), .A2(\REGISTERS[3][9] ), .B1(n852), .B2(
        \REGISTERS[9][9] ), .ZN(n383) );
  AOI22_X1 U472 ( .A1(n840), .A2(\REGISTERS[0][9] ), .B1(n7), .B2(
        \REGISTERS[19][9] ), .ZN(n382) );
  NAND4_X1 U473 ( .A1(n385), .A2(n384), .A3(n383), .A4(n382), .ZN(n396) );
  AOI22_X1 U474 ( .A1(n879), .A2(\REGISTERS[30][9] ), .B1(n3), .B2(
        \REGISTERS[2][9] ), .ZN(n389) );
  AOI22_X1 U475 ( .A1(n843), .A2(\REGISTERS[27][9] ), .B1(n29), .B2(
        \REGISTERS[11][9] ), .ZN(n388) );
  AOI22_X1 U476 ( .A1(n878), .A2(\REGISTERS[26][9] ), .B1(n19), .B2(
        \REGISTERS[4][9] ), .ZN(n387) );
  AOI22_X1 U477 ( .A1(n847), .A2(\REGISTERS[1][9] ), .B1(n6), .B2(
        \REGISTERS[24][9] ), .ZN(n386) );
  NAND4_X1 U478 ( .A1(n389), .A2(n388), .A3(n387), .A4(n386), .ZN(n395) );
  AOI22_X1 U479 ( .A1(n10), .A2(\REGISTERS[17][9] ), .B1(n13), .B2(
        \REGISTERS[12][9] ), .ZN(n393) );
  AOI22_X1 U480 ( .A1(n12), .A2(\REGISTERS[28][9] ), .B1(n2), .B2(
        \REGISTERS[23][9] ), .ZN(n392) );
  AOI22_X1 U481 ( .A1(n877), .A2(\REGISTERS[7][9] ), .B1(n23), .B2(
        \REGISTERS[16][9] ), .ZN(n391) );
  AOI22_X1 U482 ( .A1(n32), .A2(\REGISTERS[13][9] ), .B1(n30), .B2(
        \REGISTERS[25][9] ), .ZN(n390) );
  NAND4_X1 U483 ( .A1(n393), .A2(n392), .A3(n391), .A4(n390), .ZN(n394) );
  NOR4_X1 U484 ( .A1(n397), .A2(n396), .A3(n395), .A4(n394), .ZN(n398) );
  AOI22_X1 U485 ( .A1(n893), .A2(n118), .B1(n398), .B2(n35), .ZN(N256) );
  AOI22_X1 U486 ( .A1(n847), .A2(\REGISTERS[1][10] ), .B1(n858), .B2(
        \REGISTERS[22][10] ), .ZN(n402) );
  AOI22_X1 U487 ( .A1(n845), .A2(\REGISTERS[24][10] ), .B1(n844), .B2(
        \REGISTERS[31][10] ), .ZN(n401) );
  AOI22_X1 U488 ( .A1(n18), .A2(\REGISTERS[14][10] ), .B1(n856), .B2(
        \REGISTERS[12][10] ), .ZN(n400) );
  AOI22_X1 U489 ( .A1(n22), .A2(\REGISTERS[21][10] ), .B1(n870), .B2(
        \REGISTERS[16][10] ), .ZN(n399) );
  NAND4_X1 U490 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(n418) );
  AOI22_X1 U491 ( .A1(n31), .A2(\REGISTERS[10][10] ), .B1(n24), .B2(
        \REGISTERS[5][10] ), .ZN(n406) );
  AOI22_X1 U492 ( .A1(n25), .A2(\REGISTERS[15][10] ), .B1(n2), .B2(
        \REGISTERS[23][10] ), .ZN(n405) );
  AOI22_X1 U493 ( .A1(n843), .A2(\REGISTERS[27][10] ), .B1(n17), .B2(
        \REGISTERS[20][10] ), .ZN(n404) );
  AOI22_X1 U494 ( .A1(n881), .A2(\REGISTERS[25][10] ), .B1(n3), .B2(
        \REGISTERS[2][10] ), .ZN(n403) );
  NAND4_X1 U495 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(n417) );
  AOI22_X1 U496 ( .A1(n10), .A2(\REGISTERS[17][10] ), .B1(n16), .B2(
        \REGISTERS[6][10] ), .ZN(n410) );
  AOI22_X1 U497 ( .A1(n28), .A2(\REGISTERS[30][10] ), .B1(n19), .B2(
        \REGISTERS[4][10] ), .ZN(n409) );
  AOI22_X1 U498 ( .A1(n12), .A2(\REGISTERS[28][10] ), .B1(n29), .B2(
        \REGISTERS[11][10] ), .ZN(n408) );
  AOI22_X1 U499 ( .A1(n877), .A2(\REGISTERS[7][10] ), .B1(n11), .B2(
        \REGISTERS[3][10] ), .ZN(n407) );
  NAND4_X1 U500 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(n416) );
  AOI22_X1 U501 ( .A1(n32), .A2(\REGISTERS[13][10] ), .B1(n7), .B2(
        \REGISTERS[19][10] ), .ZN(n414) );
  AOI22_X1 U502 ( .A1(n840), .A2(\REGISTERS[0][10] ), .B1(n852), .B2(
        \REGISTERS[9][10] ), .ZN(n413) );
  AOI22_X1 U503 ( .A1(n27), .A2(\REGISTERS[26][10] ), .B1(n14), .B2(
        \REGISTERS[29][10] ), .ZN(n412) );
  AOI22_X1 U504 ( .A1(n20), .A2(\REGISTERS[8][10] ), .B1(n21), .B2(
        \REGISTERS[18][10] ), .ZN(n411) );
  NAND4_X1 U505 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(n415) );
  NOR4_X1 U506 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(n419) );
  AOI22_X1 U507 ( .A1(n893), .A2(n116), .B1(n419), .B2(n36), .ZN(N257) );
  AOI22_X1 U508 ( .A1(n10), .A2(\REGISTERS[17][11] ), .B1(n13), .B2(
        \REGISTERS[12][11] ), .ZN(n423) );
  AOI22_X1 U509 ( .A1(n14), .A2(\REGISTERS[29][11] ), .B1(n852), .B2(
        \REGISTERS[9][11] ), .ZN(n422) );
  AOI22_X1 U510 ( .A1(n31), .A2(\REGISTERS[10][11] ), .B1(n2), .B2(
        \REGISTERS[23][11] ), .ZN(n421) );
  AOI22_X1 U511 ( .A1(n22), .A2(\REGISTERS[21][11] ), .B1(n21), .B2(
        \REGISTERS[18][11] ), .ZN(n420) );
  NAND4_X1 U512 ( .A1(n423), .A2(n422), .A3(n421), .A4(n420), .ZN(n439) );
  AOI22_X1 U513 ( .A1(n19), .A2(\REGISTERS[4][11] ), .B1(n870), .B2(
        \REGISTERS[16][11] ), .ZN(n427) );
  AOI22_X1 U514 ( .A1(n12), .A2(\REGISTERS[28][11] ), .B1(n846), .B2(
        \REGISTERS[19][11] ), .ZN(n426) );
  AOI22_X1 U515 ( .A1(n27), .A2(\REGISTERS[26][11] ), .B1(n11), .B2(
        \REGISTERS[3][11] ), .ZN(n425) );
  AOI22_X1 U516 ( .A1(n30), .A2(\REGISTERS[25][11] ), .B1(n8), .B2(
        \REGISTERS[1][11] ), .ZN(n424) );
  NAND4_X1 U517 ( .A1(n427), .A2(n426), .A3(n425), .A4(n424), .ZN(n438) );
  AOI22_X1 U518 ( .A1(n877), .A2(\REGISTERS[7][11] ), .B1(n32), .B2(
        \REGISTERS[13][11] ), .ZN(n431) );
  AOI22_X1 U519 ( .A1(n28), .A2(\REGISTERS[30][11] ), .B1(n16), .B2(
        \REGISTERS[6][11] ), .ZN(n430) );
  AOI22_X1 U520 ( .A1(n20), .A2(\REGISTERS[8][11] ), .B1(n844), .B2(
        \REGISTERS[31][11] ), .ZN(n429) );
  AOI22_X1 U521 ( .A1(n843), .A2(\REGISTERS[27][11] ), .B1(n17), .B2(
        \REGISTERS[20][11] ), .ZN(n428) );
  NAND4_X1 U522 ( .A1(n431), .A2(n430), .A3(n429), .A4(n428), .ZN(n437) );
  AOI22_X1 U523 ( .A1(n840), .A2(\REGISTERS[0][11] ), .B1(n3), .B2(
        \REGISTERS[2][11] ), .ZN(n435) );
  AOI22_X1 U524 ( .A1(n25), .A2(\REGISTERS[15][11] ), .B1(n29), .B2(
        \REGISTERS[11][11] ), .ZN(n434) );
  AOI22_X1 U525 ( .A1(n871), .A2(\REGISTERS[5][11] ), .B1(n858), .B2(
        \REGISTERS[22][11] ), .ZN(n433) );
  AOI22_X1 U526 ( .A1(n865), .A2(\REGISTERS[14][11] ), .B1(n6), .B2(
        \REGISTERS[24][11] ), .ZN(n432) );
  NAND4_X1 U527 ( .A1(n435), .A2(n434), .A3(n433), .A4(n432), .ZN(n436) );
  NOR4_X1 U528 ( .A1(n439), .A2(n438), .A3(n437), .A4(n436), .ZN(n440) );
  AOI22_X1 U529 ( .A1(n893), .A2(n114), .B1(n440), .B2(n35), .ZN(N258) );
  AOI22_X1 U530 ( .A1(n22), .A2(\REGISTERS[21][12] ), .B1(n17), .B2(
        \REGISTERS[20][12] ), .ZN(n444) );
  AOI22_X1 U531 ( .A1(n27), .A2(\REGISTERS[26][12] ), .B1(n5), .B2(
        \REGISTERS[31][12] ), .ZN(n443) );
  AOI22_X1 U532 ( .A1(n28), .A2(\REGISTERS[30][12] ), .B1(n11), .B2(
        \REGISTERS[3][12] ), .ZN(n442) );
  AOI22_X1 U533 ( .A1(n30), .A2(\REGISTERS[25][12] ), .B1(n1), .B2(
        \REGISTERS[0][12] ), .ZN(n441) );
  NAND4_X1 U534 ( .A1(n444), .A2(n443), .A3(n442), .A4(n441), .ZN(n460) );
  AOI22_X1 U535 ( .A1(n16), .A2(\REGISTERS[6][12] ), .B1(n3), .B2(
        \REGISTERS[2][12] ), .ZN(n448) );
  AOI22_X1 U536 ( .A1(n843), .A2(\REGISTERS[27][12] ), .B1(n880), .B2(
        \REGISTERS[11][12] ), .ZN(n447) );
  AOI22_X1 U537 ( .A1(n10), .A2(\REGISTERS[17][12] ), .B1(n18), .B2(
        \REGISTERS[14][12] ), .ZN(n446) );
  AOI22_X1 U538 ( .A1(n847), .A2(\REGISTERS[1][12] ), .B1(n9), .B2(
        \REGISTERS[9][12] ), .ZN(n445) );
  NAND4_X1 U539 ( .A1(n448), .A2(n447), .A3(n446), .A4(n445), .ZN(n459) );
  AOI22_X1 U540 ( .A1(n25), .A2(\REGISTERS[15][12] ), .B1(n846), .B2(
        \REGISTERS[19][12] ), .ZN(n452) );
  AOI22_X1 U541 ( .A1(n866), .A2(\REGISTERS[4][12] ), .B1(n23), .B2(
        \REGISTERS[16][12] ), .ZN(n451) );
  AOI22_X1 U542 ( .A1(n32), .A2(\REGISTERS[13][12] ), .B1(n6), .B2(
        \REGISTERS[24][12] ), .ZN(n450) );
  AOI22_X1 U543 ( .A1(n20), .A2(\REGISTERS[8][12] ), .B1(n2), .B2(
        \REGISTERS[23][12] ), .ZN(n449) );
  NAND4_X1 U544 ( .A1(n452), .A2(n451), .A3(n450), .A4(n449), .ZN(n458) );
  AOI22_X1 U545 ( .A1(n14), .A2(\REGISTERS[29][12] ), .B1(n21), .B2(
        \REGISTERS[18][12] ), .ZN(n456) );
  AOI22_X1 U546 ( .A1(n12), .A2(\REGISTERS[28][12] ), .B1(n31), .B2(
        \REGISTERS[10][12] ), .ZN(n455) );
  AOI22_X1 U547 ( .A1(n26), .A2(\REGISTERS[7][12] ), .B1(n15), .B2(
        \REGISTERS[22][12] ), .ZN(n454) );
  AOI22_X1 U548 ( .A1(n856), .A2(\REGISTERS[12][12] ), .B1(n24), .B2(
        \REGISTERS[5][12] ), .ZN(n453) );
  NAND4_X1 U549 ( .A1(n456), .A2(n455), .A3(n454), .A4(n453), .ZN(n457) );
  NOR4_X1 U550 ( .A1(n460), .A2(n459), .A3(n458), .A4(n457), .ZN(n461) );
  AOI22_X1 U551 ( .A1(n33), .A2(n112), .B1(n461), .B2(n36), .ZN(N259) );
  AOI22_X1 U552 ( .A1(n845), .A2(\REGISTERS[24][13] ), .B1(n856), .B2(
        \REGISTERS[12][13] ), .ZN(n465) );
  AOI22_X1 U553 ( .A1(n10), .A2(\REGISTERS[17][13] ), .B1(n31), .B2(
        \REGISTERS[10][13] ), .ZN(n464) );
  AOI22_X1 U554 ( .A1(n30), .A2(\REGISTERS[25][13] ), .B1(n23), .B2(
        \REGISTERS[16][13] ), .ZN(n463) );
  AOI22_X1 U555 ( .A1(n12), .A2(\REGISTERS[28][13] ), .B1(n1), .B2(
        \REGISTERS[0][13] ), .ZN(n462) );
  NAND4_X1 U556 ( .A1(n465), .A2(n464), .A3(n463), .A4(n462), .ZN(n481) );
  AOI22_X1 U557 ( .A1(n842), .A2(\REGISTERS[2][13] ), .B1(n5), .B2(
        \REGISTERS[31][13] ), .ZN(n469) );
  AOI22_X1 U558 ( .A1(n2), .A2(\REGISTERS[23][13] ), .B1(n15), .B2(
        \REGISTERS[22][13] ), .ZN(n468) );
  AOI22_X1 U559 ( .A1(n32), .A2(\REGISTERS[13][13] ), .B1(n880), .B2(
        \REGISTERS[11][13] ), .ZN(n467) );
  AOI22_X1 U560 ( .A1(n846), .A2(\REGISTERS[19][13] ), .B1(n9), .B2(
        \REGISTERS[9][13] ), .ZN(n466) );
  NAND4_X1 U561 ( .A1(n469), .A2(n468), .A3(n467), .A4(n466), .ZN(n480) );
  AOI22_X1 U562 ( .A1(n876), .A2(\REGISTERS[15][13] ), .B1(n4), .B2(
        \REGISTERS[27][13] ), .ZN(n473) );
  AOI22_X1 U563 ( .A1(n867), .A2(\REGISTERS[8][13] ), .B1(n871), .B2(
        \REGISTERS[5][13] ), .ZN(n472) );
  AOI22_X1 U564 ( .A1(n14), .A2(\REGISTERS[29][13] ), .B1(n864), .B2(
        \REGISTERS[20][13] ), .ZN(n471) );
  AOI22_X1 U565 ( .A1(n859), .A2(\REGISTERS[6][13] ), .B1(n18), .B2(
        \REGISTERS[14][13] ), .ZN(n470) );
  NAND4_X1 U566 ( .A1(n473), .A2(n472), .A3(n471), .A4(n470), .ZN(n479) );
  AOI22_X1 U567 ( .A1(n847), .A2(\REGISTERS[1][13] ), .B1(n854), .B2(
        \REGISTERS[3][13] ), .ZN(n477) );
  AOI22_X1 U568 ( .A1(n26), .A2(\REGISTERS[7][13] ), .B1(n19), .B2(
        \REGISTERS[4][13] ), .ZN(n476) );
  AOI22_X1 U569 ( .A1(n27), .A2(\REGISTERS[26][13] ), .B1(n21), .B2(
        \REGISTERS[18][13] ), .ZN(n475) );
  AOI22_X1 U570 ( .A1(n28), .A2(\REGISTERS[30][13] ), .B1(n22), .B2(
        \REGISTERS[21][13] ), .ZN(n474) );
  NAND4_X1 U571 ( .A1(n477), .A2(n476), .A3(n475), .A4(n474), .ZN(n478) );
  NOR4_X1 U572 ( .A1(n481), .A2(n480), .A3(n479), .A4(n478), .ZN(n482) );
  AOI22_X1 U573 ( .A1(n33), .A2(n110), .B1(n482), .B2(n35), .ZN(N260) );
  AOI22_X1 U574 ( .A1(n10), .A2(\REGISTERS[17][14] ), .B1(n23), .B2(
        \REGISTERS[16][14] ), .ZN(n486) );
  AOI22_X1 U575 ( .A1(n30), .A2(\REGISTERS[25][14] ), .B1(n864), .B2(
        \REGISTERS[20][14] ), .ZN(n485) );
  AOI22_X1 U576 ( .A1(n14), .A2(\REGISTERS[29][14] ), .B1(n1), .B2(
        \REGISTERS[0][14] ), .ZN(n484) );
  AOI22_X1 U577 ( .A1(n7), .A2(\REGISTERS[19][14] ), .B1(n13), .B2(
        \REGISTERS[12][14] ), .ZN(n483) );
  NAND4_X1 U578 ( .A1(n486), .A2(n485), .A3(n484), .A4(n483), .ZN(n502) );
  AOI22_X1 U579 ( .A1(n866), .A2(\REGISTERS[4][14] ), .B1(n15), .B2(
        \REGISTERS[22][14] ), .ZN(n490) );
  AOI22_X1 U580 ( .A1(n27), .A2(\REGISTERS[26][14] ), .B1(n25), .B2(
        \REGISTERS[15][14] ), .ZN(n489) );
  AOI22_X1 U581 ( .A1(n859), .A2(\REGISTERS[6][14] ), .B1(n6), .B2(
        \REGISTERS[24][14] ), .ZN(n488) );
  AOI22_X1 U582 ( .A1(n880), .A2(\REGISTERS[11][14] ), .B1(n9), .B2(
        \REGISTERS[9][14] ), .ZN(n487) );
  NAND4_X1 U583 ( .A1(n490), .A2(n489), .A3(n488), .A4(n487), .ZN(n501) );
  AOI22_X1 U584 ( .A1(n12), .A2(\REGISTERS[28][14] ), .B1(n8), .B2(
        \REGISTERS[1][14] ), .ZN(n494) );
  AOI22_X1 U585 ( .A1(n842), .A2(\REGISTERS[2][14] ), .B1(n5), .B2(
        \REGISTERS[31][14] ), .ZN(n493) );
  AOI22_X1 U586 ( .A1(n26), .A2(\REGISTERS[7][14] ), .B1(n2), .B2(
        \REGISTERS[23][14] ), .ZN(n492) );
  AOI22_X1 U587 ( .A1(n28), .A2(\REGISTERS[30][14] ), .B1(n4), .B2(
        \REGISTERS[27][14] ), .ZN(n491) );
  NAND4_X1 U588 ( .A1(n494), .A2(n493), .A3(n492), .A4(n491), .ZN(n500) );
  AOI22_X1 U589 ( .A1(n31), .A2(\REGISTERS[10][14] ), .B1(n20), .B2(
        \REGISTERS[8][14] ), .ZN(n498) );
  AOI22_X1 U590 ( .A1(n868), .A2(\REGISTERS[18][14] ), .B1(n871), .B2(
        \REGISTERS[5][14] ), .ZN(n497) );
  AOI22_X1 U591 ( .A1(n869), .A2(\REGISTERS[21][14] ), .B1(n18), .B2(
        \REGISTERS[14][14] ), .ZN(n496) );
  AOI22_X1 U592 ( .A1(n32), .A2(\REGISTERS[13][14] ), .B1(n854), .B2(
        \REGISTERS[3][14] ), .ZN(n495) );
  NAND4_X1 U593 ( .A1(n498), .A2(n497), .A3(n496), .A4(n495), .ZN(n499) );
  NOR4_X1 U594 ( .A1(n502), .A2(n501), .A3(n500), .A4(n499), .ZN(n503) );
  AOI22_X1 U595 ( .A1(n33), .A2(n108), .B1(n503), .B2(n36), .ZN(N261) );
  AOI22_X1 U596 ( .A1(n4), .A2(\REGISTERS[27][15] ), .B1(n17), .B2(
        \REGISTERS[20][15] ), .ZN(n507) );
  AOI22_X1 U597 ( .A1(n30), .A2(\REGISTERS[25][15] ), .B1(n14), .B2(
        \REGISTERS[29][15] ), .ZN(n506) );
  AOI22_X1 U598 ( .A1(n854), .A2(\REGISTERS[3][15] ), .B1(n13), .B2(
        \REGISTERS[12][15] ), .ZN(n505) );
  AOI22_X1 U599 ( .A1(n32), .A2(\REGISTERS[13][15] ), .B1(n12), .B2(
        \REGISTERS[28][15] ), .ZN(n504) );
  NAND4_X1 U600 ( .A1(n507), .A2(n506), .A3(n505), .A4(n504), .ZN(n523) );
  AOI22_X1 U601 ( .A1(n876), .A2(\REGISTERS[15][15] ), .B1(n21), .B2(
        \REGISTERS[18][15] ), .ZN(n511) );
  AOI22_X1 U602 ( .A1(n846), .A2(\REGISTERS[19][15] ), .B1(n9), .B2(
        \REGISTERS[9][15] ), .ZN(n510) );
  AOI22_X1 U603 ( .A1(n858), .A2(\REGISTERS[22][15] ), .B1(n23), .B2(
        \REGISTERS[16][15] ), .ZN(n509) );
  AOI22_X1 U604 ( .A1(n840), .A2(\REGISTERS[0][15] ), .B1(n8), .B2(
        \REGISTERS[1][15] ), .ZN(n508) );
  NAND4_X1 U605 ( .A1(n511), .A2(n510), .A3(n509), .A4(n508), .ZN(n522) );
  AOI22_X1 U606 ( .A1(n26), .A2(\REGISTERS[7][15] ), .B1(n18), .B2(
        \REGISTERS[14][15] ), .ZN(n515) );
  AOI22_X1 U607 ( .A1(n22), .A2(\REGISTERS[21][15] ), .B1(n16), .B2(
        \REGISTERS[6][15] ), .ZN(n514) );
  AOI22_X1 U608 ( .A1(n845), .A2(\REGISTERS[24][15] ), .B1(n24), .B2(
        \REGISTERS[5][15] ), .ZN(n513) );
  AOI22_X1 U609 ( .A1(n10), .A2(\REGISTERS[17][15] ), .B1(n842), .B2(
        \REGISTERS[2][15] ), .ZN(n512) );
  NAND4_X1 U610 ( .A1(n515), .A2(n514), .A3(n513), .A4(n512), .ZN(n521) );
  AOI22_X1 U611 ( .A1(n867), .A2(\REGISTERS[8][15] ), .B1(n5), .B2(
        \REGISTERS[31][15] ), .ZN(n519) );
  AOI22_X1 U612 ( .A1(n28), .A2(\REGISTERS[30][15] ), .B1(n2), .B2(
        \REGISTERS[23][15] ), .ZN(n518) );
  AOI22_X1 U613 ( .A1(n866), .A2(\REGISTERS[4][15] ), .B1(n29), .B2(
        \REGISTERS[11][15] ), .ZN(n517) );
  AOI22_X1 U614 ( .A1(n27), .A2(\REGISTERS[26][15] ), .B1(n31), .B2(
        \REGISTERS[10][15] ), .ZN(n516) );
  NAND4_X1 U615 ( .A1(n519), .A2(n518), .A3(n517), .A4(n516), .ZN(n520) );
  NOR4_X1 U616 ( .A1(n523), .A2(n522), .A3(n521), .A4(n520), .ZN(n524) );
  AOI22_X1 U617 ( .A1(n33), .A2(n106), .B1(n524), .B2(n35), .ZN(N262) );
  AOI22_X1 U618 ( .A1(n853), .A2(\REGISTERS[17][16] ), .B1(n23), .B2(
        \REGISTERS[16][16] ), .ZN(n528) );
  AOI22_X1 U619 ( .A1(n30), .A2(\REGISTERS[25][16] ), .B1(n13), .B2(
        \REGISTERS[12][16] ), .ZN(n527) );
  AOI22_X1 U620 ( .A1(n26), .A2(\REGISTERS[7][16] ), .B1(n868), .B2(
        \REGISTERS[18][16] ), .ZN(n526) );
  AOI22_X1 U621 ( .A1(n866), .A2(\REGISTERS[4][16] ), .B1(n5), .B2(
        \REGISTERS[31][16] ), .ZN(n525) );
  NAND4_X1 U622 ( .A1(n528), .A2(n527), .A3(n526), .A4(n525), .ZN(n544) );
  AOI22_X1 U623 ( .A1(n859), .A2(\REGISTERS[6][16] ), .B1(n9), .B2(
        \REGISTERS[9][16] ), .ZN(n532) );
  AOI22_X1 U624 ( .A1(n32), .A2(\REGISTERS[13][16] ), .B1(n842), .B2(
        \REGISTERS[2][16] ), .ZN(n531) );
  AOI22_X1 U625 ( .A1(n14), .A2(\REGISTERS[29][16] ), .B1(n4), .B2(
        \REGISTERS[27][16] ), .ZN(n530) );
  AOI22_X1 U626 ( .A1(n865), .A2(\REGISTERS[14][16] ), .B1(n7), .B2(
        \REGISTERS[19][16] ), .ZN(n529) );
  NAND4_X1 U627 ( .A1(n532), .A2(n531), .A3(n530), .A4(n529), .ZN(n543) );
  AOI22_X1 U628 ( .A1(n876), .A2(\REGISTERS[15][16] ), .B1(n17), .B2(
        \REGISTERS[20][16] ), .ZN(n536) );
  AOI22_X1 U629 ( .A1(n2), .A2(\REGISTERS[23][16] ), .B1(n29), .B2(
        \REGISTERS[11][16] ), .ZN(n535) );
  AOI22_X1 U630 ( .A1(n31), .A2(\REGISTERS[10][16] ), .B1(n1), .B2(
        \REGISTERS[0][16] ), .ZN(n534) );
  AOI22_X1 U631 ( .A1(n8), .A2(\REGISTERS[1][16] ), .B1(n15), .B2(
        \REGISTERS[22][16] ), .ZN(n533) );
  NAND4_X1 U632 ( .A1(n536), .A2(n535), .A3(n534), .A4(n533), .ZN(n542) );
  AOI22_X1 U633 ( .A1(n28), .A2(\REGISTERS[30][16] ), .B1(n20), .B2(
        \REGISTERS[8][16] ), .ZN(n540) );
  AOI22_X1 U634 ( .A1(n27), .A2(\REGISTERS[26][16] ), .B1(n24), .B2(
        \REGISTERS[5][16] ), .ZN(n539) );
  AOI22_X1 U635 ( .A1(n12), .A2(\REGISTERS[28][16] ), .B1(n22), .B2(
        \REGISTERS[21][16] ), .ZN(n538) );
  AOI22_X1 U636 ( .A1(n845), .A2(\REGISTERS[24][16] ), .B1(n11), .B2(
        \REGISTERS[3][16] ), .ZN(n537) );
  NAND4_X1 U637 ( .A1(n540), .A2(n539), .A3(n538), .A4(n537), .ZN(n541) );
  NOR4_X1 U638 ( .A1(n544), .A2(n543), .A3(n542), .A4(n541), .ZN(n545) );
  AOI22_X1 U639 ( .A1(n33), .A2(n104), .B1(n545), .B2(n36), .ZN(N263) );
  AOI22_X1 U640 ( .A1(n876), .A2(\REGISTERS[15][17] ), .B1(n24), .B2(
        \REGISTERS[5][17] ), .ZN(n549) );
  AOI22_X1 U641 ( .A1(n32), .A2(\REGISTERS[13][17] ), .B1(n3), .B2(
        \REGISTERS[2][17] ), .ZN(n548) );
  AOI22_X1 U642 ( .A1(n859), .A2(\REGISTERS[6][17] ), .B1(n5), .B2(
        \REGISTERS[31][17] ), .ZN(n547) );
  AOI22_X1 U643 ( .A1(n868), .A2(\REGISTERS[18][17] ), .B1(n6), .B2(
        \REGISTERS[24][17] ), .ZN(n546) );
  NAND4_X1 U644 ( .A1(n549), .A2(n548), .A3(n547), .A4(n546), .ZN(n565) );
  AOI22_X1 U645 ( .A1(n854), .A2(\REGISTERS[3][17] ), .B1(n15), .B2(
        \REGISTERS[22][17] ), .ZN(n553) );
  AOI22_X1 U646 ( .A1(n14), .A2(\REGISTERS[29][17] ), .B1(n18), .B2(
        \REGISTERS[14][17] ), .ZN(n552) );
  AOI22_X1 U647 ( .A1(n1), .A2(\REGISTERS[0][17] ), .B1(n23), .B2(
        \REGISTERS[16][17] ), .ZN(n551) );
  AOI22_X1 U648 ( .A1(n853), .A2(\REGISTERS[17][17] ), .B1(n31), .B2(
        \REGISTERS[10][17] ), .ZN(n550) );
  NAND4_X1 U649 ( .A1(n553), .A2(n552), .A3(n551), .A4(n550), .ZN(n564) );
  AOI22_X1 U650 ( .A1(n869), .A2(\REGISTERS[21][17] ), .B1(n9), .B2(
        \REGISTERS[9][17] ), .ZN(n557) );
  AOI22_X1 U651 ( .A1(n28), .A2(\REGISTERS[30][17] ), .B1(n27), .B2(
        \REGISTERS[26][17] ), .ZN(n556) );
  AOI22_X1 U652 ( .A1(n843), .A2(\REGISTERS[27][17] ), .B1(n19), .B2(
        \REGISTERS[4][17] ), .ZN(n555) );
  AOI22_X1 U653 ( .A1(n30), .A2(\REGISTERS[25][17] ), .B1(n7), .B2(
        \REGISTERS[19][17] ), .ZN(n554) );
  NAND4_X1 U654 ( .A1(n557), .A2(n556), .A3(n555), .A4(n554), .ZN(n563) );
  AOI22_X1 U655 ( .A1(n855), .A2(\REGISTERS[28][17] ), .B1(n29), .B2(
        \REGISTERS[11][17] ), .ZN(n561) );
  AOI22_X1 U656 ( .A1(n26), .A2(\REGISTERS[7][17] ), .B1(n17), .B2(
        \REGISTERS[20][17] ), .ZN(n560) );
  AOI22_X1 U657 ( .A1(n867), .A2(\REGISTERS[8][17] ), .B1(n2), .B2(
        \REGISTERS[23][17] ), .ZN(n559) );
  AOI22_X1 U658 ( .A1(n847), .A2(\REGISTERS[1][17] ), .B1(n13), .B2(
        \REGISTERS[12][17] ), .ZN(n558) );
  NAND4_X1 U659 ( .A1(n561), .A2(n560), .A3(n559), .A4(n558), .ZN(n562) );
  NOR4_X1 U660 ( .A1(n565), .A2(n564), .A3(n563), .A4(n562), .ZN(n566) );
  AOI22_X1 U661 ( .A1(n33), .A2(n102), .B1(n566), .B2(n35), .ZN(N264) );
  AOI22_X1 U662 ( .A1(n859), .A2(\REGISTERS[6][18] ), .B1(n29), .B2(
        \REGISTERS[11][18] ), .ZN(n570) );
  AOI22_X1 U663 ( .A1(n883), .A2(\REGISTERS[13][18] ), .B1(n1), .B2(
        \REGISTERS[0][18] ), .ZN(n569) );
  AOI22_X1 U664 ( .A1(n871), .A2(\REGISTERS[5][18] ), .B1(n15), .B2(
        \REGISTERS[22][18] ), .ZN(n568) );
  AOI22_X1 U665 ( .A1(n14), .A2(\REGISTERS[29][18] ), .B1(n6), .B2(
        \REGISTERS[24][18] ), .ZN(n567) );
  NAND4_X1 U666 ( .A1(n570), .A2(n569), .A3(n568), .A4(n567), .ZN(n586) );
  AOI22_X1 U667 ( .A1(n28), .A2(\REGISTERS[30][18] ), .B1(n12), .B2(
        \REGISTERS[28][18] ), .ZN(n574) );
  AOI22_X1 U668 ( .A1(n865), .A2(\REGISTERS[14][18] ), .B1(n13), .B2(
        \REGISTERS[12][18] ), .ZN(n573) );
  AOI22_X1 U669 ( .A1(n867), .A2(\REGISTERS[8][18] ), .B1(n23), .B2(
        \REGISTERS[16][18] ), .ZN(n572) );
  AOI22_X1 U670 ( .A1(n841), .A2(\REGISTERS[23][18] ), .B1(n9), .B2(
        \REGISTERS[9][18] ), .ZN(n571) );
  NAND4_X1 U671 ( .A1(n574), .A2(n573), .A3(n572), .A4(n571), .ZN(n585) );
  AOI22_X1 U672 ( .A1(n854), .A2(\REGISTERS[3][18] ), .B1(n5), .B2(
        \REGISTERS[31][18] ), .ZN(n578) );
  AOI22_X1 U673 ( .A1(n31), .A2(\REGISTERS[10][18] ), .B1(n7), .B2(
        \REGISTERS[19][18] ), .ZN(n577) );
  AOI22_X1 U674 ( .A1(n26), .A2(\REGISTERS[7][18] ), .B1(n25), .B2(
        \REGISTERS[15][18] ), .ZN(n576) );
  AOI22_X1 U675 ( .A1(n27), .A2(\REGISTERS[26][18] ), .B1(n22), .B2(
        \REGISTERS[21][18] ), .ZN(n575) );
  NAND4_X1 U676 ( .A1(n578), .A2(n577), .A3(n576), .A4(n575), .ZN(n584) );
  AOI22_X1 U677 ( .A1(n864), .A2(\REGISTERS[20][18] ), .B1(n19), .B2(
        \REGISTERS[4][18] ), .ZN(n582) );
  AOI22_X1 U678 ( .A1(n30), .A2(\REGISTERS[25][18] ), .B1(n8), .B2(
        \REGISTERS[1][18] ), .ZN(n581) );
  AOI22_X1 U679 ( .A1(n853), .A2(\REGISTERS[17][18] ), .B1(n868), .B2(
        \REGISTERS[18][18] ), .ZN(n580) );
  AOI22_X1 U680 ( .A1(n4), .A2(\REGISTERS[27][18] ), .B1(n3), .B2(
        \REGISTERS[2][18] ), .ZN(n579) );
  NAND4_X1 U681 ( .A1(n582), .A2(n581), .A3(n580), .A4(n579), .ZN(n583) );
  NOR4_X1 U682 ( .A1(n586), .A2(n585), .A3(n584), .A4(n583), .ZN(n587) );
  AOI22_X1 U683 ( .A1(n33), .A2(n100), .B1(n587), .B2(n36), .ZN(N265) );
  AOI22_X1 U684 ( .A1(n26), .A2(\REGISTERS[7][19] ), .B1(n4), .B2(
        \REGISTERS[27][19] ), .ZN(n591) );
  AOI22_X1 U685 ( .A1(n865), .A2(\REGISTERS[14][19] ), .B1(n21), .B2(
        \REGISTERS[18][19] ), .ZN(n590) );
  AOI22_X1 U686 ( .A1(n867), .A2(\REGISTERS[8][19] ), .B1(n7), .B2(
        \REGISTERS[19][19] ), .ZN(n589) );
  AOI22_X1 U687 ( .A1(n28), .A2(\REGISTERS[30][19] ), .B1(n29), .B2(
        \REGISTERS[11][19] ), .ZN(n588) );
  NAND4_X1 U688 ( .A1(n591), .A2(n590), .A3(n589), .A4(n588), .ZN(n607) );
  AOI22_X1 U689 ( .A1(n883), .A2(\REGISTERS[13][19] ), .B1(n8), .B2(
        \REGISTERS[1][19] ), .ZN(n595) );
  AOI22_X1 U690 ( .A1(n30), .A2(\REGISTERS[25][19] ), .B1(n15), .B2(
        \REGISTERS[22][19] ), .ZN(n594) );
  AOI22_X1 U691 ( .A1(n866), .A2(\REGISTERS[4][19] ), .B1(n9), .B2(
        \REGISTERS[9][19] ), .ZN(n593) );
  AOI22_X1 U692 ( .A1(n876), .A2(\REGISTERS[15][19] ), .B1(n5), .B2(
        \REGISTERS[31][19] ), .ZN(n592) );
  NAND4_X1 U693 ( .A1(n595), .A2(n594), .A3(n593), .A4(n592), .ZN(n606) );
  AOI22_X1 U694 ( .A1(n882), .A2(\REGISTERS[10][19] ), .B1(n1), .B2(
        \REGISTERS[0][19] ), .ZN(n599) );
  AOI22_X1 U695 ( .A1(n853), .A2(\REGISTERS[17][19] ), .B1(n2), .B2(
        \REGISTERS[23][19] ), .ZN(n598) );
  AOI22_X1 U696 ( .A1(n869), .A2(\REGISTERS[21][19] ), .B1(n17), .B2(
        \REGISTERS[20][19] ), .ZN(n597) );
  AOI22_X1 U697 ( .A1(n11), .A2(\REGISTERS[3][19] ), .B1(n13), .B2(
        \REGISTERS[12][19] ), .ZN(n596) );
  NAND4_X1 U698 ( .A1(n599), .A2(n598), .A3(n597), .A4(n596), .ZN(n605) );
  AOI22_X1 U699 ( .A1(n878), .A2(\REGISTERS[26][19] ), .B1(n23), .B2(
        \REGISTERS[16][19] ), .ZN(n603) );
  AOI22_X1 U700 ( .A1(n845), .A2(\REGISTERS[24][19] ), .B1(n3), .B2(
        \REGISTERS[2][19] ), .ZN(n602) );
  AOI22_X1 U701 ( .A1(n857), .A2(\REGISTERS[29][19] ), .B1(n24), .B2(
        \REGISTERS[5][19] ), .ZN(n601) );
  AOI22_X1 U702 ( .A1(n855), .A2(\REGISTERS[28][19] ), .B1(n16), .B2(
        \REGISTERS[6][19] ), .ZN(n600) );
  NAND4_X1 U703 ( .A1(n603), .A2(n602), .A3(n601), .A4(n600), .ZN(n604) );
  NOR4_X1 U704 ( .A1(n607), .A2(n606), .A3(n605), .A4(n604), .ZN(n608) );
  AOI22_X1 U705 ( .A1(n33), .A2(n98), .B1(n608), .B2(n36), .ZN(N266) );
  AOI22_X1 U706 ( .A1(n878), .A2(\REGISTERS[26][20] ), .B1(n10), .B2(
        \REGISTERS[17][20] ), .ZN(n612) );
  AOI22_X1 U707 ( .A1(n869), .A2(\REGISTERS[21][20] ), .B1(n8), .B2(
        \REGISTERS[1][20] ), .ZN(n611) );
  AOI22_X1 U708 ( .A1(n26), .A2(\REGISTERS[7][20] ), .B1(n4), .B2(
        \REGISTERS[27][20] ), .ZN(n610) );
  AOI22_X1 U709 ( .A1(n879), .A2(\REGISTERS[30][20] ), .B1(n14), .B2(
        \REGISTERS[29][20] ), .ZN(n609) );
  NAND4_X1 U710 ( .A1(n612), .A2(n611), .A3(n610), .A4(n609), .ZN(n628) );
  AOI22_X1 U711 ( .A1(n882), .A2(\REGISTERS[10][20] ), .B1(n18), .B2(
        \REGISTERS[14][20] ), .ZN(n616) );
  AOI22_X1 U712 ( .A1(n854), .A2(\REGISTERS[3][20] ), .B1(n3), .B2(
        \REGISTERS[2][20] ), .ZN(n615) );
  AOI22_X1 U713 ( .A1(n841), .A2(\REGISTERS[23][20] ), .B1(n15), .B2(
        \REGISTERS[22][20] ), .ZN(n614) );
  AOI22_X1 U714 ( .A1(n846), .A2(\REGISTERS[19][20] ), .B1(n29), .B2(
        \REGISTERS[11][20] ), .ZN(n613) );
  NAND4_X1 U715 ( .A1(n616), .A2(n615), .A3(n614), .A4(n613), .ZN(n627) );
  AOI22_X1 U716 ( .A1(n881), .A2(\REGISTERS[25][20] ), .B1(n13), .B2(
        \REGISTERS[12][20] ), .ZN(n620) );
  AOI22_X1 U717 ( .A1(n25), .A2(\REGISTERS[15][20] ), .B1(n17), .B2(
        \REGISTERS[20][20] ), .ZN(n619) );
  AOI22_X1 U718 ( .A1(n859), .A2(\REGISTERS[6][20] ), .B1(n21), .B2(
        \REGISTERS[18][20] ), .ZN(n618) );
  AOI22_X1 U719 ( .A1(n883), .A2(\REGISTERS[13][20] ), .B1(n12), .B2(
        \REGISTERS[28][20] ), .ZN(n617) );
  NAND4_X1 U720 ( .A1(n620), .A2(n619), .A3(n618), .A4(n617), .ZN(n626) );
  AOI22_X1 U721 ( .A1(n867), .A2(\REGISTERS[8][20] ), .B1(n24), .B2(
        \REGISTERS[5][20] ), .ZN(n624) );
  AOI22_X1 U722 ( .A1(n866), .A2(\REGISTERS[4][20] ), .B1(n852), .B2(
        \REGISTERS[9][20] ), .ZN(n623) );
  AOI22_X1 U723 ( .A1(n1), .A2(\REGISTERS[0][20] ), .B1(n6), .B2(
        \REGISTERS[24][20] ), .ZN(n622) );
  AOI22_X1 U724 ( .A1(n870), .A2(\REGISTERS[16][20] ), .B1(n844), .B2(
        \REGISTERS[31][20] ), .ZN(n621) );
  NAND4_X1 U725 ( .A1(n624), .A2(n623), .A3(n622), .A4(n621), .ZN(n625) );
  NOR4_X1 U726 ( .A1(n628), .A2(n627), .A3(n626), .A4(n625), .ZN(n629) );
  AOI22_X1 U727 ( .A1(n33), .A2(n96), .B1(n629), .B2(n35), .ZN(N267) );
  AOI22_X1 U728 ( .A1(n854), .A2(\REGISTERS[3][21] ), .B1(n15), .B2(
        \REGISTERS[22][21] ), .ZN(n633) );
  AOI22_X1 U729 ( .A1(n856), .A2(\REGISTERS[12][21] ), .B1(n5), .B2(
        \REGISTERS[31][21] ), .ZN(n632) );
  AOI22_X1 U730 ( .A1(n857), .A2(\REGISTERS[29][21] ), .B1(n17), .B2(
        \REGISTERS[20][21] ), .ZN(n631) );
  AOI22_X1 U731 ( .A1(n855), .A2(\REGISTERS[28][21] ), .B1(n9), .B2(
        \REGISTERS[9][21] ), .ZN(n630) );
  NAND4_X1 U732 ( .A1(n633), .A2(n632), .A3(n631), .A4(n630), .ZN(n649) );
  AOI22_X1 U733 ( .A1(n20), .A2(\REGISTERS[8][21] ), .B1(n4), .B2(
        \REGISTERS[27][21] ), .ZN(n637) );
  AOI22_X1 U734 ( .A1(n869), .A2(\REGISTERS[21][21] ), .B1(n18), .B2(
        \REGISTERS[14][21] ), .ZN(n636) );
  AOI22_X1 U735 ( .A1(n846), .A2(\REGISTERS[19][21] ), .B1(n24), .B2(
        \REGISTERS[5][21] ), .ZN(n635) );
  AOI22_X1 U736 ( .A1(n26), .A2(\REGISTERS[7][21] ), .B1(n25), .B2(
        \REGISTERS[15][21] ), .ZN(n634) );
  NAND4_X1 U737 ( .A1(n637), .A2(n636), .A3(n635), .A4(n634), .ZN(n648) );
  AOI22_X1 U738 ( .A1(n881), .A2(\REGISTERS[25][21] ), .B1(n3), .B2(
        \REGISTERS[2][21] ), .ZN(n641) );
  AOI22_X1 U739 ( .A1(n879), .A2(\REGISTERS[30][21] ), .B1(n8), .B2(
        \REGISTERS[1][21] ), .ZN(n640) );
  AOI22_X1 U740 ( .A1(n883), .A2(\REGISTERS[13][21] ), .B1(n10), .B2(
        \REGISTERS[17][21] ), .ZN(n639) );
  AOI22_X1 U741 ( .A1(n840), .A2(\REGISTERS[0][21] ), .B1(n19), .B2(
        \REGISTERS[4][21] ), .ZN(n638) );
  NAND4_X1 U742 ( .A1(n641), .A2(n640), .A3(n639), .A4(n638), .ZN(n647) );
  AOI22_X1 U743 ( .A1(n882), .A2(\REGISTERS[10][21] ), .B1(n6), .B2(
        \REGISTERS[24][21] ), .ZN(n645) );
  AOI22_X1 U744 ( .A1(n16), .A2(\REGISTERS[6][21] ), .B1(n21), .B2(
        \REGISTERS[18][21] ), .ZN(n644) );
  AOI22_X1 U745 ( .A1(n878), .A2(\REGISTERS[26][21] ), .B1(n2), .B2(
        \REGISTERS[23][21] ), .ZN(n643) );
  AOI22_X1 U746 ( .A1(n880), .A2(\REGISTERS[11][21] ), .B1(n23), .B2(
        \REGISTERS[16][21] ), .ZN(n642) );
  NAND4_X1 U747 ( .A1(n645), .A2(n644), .A3(n643), .A4(n642), .ZN(n646) );
  NOR4_X1 U748 ( .A1(n649), .A2(n648), .A3(n647), .A4(n646), .ZN(n650) );
  AOI22_X1 U749 ( .A1(n33), .A2(n1781), .B1(n650), .B2(n36), .ZN(N268) );
  AOI22_X1 U750 ( .A1(n877), .A2(\REGISTERS[7][22] ), .B1(n16), .B2(
        \REGISTERS[6][22] ), .ZN(n654) );
  AOI22_X1 U751 ( .A1(n853), .A2(\REGISTERS[17][22] ), .B1(n4), .B2(
        \REGISTERS[27][22] ), .ZN(n653) );
  AOI22_X1 U752 ( .A1(n6), .A2(\REGISTERS[24][22] ), .B1(n24), .B2(
        \REGISTERS[5][22] ), .ZN(n652) );
  AOI22_X1 U753 ( .A1(n856), .A2(\REGISTERS[12][22] ), .B1(n844), .B2(
        \REGISTERS[31][22] ), .ZN(n651) );
  NAND4_X1 U754 ( .A1(n654), .A2(n653), .A3(n652), .A4(n651), .ZN(n670) );
  AOI22_X1 U755 ( .A1(n878), .A2(\REGISTERS[26][22] ), .B1(n32), .B2(
        \REGISTERS[13][22] ), .ZN(n658) );
  AOI22_X1 U756 ( .A1(n865), .A2(\REGISTERS[14][22] ), .B1(n11), .B2(
        \REGISTERS[3][22] ), .ZN(n657) );
  AOI22_X1 U757 ( .A1(n22), .A2(\REGISTERS[21][22] ), .B1(n21), .B2(
        \REGISTERS[18][22] ), .ZN(n656) );
  AOI22_X1 U758 ( .A1(n841), .A2(\REGISTERS[23][22] ), .B1(n19), .B2(
        \REGISTERS[4][22] ), .ZN(n655) );
  NAND4_X1 U759 ( .A1(n658), .A2(n657), .A3(n656), .A4(n655), .ZN(n669) );
  AOI22_X1 U760 ( .A1(n842), .A2(\REGISTERS[2][22] ), .B1(n29), .B2(
        \REGISTERS[11][22] ), .ZN(n662) );
  AOI22_X1 U761 ( .A1(n881), .A2(\REGISTERS[25][22] ), .B1(n31), .B2(
        \REGISTERS[10][22] ), .ZN(n661) );
  AOI22_X1 U762 ( .A1(n879), .A2(\REGISTERS[30][22] ), .B1(n25), .B2(
        \REGISTERS[15][22] ), .ZN(n660) );
  AOI22_X1 U763 ( .A1(n867), .A2(\REGISTERS[8][22] ), .B1(n17), .B2(
        \REGISTERS[20][22] ), .ZN(n659) );
  NAND4_X1 U764 ( .A1(n662), .A2(n661), .A3(n660), .A4(n659), .ZN(n668) );
  AOI22_X1 U765 ( .A1(n857), .A2(\REGISTERS[29][22] ), .B1(n7), .B2(
        \REGISTERS[19][22] ), .ZN(n666) );
  AOI22_X1 U766 ( .A1(n870), .A2(\REGISTERS[16][22] ), .B1(n852), .B2(
        \REGISTERS[9][22] ), .ZN(n665) );
  AOI22_X1 U767 ( .A1(n840), .A2(\REGISTERS[0][22] ), .B1(n858), .B2(
        \REGISTERS[22][22] ), .ZN(n664) );
  AOI22_X1 U768 ( .A1(n855), .A2(\REGISTERS[28][22] ), .B1(n847), .B2(
        \REGISTERS[1][22] ), .ZN(n663) );
  NAND4_X1 U769 ( .A1(n666), .A2(n665), .A3(n664), .A4(n663), .ZN(n667) );
  NOR4_X1 U770 ( .A1(n670), .A2(n669), .A3(n668), .A4(n667), .ZN(n671) );
  AOI22_X1 U771 ( .A1(n33), .A2(n92), .B1(n671), .B2(n36), .ZN(N269) );
  AOI22_X1 U772 ( .A1(n18), .A2(\REGISTERS[14][23] ), .B1(n24), .B2(
        \REGISTERS[5][23] ), .ZN(n675) );
  AOI22_X1 U773 ( .A1(n877), .A2(\REGISTERS[7][23] ), .B1(n27), .B2(
        \REGISTERS[26][23] ), .ZN(n674) );
  AOI22_X1 U774 ( .A1(n881), .A2(\REGISTERS[25][23] ), .B1(n7), .B2(
        \REGISTERS[19][23] ), .ZN(n673) );
  AOI22_X1 U775 ( .A1(n840), .A2(\REGISTERS[0][23] ), .B1(n17), .B2(
        \REGISTERS[20][23] ), .ZN(n672) );
  NAND4_X1 U776 ( .A1(n675), .A2(n674), .A3(n673), .A4(n672), .ZN(n691) );
  AOI22_X1 U777 ( .A1(n845), .A2(\REGISTERS[24][23] ), .B1(n852), .B2(
        \REGISTERS[9][23] ), .ZN(n679) );
  AOI22_X1 U778 ( .A1(n20), .A2(\REGISTERS[8][23] ), .B1(n844), .B2(
        \REGISTERS[31][23] ), .ZN(n678) );
  AOI22_X1 U779 ( .A1(n8), .A2(\REGISTERS[1][23] ), .B1(n21), .B2(
        \REGISTERS[18][23] ), .ZN(n677) );
  AOI22_X1 U780 ( .A1(n843), .A2(\REGISTERS[27][23] ), .B1(n11), .B2(
        \REGISTERS[3][23] ), .ZN(n676) );
  NAND4_X1 U781 ( .A1(n679), .A2(n678), .A3(n677), .A4(n676), .ZN(n690) );
  AOI22_X1 U782 ( .A1(n841), .A2(\REGISTERS[23][23] ), .B1(n870), .B2(
        \REGISTERS[16][23] ), .ZN(n683) );
  AOI22_X1 U783 ( .A1(n855), .A2(\REGISTERS[28][23] ), .B1(n25), .B2(
        \REGISTERS[15][23] ), .ZN(n682) );
  AOI22_X1 U784 ( .A1(n880), .A2(\REGISTERS[11][23] ), .B1(n858), .B2(
        \REGISTERS[22][23] ), .ZN(n681) );
  AOI22_X1 U785 ( .A1(n857), .A2(\REGISTERS[29][23] ), .B1(n19), .B2(
        \REGISTERS[4][23] ), .ZN(n680) );
  NAND4_X1 U786 ( .A1(n683), .A2(n682), .A3(n681), .A4(n680), .ZN(n689) );
  AOI22_X1 U787 ( .A1(n859), .A2(\REGISTERS[6][23] ), .B1(n13), .B2(
        \REGISTERS[12][23] ), .ZN(n687) );
  AOI22_X1 U788 ( .A1(n10), .A2(\REGISTERS[17][23] ), .B1(n3), .B2(
        \REGISTERS[2][23] ), .ZN(n686) );
  AOI22_X1 U789 ( .A1(n879), .A2(\REGISTERS[30][23] ), .B1(n31), .B2(
        \REGISTERS[10][23] ), .ZN(n685) );
  AOI22_X1 U790 ( .A1(n883), .A2(\REGISTERS[13][23] ), .B1(n22), .B2(
        \REGISTERS[21][23] ), .ZN(n684) );
  NAND4_X1 U791 ( .A1(n687), .A2(n686), .A3(n685), .A4(n684), .ZN(n688) );
  NOR4_X1 U792 ( .A1(n691), .A2(n690), .A3(n689), .A4(n688), .ZN(n692) );
  AOI22_X1 U793 ( .A1(n33), .A2(n90), .B1(n692), .B2(n36), .ZN(N270) );
  AOI22_X1 U794 ( .A1(n867), .A2(\REGISTERS[8][24] ), .B1(n3), .B2(
        \REGISTERS[2][24] ), .ZN(n696) );
  AOI22_X1 U795 ( .A1(n881), .A2(\REGISTERS[25][24] ), .B1(n18), .B2(
        \REGISTERS[14][24] ), .ZN(n695) );
  AOI22_X1 U796 ( .A1(n853), .A2(\REGISTERS[17][24] ), .B1(n4), .B2(
        \REGISTERS[27][24] ), .ZN(n694) );
  AOI22_X1 U797 ( .A1(n879), .A2(\REGISTERS[30][24] ), .B1(n27), .B2(
        \REGISTERS[26][24] ), .ZN(n693) );
  NAND4_X1 U798 ( .A1(n696), .A2(n695), .A3(n694), .A4(n693), .ZN(n712) );
  AOI22_X1 U799 ( .A1(n856), .A2(\REGISTERS[12][24] ), .B1(n5), .B2(
        \REGISTERS[31][24] ), .ZN(n700) );
  AOI22_X1 U800 ( .A1(n871), .A2(\REGISTERS[5][24] ), .B1(n870), .B2(
        \REGISTERS[16][24] ), .ZN(n699) );
  AOI22_X1 U801 ( .A1(n26), .A2(\REGISTERS[7][24] ), .B1(n858), .B2(
        \REGISTERS[22][24] ), .ZN(n698) );
  AOI22_X1 U802 ( .A1(n882), .A2(\REGISTERS[10][24] ), .B1(n8), .B2(
        \REGISTERS[1][24] ), .ZN(n697) );
  NAND4_X1 U803 ( .A1(n700), .A2(n699), .A3(n698), .A4(n697), .ZN(n711) );
  AOI22_X1 U804 ( .A1(n869), .A2(\REGISTERS[21][24] ), .B1(n11), .B2(
        \REGISTERS[3][24] ), .ZN(n704) );
  AOI22_X1 U805 ( .A1(n841), .A2(\REGISTERS[23][24] ), .B1(n7), .B2(
        \REGISTERS[19][24] ), .ZN(n703) );
  AOI22_X1 U806 ( .A1(n857), .A2(\REGISTERS[29][24] ), .B1(n21), .B2(
        \REGISTERS[18][24] ), .ZN(n702) );
  AOI22_X1 U807 ( .A1(n880), .A2(\REGISTERS[11][24] ), .B1(n9), .B2(
        \REGISTERS[9][24] ), .ZN(n701) );
  NAND4_X1 U808 ( .A1(n704), .A2(n703), .A3(n702), .A4(n701), .ZN(n710) );
  AOI22_X1 U809 ( .A1(n864), .A2(\REGISTERS[20][24] ), .B1(n6), .B2(
        \REGISTERS[24][24] ), .ZN(n708) );
  AOI22_X1 U810 ( .A1(n876), .A2(\REGISTERS[15][24] ), .B1(n1), .B2(
        \REGISTERS[0][24] ), .ZN(n707) );
  AOI22_X1 U811 ( .A1(n883), .A2(\REGISTERS[13][24] ), .B1(n19), .B2(
        \REGISTERS[4][24] ), .ZN(n706) );
  AOI22_X1 U812 ( .A1(n855), .A2(\REGISTERS[28][24] ), .B1(n16), .B2(
        \REGISTERS[6][24] ), .ZN(n705) );
  NAND4_X1 U813 ( .A1(n708), .A2(n707), .A3(n706), .A4(n705), .ZN(n709) );
  NOR4_X1 U814 ( .A1(n712), .A2(n711), .A3(n710), .A4(n709), .ZN(n713) );
  AOI22_X1 U815 ( .A1(n34), .A2(n1780), .B1(n713), .B2(n36), .ZN(N271) );
  AOI22_X1 U816 ( .A1(n2), .A2(\REGISTERS[23][25] ), .B1(n24), .B2(
        \REGISTERS[5][25] ), .ZN(n717) );
  AOI22_X1 U817 ( .A1(n879), .A2(\REGISTERS[30][25] ), .B1(n29), .B2(
        \REGISTERS[11][25] ), .ZN(n716) );
  AOI22_X1 U818 ( .A1(n12), .A2(\REGISTERS[28][25] ), .B1(n20), .B2(
        \REGISTERS[8][25] ), .ZN(n715) );
  AOI22_X1 U819 ( .A1(n25), .A2(\REGISTERS[15][25] ), .B1(n7), .B2(
        \REGISTERS[19][25] ), .ZN(n714) );
  NAND4_X1 U820 ( .A1(n717), .A2(n716), .A3(n715), .A4(n714), .ZN(n733) );
  AOI22_X1 U821 ( .A1(n10), .A2(\REGISTERS[17][25] ), .B1(n21), .B2(
        \REGISTERS[18][25] ), .ZN(n721) );
  AOI22_X1 U822 ( .A1(n878), .A2(\REGISTERS[26][25] ), .B1(n6), .B2(
        \REGISTERS[24][25] ), .ZN(n720) );
  AOI22_X1 U823 ( .A1(n856), .A2(\REGISTERS[12][25] ), .B1(n9), .B2(
        \REGISTERS[9][25] ), .ZN(n719) );
  AOI22_X1 U824 ( .A1(n1), .A2(\REGISTERS[0][25] ), .B1(n5), .B2(
        \REGISTERS[31][25] ), .ZN(n718) );
  NAND4_X1 U825 ( .A1(n721), .A2(n720), .A3(n719), .A4(n718), .ZN(n732) );
  AOI22_X1 U826 ( .A1(n865), .A2(\REGISTERS[14][25] ), .B1(n4), .B2(
        \REGISTERS[27][25] ), .ZN(n725) );
  AOI22_X1 U827 ( .A1(n881), .A2(\REGISTERS[25][25] ), .B1(n11), .B2(
        \REGISTERS[3][25] ), .ZN(n724) );
  AOI22_X1 U828 ( .A1(n882), .A2(\REGISTERS[10][25] ), .B1(n19), .B2(
        \REGISTERS[4][25] ), .ZN(n723) );
  AOI22_X1 U829 ( .A1(n842), .A2(\REGISTERS[2][25] ), .B1(n858), .B2(
        \REGISTERS[22][25] ), .ZN(n722) );
  NAND4_X1 U830 ( .A1(n725), .A2(n724), .A3(n723), .A4(n722), .ZN(n731) );
  AOI22_X1 U831 ( .A1(n857), .A2(\REGISTERS[29][25] ), .B1(n17), .B2(
        \REGISTERS[20][25] ), .ZN(n729) );
  AOI22_X1 U832 ( .A1(n26), .A2(\REGISTERS[7][25] ), .B1(n22), .B2(
        \REGISTERS[21][25] ), .ZN(n728) );
  AOI22_X1 U833 ( .A1(n883), .A2(\REGISTERS[13][25] ), .B1(n16), .B2(
        \REGISTERS[6][25] ), .ZN(n727) );
  AOI22_X1 U834 ( .A1(n847), .A2(\REGISTERS[1][25] ), .B1(n870), .B2(
        \REGISTERS[16][25] ), .ZN(n726) );
  NAND4_X1 U835 ( .A1(n729), .A2(n728), .A3(n727), .A4(n726), .ZN(n730) );
  NOR4_X1 U836 ( .A1(n733), .A2(n732), .A3(n731), .A4(n730), .ZN(n734) );
  AOI22_X1 U837 ( .A1(n34), .A2(n86), .B1(n734), .B2(n35), .ZN(N272) );
  AOI22_X1 U838 ( .A1(n14), .A2(\REGISTERS[29][26] ), .B1(n870), .B2(
        \REGISTERS[16][26] ), .ZN(n738) );
  AOI22_X1 U839 ( .A1(n6), .A2(\REGISTERS[24][26] ), .B1(n858), .B2(
        \REGISTERS[22][26] ), .ZN(n737) );
  AOI22_X1 U840 ( .A1(n855), .A2(\REGISTERS[28][26] ), .B1(n29), .B2(
        \REGISTERS[11][26] ), .ZN(n736) );
  AOI22_X1 U841 ( .A1(n18), .A2(\REGISTERS[14][26] ), .B1(n5), .B2(
        \REGISTERS[31][26] ), .ZN(n735) );
  NAND4_X1 U842 ( .A1(n738), .A2(n737), .A3(n736), .A4(n735), .ZN(n754) );
  AOI22_X1 U843 ( .A1(n8), .A2(\REGISTERS[1][26] ), .B1(n13), .B2(
        \REGISTERS[12][26] ), .ZN(n742) );
  AOI22_X1 U844 ( .A1(n864), .A2(\REGISTERS[20][26] ), .B1(n9), .B2(
        \REGISTERS[9][26] ), .ZN(n741) );
  AOI22_X1 U845 ( .A1(n30), .A2(\REGISTERS[25][26] ), .B1(n3), .B2(
        \REGISTERS[2][26] ), .ZN(n740) );
  AOI22_X1 U846 ( .A1(n32), .A2(\REGISTERS[13][26] ), .B1(n846), .B2(
        \REGISTERS[19][26] ), .ZN(n739) );
  NAND4_X1 U847 ( .A1(n742), .A2(n741), .A3(n740), .A4(n739), .ZN(n753) );
  AOI22_X1 U848 ( .A1(n26), .A2(\REGISTERS[7][26] ), .B1(n11), .B2(
        \REGISTERS[3][26] ), .ZN(n746) );
  AOI22_X1 U849 ( .A1(n841), .A2(\REGISTERS[23][26] ), .B1(n24), .B2(
        \REGISTERS[5][26] ), .ZN(n745) );
  AOI22_X1 U850 ( .A1(n31), .A2(\REGISTERS[10][26] ), .B1(n19), .B2(
        \REGISTERS[4][26] ), .ZN(n744) );
  AOI22_X1 U851 ( .A1(n876), .A2(\REGISTERS[15][26] ), .B1(n4), .B2(
        \REGISTERS[27][26] ), .ZN(n743) );
  NAND4_X1 U852 ( .A1(n746), .A2(n745), .A3(n744), .A4(n743), .ZN(n752) );
  AOI22_X1 U853 ( .A1(n879), .A2(\REGISTERS[30][26] ), .B1(n1), .B2(
        \REGISTERS[0][26] ), .ZN(n750) );
  AOI22_X1 U854 ( .A1(n878), .A2(\REGISTERS[26][26] ), .B1(n16), .B2(
        \REGISTERS[6][26] ), .ZN(n749) );
  AOI22_X1 U855 ( .A1(n22), .A2(\REGISTERS[21][26] ), .B1(n20), .B2(
        \REGISTERS[8][26] ), .ZN(n748) );
  AOI22_X1 U856 ( .A1(n853), .A2(\REGISTERS[17][26] ), .B1(n21), .B2(
        \REGISTERS[18][26] ), .ZN(n747) );
  NAND4_X1 U857 ( .A1(n750), .A2(n749), .A3(n748), .A4(n747), .ZN(n751) );
  NOR4_X1 U858 ( .A1(n754), .A2(n753), .A3(n752), .A4(n751), .ZN(n755) );
  AOI22_X1 U859 ( .A1(n34), .A2(n84), .B1(n755), .B2(n35), .ZN(N273) );
  AOI22_X1 U860 ( .A1(n27), .A2(\REGISTERS[26][27] ), .B1(n8), .B2(
        \REGISTERS[1][27] ), .ZN(n759) );
  AOI22_X1 U861 ( .A1(n26), .A2(\REGISTERS[7][27] ), .B1(n10), .B2(
        \REGISTERS[17][27] ), .ZN(n758) );
  AOI22_X1 U862 ( .A1(n868), .A2(\REGISTERS[18][27] ), .B1(n871), .B2(
        \REGISTERS[5][27] ), .ZN(n757) );
  AOI22_X1 U863 ( .A1(n2), .A2(\REGISTERS[23][27] ), .B1(n842), .B2(
        \REGISTERS[2][27] ), .ZN(n756) );
  NAND4_X1 U864 ( .A1(n759), .A2(n758), .A3(n757), .A4(n756), .ZN(n775) );
  AOI22_X1 U865 ( .A1(n882), .A2(\REGISTERS[10][27] ), .B1(n15), .B2(
        \REGISTERS[22][27] ), .ZN(n763) );
  AOI22_X1 U866 ( .A1(n846), .A2(\REGISTERS[19][27] ), .B1(n856), .B2(
        \REGISTERS[12][27] ), .ZN(n762) );
  AOI22_X1 U867 ( .A1(n857), .A2(\REGISTERS[29][27] ), .B1(n880), .B2(
        \REGISTERS[11][27] ), .ZN(n761) );
  AOI22_X1 U868 ( .A1(n845), .A2(\REGISTERS[24][27] ), .B1(n9), .B2(
        \REGISTERS[9][27] ), .ZN(n760) );
  NAND4_X1 U869 ( .A1(n763), .A2(n762), .A3(n761), .A4(n760), .ZN(n774) );
  AOI22_X1 U870 ( .A1(n883), .A2(\REGISTERS[13][27] ), .B1(n17), .B2(
        \REGISTERS[20][27] ), .ZN(n767) );
  AOI22_X1 U871 ( .A1(n854), .A2(\REGISTERS[3][27] ), .B1(n5), .B2(
        \REGISTERS[31][27] ), .ZN(n766) );
  AOI22_X1 U872 ( .A1(n12), .A2(\REGISTERS[28][27] ), .B1(n25), .B2(
        \REGISTERS[15][27] ), .ZN(n765) );
  AOI22_X1 U873 ( .A1(n28), .A2(\REGISTERS[30][27] ), .B1(n18), .B2(
        \REGISTERS[14][27] ), .ZN(n764) );
  NAND4_X1 U874 ( .A1(n767), .A2(n766), .A3(n765), .A4(n764), .ZN(n773) );
  AOI22_X1 U875 ( .A1(n16), .A2(\REGISTERS[6][27] ), .B1(n4), .B2(
        \REGISTERS[27][27] ), .ZN(n771) );
  AOI22_X1 U876 ( .A1(n866), .A2(\REGISTERS[4][27] ), .B1(n23), .B2(
        \REGISTERS[16][27] ), .ZN(n770) );
  AOI22_X1 U877 ( .A1(n881), .A2(\REGISTERS[25][27] ), .B1(n1), .B2(
        \REGISTERS[0][27] ), .ZN(n769) );
  AOI22_X1 U878 ( .A1(n869), .A2(\REGISTERS[21][27] ), .B1(n20), .B2(
        \REGISTERS[8][27] ), .ZN(n768) );
  NAND4_X1 U879 ( .A1(n771), .A2(n770), .A3(n769), .A4(n768), .ZN(n772) );
  NOR4_X1 U880 ( .A1(n775), .A2(n774), .A3(n773), .A4(n772), .ZN(n776) );
  AOI22_X1 U881 ( .A1(n34), .A2(n1779), .B1(n776), .B2(n35), .ZN(N274) );
  AOI22_X1 U882 ( .A1(n32), .A2(\REGISTERS[13][28] ), .B1(n868), .B2(
        \REGISTERS[18][28] ), .ZN(n780) );
  AOI22_X1 U883 ( .A1(n840), .A2(\REGISTERS[0][28] ), .B1(n870), .B2(
        \REGISTERS[16][28] ), .ZN(n779) );
  AOI22_X1 U884 ( .A1(n6), .A2(\REGISTERS[24][28] ), .B1(n858), .B2(
        \REGISTERS[22][28] ), .ZN(n778) );
  AOI22_X1 U885 ( .A1(n4), .A2(\REGISTERS[27][28] ), .B1(n17), .B2(
        \REGISTERS[20][28] ), .ZN(n777) );
  NAND4_X1 U886 ( .A1(n780), .A2(n779), .A3(n778), .A4(n777), .ZN(n796) );
  AOI22_X1 U887 ( .A1(n22), .A2(\REGISTERS[21][28] ), .B1(n19), .B2(
        \REGISTERS[4][28] ), .ZN(n784) );
  AOI22_X1 U888 ( .A1(n859), .A2(\REGISTERS[6][28] ), .B1(n5), .B2(
        \REGISTERS[31][28] ), .ZN(n783) );
  AOI22_X1 U889 ( .A1(n31), .A2(\REGISTERS[10][28] ), .B1(n20), .B2(
        \REGISTERS[8][28] ), .ZN(n782) );
  AOI22_X1 U890 ( .A1(n25), .A2(\REGISTERS[15][28] ), .B1(n13), .B2(
        \REGISTERS[12][28] ), .ZN(n781) );
  NAND4_X1 U891 ( .A1(n784), .A2(n783), .A3(n782), .A4(n781), .ZN(n795) );
  AOI22_X1 U892 ( .A1(n26), .A2(\REGISTERS[7][28] ), .B1(n9), .B2(
        \REGISTERS[9][28] ), .ZN(n788) );
  AOI22_X1 U893 ( .A1(n847), .A2(\REGISTERS[1][28] ), .B1(n3), .B2(
        \REGISTERS[2][28] ), .ZN(n787) );
  AOI22_X1 U894 ( .A1(n865), .A2(\REGISTERS[14][28] ), .B1(n2), .B2(
        \REGISTERS[23][28] ), .ZN(n786) );
  AOI22_X1 U895 ( .A1(n14), .A2(\REGISTERS[29][28] ), .B1(n7), .B2(
        \REGISTERS[19][28] ), .ZN(n785) );
  NAND4_X1 U896 ( .A1(n788), .A2(n787), .A3(n786), .A4(n785), .ZN(n794) );
  AOI22_X1 U897 ( .A1(n879), .A2(\REGISTERS[30][28] ), .B1(n11), .B2(
        \REGISTERS[3][28] ), .ZN(n792) );
  AOI22_X1 U898 ( .A1(n855), .A2(\REGISTERS[28][28] ), .B1(n29), .B2(
        \REGISTERS[11][28] ), .ZN(n791) );
  AOI22_X1 U899 ( .A1(n10), .A2(\REGISTERS[17][28] ), .B1(n24), .B2(
        \REGISTERS[5][28] ), .ZN(n790) );
  AOI22_X1 U900 ( .A1(n878), .A2(\REGISTERS[26][28] ), .B1(n30), .B2(
        \REGISTERS[25][28] ), .ZN(n789) );
  NAND4_X1 U901 ( .A1(n792), .A2(n791), .A3(n790), .A4(n789), .ZN(n793) );
  NOR4_X1 U902 ( .A1(n796), .A2(n795), .A3(n794), .A4(n793), .ZN(n797) );
  AOI22_X1 U903 ( .A1(n34), .A2(n80), .B1(n797), .B2(n35), .ZN(N275) );
  AOI22_X1 U904 ( .A1(n845), .A2(\REGISTERS[24][29] ), .B1(n24), .B2(
        \REGISTERS[5][29] ), .ZN(n801) );
  AOI22_X1 U905 ( .A1(n30), .A2(\REGISTERS[25][29] ), .B1(n8), .B2(
        \REGISTERS[1][29] ), .ZN(n800) );
  AOI22_X1 U906 ( .A1(n853), .A2(\REGISTERS[17][29] ), .B1(n23), .B2(
        \REGISTERS[16][29] ), .ZN(n799) );
  AOI22_X1 U907 ( .A1(n20), .A2(\REGISTERS[8][29] ), .B1(n9), .B2(
        \REGISTERS[9][29] ), .ZN(n798) );
  NAND4_X1 U908 ( .A1(n801), .A2(n800), .A3(n799), .A4(n798), .ZN(n817) );
  AOI22_X1 U909 ( .A1(n876), .A2(\REGISTERS[15][29] ), .B1(n1), .B2(
        \REGISTERS[0][29] ), .ZN(n805) );
  AOI22_X1 U910 ( .A1(n12), .A2(\REGISTERS[28][29] ), .B1(n880), .B2(
        \REGISTERS[11][29] ), .ZN(n804) );
  AOI22_X1 U911 ( .A1(n16), .A2(\REGISTERS[6][29] ), .B1(n13), .B2(
        \REGISTERS[12][29] ), .ZN(n803) );
  AOI22_X1 U912 ( .A1(n846), .A2(\REGISTERS[19][29] ), .B1(n19), .B2(
        \REGISTERS[4][29] ), .ZN(n802) );
  NAND4_X1 U913 ( .A1(n805), .A2(n804), .A3(n803), .A4(n802), .ZN(n816) );
  AOI22_X1 U914 ( .A1(n882), .A2(\REGISTERS[10][29] ), .B1(n15), .B2(
        \REGISTERS[22][29] ), .ZN(n809) );
  AOI22_X1 U915 ( .A1(n26), .A2(\REGISTERS[7][29] ), .B1(n22), .B2(
        \REGISTERS[21][29] ), .ZN(n808) );
  AOI22_X1 U916 ( .A1(n883), .A2(\REGISTERS[13][29] ), .B1(n11), .B2(
        \REGISTERS[3][29] ), .ZN(n807) );
  AOI22_X1 U917 ( .A1(n28), .A2(\REGISTERS[30][29] ), .B1(n21), .B2(
        \REGISTERS[18][29] ), .ZN(n806) );
  NAND4_X1 U918 ( .A1(n809), .A2(n808), .A3(n807), .A4(n806), .ZN(n815) );
  AOI22_X1 U919 ( .A1(n27), .A2(\REGISTERS[26][29] ), .B1(n14), .B2(
        \REGISTERS[29][29] ), .ZN(n813) );
  AOI22_X1 U920 ( .A1(n18), .A2(\REGISTERS[14][29] ), .B1(n5), .B2(
        \REGISTERS[31][29] ), .ZN(n812) );
  AOI22_X1 U921 ( .A1(n843), .A2(\REGISTERS[27][29] ), .B1(n842), .B2(
        \REGISTERS[2][29] ), .ZN(n811) );
  AOI22_X1 U922 ( .A1(n841), .A2(\REGISTERS[23][29] ), .B1(n864), .B2(
        \REGISTERS[20][29] ), .ZN(n810) );
  NAND4_X1 U923 ( .A1(n813), .A2(n812), .A3(n811), .A4(n810), .ZN(n814) );
  NOR4_X1 U924 ( .A1(n817), .A2(n816), .A3(n815), .A4(n814), .ZN(n818) );
  AOI22_X1 U925 ( .A1(n34), .A2(n1777), .B1(n818), .B2(n35), .ZN(N276) );
  AOI22_X1 U926 ( .A1(n879), .A2(\REGISTERS[30][30] ), .B1(n856), .B2(
        \REGISTERS[12][30] ), .ZN(n822) );
  AOI22_X1 U927 ( .A1(n859), .A2(\REGISTERS[6][30] ), .B1(n871), .B2(
        \REGISTERS[5][30] ), .ZN(n821) );
  AOI22_X1 U928 ( .A1(n32), .A2(\REGISTERS[13][30] ), .B1(n8), .B2(
        \REGISTERS[1][30] ), .ZN(n820) );
  AOI22_X1 U929 ( .A1(n31), .A2(\REGISTERS[10][30] ), .B1(n858), .B2(
        \REGISTERS[22][30] ), .ZN(n819) );
  NAND4_X1 U930 ( .A1(n822), .A2(n821), .A3(n820), .A4(n819), .ZN(n838) );
  AOI22_X1 U931 ( .A1(n2), .A2(\REGISTERS[23][30] ), .B1(n5), .B2(
        \REGISTERS[31][30] ), .ZN(n826) );
  AOI22_X1 U932 ( .A1(n878), .A2(\REGISTERS[26][30] ), .B1(n870), .B2(
        \REGISTERS[16][30] ), .ZN(n825) );
  AOI22_X1 U933 ( .A1(n26), .A2(\REGISTERS[7][30] ), .B1(n19), .B2(
        \REGISTERS[4][30] ), .ZN(n824) );
  AOI22_X1 U934 ( .A1(n857), .A2(\REGISTERS[29][30] ), .B1(n7), .B2(
        \REGISTERS[19][30] ), .ZN(n823) );
  NAND4_X1 U935 ( .A1(n826), .A2(n825), .A3(n824), .A4(n823), .ZN(n837) );
  AOI22_X1 U936 ( .A1(n17), .A2(\REGISTERS[20][30] ), .B1(n6), .B2(
        \REGISTERS[24][30] ), .ZN(n830) );
  AOI22_X1 U937 ( .A1(n881), .A2(\REGISTERS[25][30] ), .B1(n25), .B2(
        \REGISTERS[15][30] ), .ZN(n829) );
  AOI22_X1 U938 ( .A1(n1), .A2(\REGISTERS[0][30] ), .B1(n868), .B2(
        \REGISTERS[18][30] ), .ZN(n828) );
  AOI22_X1 U939 ( .A1(n869), .A2(\REGISTERS[21][30] ), .B1(n11), .B2(
        \REGISTERS[3][30] ), .ZN(n827) );
  NAND4_X1 U940 ( .A1(n830), .A2(n829), .A3(n828), .A4(n827), .ZN(n836) );
  AOI22_X1 U941 ( .A1(n867), .A2(\REGISTERS[8][30] ), .B1(n29), .B2(
        \REGISTERS[11][30] ), .ZN(n834) );
  AOI22_X1 U942 ( .A1(n865), .A2(\REGISTERS[14][30] ), .B1(n4), .B2(
        \REGISTERS[27][30] ), .ZN(n833) );
  AOI22_X1 U943 ( .A1(n855), .A2(\REGISTERS[28][30] ), .B1(n10), .B2(
        \REGISTERS[17][30] ), .ZN(n832) );
  AOI22_X1 U944 ( .A1(n842), .A2(\REGISTERS[2][30] ), .B1(n9), .B2(
        \REGISTERS[9][30] ), .ZN(n831) );
  NAND4_X1 U945 ( .A1(n834), .A2(n833), .A3(n832), .A4(n831), .ZN(n835) );
  NOR4_X1 U946 ( .A1(n838), .A2(n837), .A3(n836), .A4(n835), .ZN(n839) );
  AOI22_X1 U947 ( .A1(n34), .A2(n76), .B1(n839), .B2(n35), .ZN(N277) );
  AOI22_X1 U948 ( .A1(n2), .A2(\REGISTERS[23][31] ), .B1(n1), .B2(
        \REGISTERS[0][31] ), .ZN(n851) );
  AOI22_X1 U949 ( .A1(n843), .A2(\REGISTERS[27][31] ), .B1(n3), .B2(
        \REGISTERS[2][31] ), .ZN(n850) );
  AOI22_X1 U950 ( .A1(n845), .A2(\REGISTERS[24][31] ), .B1(n5), .B2(
        \REGISTERS[31][31] ), .ZN(n849) );
  AOI22_X1 U951 ( .A1(n847), .A2(\REGISTERS[1][31] ), .B1(n7), .B2(
        \REGISTERS[19][31] ), .ZN(n848) );
  NAND4_X1 U952 ( .A1(n851), .A2(n850), .A3(n849), .A4(n848), .ZN(n891) );
  AOI22_X1 U953 ( .A1(n10), .A2(\REGISTERS[17][31] ), .B1(n9), .B2(
        \REGISTERS[9][31] ), .ZN(n863) );
  AOI22_X1 U954 ( .A1(n12), .A2(\REGISTERS[28][31] ), .B1(n11), .B2(
        \REGISTERS[3][31] ), .ZN(n862) );
  AOI22_X1 U955 ( .A1(n14), .A2(\REGISTERS[29][31] ), .B1(n13), .B2(
        \REGISTERS[12][31] ), .ZN(n861) );
  AOI22_X1 U956 ( .A1(n16), .A2(\REGISTERS[6][31] ), .B1(n15), .B2(
        \REGISTERS[22][31] ), .ZN(n860) );
  NAND4_X1 U957 ( .A1(n863), .A2(n862), .A3(n861), .A4(n860), .ZN(n890) );
  AOI22_X1 U958 ( .A1(n865), .A2(\REGISTERS[14][31] ), .B1(n17), .B2(
        \REGISTERS[20][31] ), .ZN(n875) );
  AOI22_X1 U959 ( .A1(n20), .A2(\REGISTERS[8][31] ), .B1(n866), .B2(
        \REGISTERS[4][31] ), .ZN(n874) );
  AOI22_X1 U960 ( .A1(n869), .A2(\REGISTERS[21][31] ), .B1(n21), .B2(
        \REGISTERS[18][31] ), .ZN(n873) );
  AOI22_X1 U961 ( .A1(n871), .A2(\REGISTERS[5][31] ), .B1(n23), .B2(
        \REGISTERS[16][31] ), .ZN(n872) );
  NAND4_X1 U962 ( .A1(n875), .A2(n874), .A3(n873), .A4(n872), .ZN(n889) );
  AOI22_X1 U963 ( .A1(n26), .A2(\REGISTERS[7][31] ), .B1(n25), .B2(
        \REGISTERS[15][31] ), .ZN(n887) );
  AOI22_X1 U964 ( .A1(n28), .A2(\REGISTERS[30][31] ), .B1(n27), .B2(
        \REGISTERS[26][31] ), .ZN(n886) );
  AOI22_X1 U965 ( .A1(n30), .A2(\REGISTERS[25][31] ), .B1(n29), .B2(
        \REGISTERS[11][31] ), .ZN(n885) );
  AOI22_X1 U966 ( .A1(n32), .A2(\REGISTERS[13][31] ), .B1(n31), .B2(
        \REGISTERS[10][31] ), .ZN(n884) );
  NAND4_X1 U967 ( .A1(n887), .A2(n886), .A3(n885), .A4(n884), .ZN(n888) );
  NOR4_X1 U968 ( .A1(n891), .A2(n890), .A3(n889), .A4(n888), .ZN(n892) );
  AOI22_X1 U969 ( .A1(n34), .A2(n74), .B1(n892), .B2(n35), .ZN(N278) );
  OAI221_X1 U970 ( .B1(ADD_WR[4]), .B2(n912), .C1(n894), .C2(ADD_RD2[4]), .A(
        WR), .ZN(n903) );
  AOI22_X1 U971 ( .A1(n897), .A2(ADD_RD2[3]), .B1(ADD_RD2[1]), .B2(n896), .ZN(
        n895) );
  OAI221_X1 U972 ( .B1(n897), .B2(ADD_RD2[3]), .C1(n896), .C2(ADD_RD2[1]), .A(
        n895), .ZN(n902) );
  AOI22_X1 U973 ( .A1(n900), .A2(ADD_RD2[2]), .B1(n899), .B2(ADD_RD2[0]), .ZN(
        n898) );
  OAI221_X1 U974 ( .B1(n900), .B2(ADD_RD2[2]), .C1(n899), .C2(ADD_RD2[0]), .A(
        n898), .ZN(n901) );
  INV_X1 U975 ( .A(ADD_RD2[2]), .ZN(n904) );
  NAND2_X1 U976 ( .A1(ADD_RD2[1]), .A2(n904), .ZN(n927) );
  INV_X1 U977 ( .A(ADD_RD2[3]), .ZN(n906) );
  NAND3_X1 U978 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[0]), .A3(n906), .ZN(n924) );
  NOR2_X1 U979 ( .A1(n927), .A2(n924), .ZN(n1603) );
  INV_X1 U980 ( .A(ADD_RD2[1]), .ZN(n905) );
  NAND2_X1 U981 ( .A1(n904), .A2(n905), .ZN(n930) );
  NAND3_X1 U982 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n912), .ZN(n919) );
  NOR2_X1 U983 ( .A1(n930), .A2(n919), .ZN(n1579) );
  AOI22_X1 U984 ( .A1(\REGISTERS[19][0] ), .A2(n58), .B1(\REGISTERS[9][0] ), 
        .B2(n42), .ZN(n911) );
  NAND2_X1 U985 ( .A1(ADD_RD2[2]), .A2(ADD_RD2[1]), .ZN(n925) );
  NOR2_X1 U986 ( .A1(n924), .A2(n925), .ZN(n1589) );
  NAND2_X1 U987 ( .A1(ADD_RD2[2]), .A2(n905), .ZN(n933) );
  NOR2_X1 U988 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .ZN(n907) );
  NAND2_X1 U989 ( .A1(ADD_RD2[4]), .A2(n907), .ZN(n929) );
  NOR2_X1 U990 ( .A1(n933), .A2(n929), .ZN(n1615) );
  AOI22_X1 U991 ( .A1(\REGISTERS[23][0] ), .A2(n48), .B1(\REGISTERS[20][0] ), 
        .B2(n66), .ZN(n910) );
  INV_X1 U992 ( .A(ADD_RD2[0]), .ZN(n913) );
  NAND3_X1 U993 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .A3(n913), .ZN(n931) );
  NOR2_X1 U994 ( .A1(n925), .A2(n931), .ZN(n1614) );
  NAND3_X1 U995 ( .A1(ADD_RD2[0]), .A2(n912), .A3(n906), .ZN(n932) );
  NOR2_X1 U996 ( .A1(n927), .A2(n932), .ZN(n1591) );
  AOI22_X1 U997 ( .A1(\REGISTERS[30][0] ), .A2(n65), .B1(\REGISTERS[3][0] ), 
        .B2(n50), .ZN(n909) );
  NAND2_X1 U998 ( .A1(n907), .A2(n912), .ZN(n928) );
  NOR2_X1 U999 ( .A1(n930), .A2(n928), .ZN(n1613) );
  NAND3_X1 U1000 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(ADD_RD2[3]), .ZN(n918) );
  NOR2_X1 U1001 ( .A1(n925), .A2(n918), .ZN(n1599) );
  AOI22_X1 U1002 ( .A1(\REGISTERS[0][0] ), .A2(n64), .B1(\REGISTERS[31][0] ), 
        .B2(n54), .ZN(n908) );
  NAND4_X1 U1003 ( .A1(n911), .A2(n910), .A3(n909), .A4(n908), .ZN(n941) );
  NOR2_X1 U1004 ( .A1(n927), .A2(n931), .ZN(n1602) );
  NAND3_X1 U1005 ( .A1(ADD_RD2[3]), .A2(n913), .A3(n912), .ZN(n926) );
  NOR2_X1 U1006 ( .A1(n927), .A2(n926), .ZN(n1578) );
  AOI22_X1 U1007 ( .A1(\REGISTERS[26][0] ), .A2(n57), .B1(\REGISTERS[10][0] ), 
        .B2(n41), .ZN(n917) );
  NOR2_X1 U1008 ( .A1(n925), .A2(n928), .ZN(n1616) );
  NOR2_X1 U1009 ( .A1(n925), .A2(n926), .ZN(n1581) );
  AOI22_X1 U1010 ( .A1(\REGISTERS[6][0] ), .A2(n67), .B1(\REGISTERS[14][0] ), 
        .B2(n44), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(n919), .A2(n933), .ZN(n1586) );
  NOR2_X1 U1012 ( .A1(n933), .A2(n918), .ZN(n1617) );
  AOI22_X1 U1013 ( .A1(\REGISTERS[13][0] ), .A2(n1586), .B1(\REGISTERS[29][0] ), .B2(n68), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(n930), .A2(n932), .ZN(n1576) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n927), .ZN(n1590) );
  AOI22_X1 U1016 ( .A1(\REGISTERS[1][0] ), .A2(n39), .B1(\REGISTERS[11][0] ), 
        .B2(n49), .ZN(n914) );
  NAND4_X1 U1017 ( .A1(n917), .A2(n916), .A3(n915), .A4(n914), .ZN(n940) );
  NOR2_X1 U1018 ( .A1(n930), .A2(n918), .ZN(n1610) );
  NOR2_X1 U1019 ( .A1(n927), .A2(n918), .ZN(n1577) );
  AOI22_X1 U1020 ( .A1(\REGISTERS[25][0] ), .A2(n1610), .B1(\REGISTERS[27][0] ), .B2(n40), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n925), .ZN(n1600) );
  NOR2_X1 U1022 ( .A1(n930), .A2(n931), .ZN(n1588) );
  AOI22_X1 U1023 ( .A1(\REGISTERS[15][0] ), .A2(n55), .B1(\REGISTERS[24][0] ), 
        .B2(n47), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n932), .ZN(n1580) );
  NOR2_X1 U1025 ( .A1(n930), .A2(n926), .ZN(n1575) );
  AOI22_X1 U1026 ( .A1(\REGISTERS[7][0] ), .A2(n1580), .B1(\REGISTERS[8][0] ), 
        .B2(n38), .ZN(n921) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n924), .ZN(n1593) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n929), .ZN(n1604) );
  AOI22_X1 U1029 ( .A1(\REGISTERS[17][0] ), .A2(n52), .B1(\REGISTERS[18][0] ), 
        .B2(n59), .ZN(n920) );
  NAND4_X1 U1030 ( .A1(n923), .A2(n922), .A3(n921), .A4(n920), .ZN(n939) );
  NOR2_X1 U1031 ( .A1(n924), .A2(n933), .ZN(n1598) );
  NOR2_X1 U1032 ( .A1(n925), .A2(n929), .ZN(n1592) );
  AOI22_X1 U1033 ( .A1(\REGISTERS[21][0] ), .A2(n53), .B1(\REGISTERS[22][0] ), 
        .B2(n51), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n926), .ZN(n1601) );
  NOR2_X1 U1035 ( .A1(n927), .A2(n928), .ZN(n1587) );
  AOI22_X1 U1036 ( .A1(\REGISTERS[12][0] ), .A2(n56), .B1(\REGISTERS[2][0] ), 
        .B2(n46), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n933), .A2(n928), .ZN(n1574) );
  NOR2_X1 U1038 ( .A1(n930), .A2(n929), .ZN(n1612) );
  AOI22_X1 U1039 ( .A1(\REGISTERS[4][0] ), .A2(n1574), .B1(\REGISTERS[16][0] ), 
        .B2(n63), .ZN(n935) );
  NOR2_X1 U1040 ( .A1(n933), .A2(n931), .ZN(n1605) );
  NOR2_X1 U1041 ( .A1(n933), .A2(n932), .ZN(n1611) );
  AOI22_X1 U1042 ( .A1(\REGISTERS[28][0] ), .A2(n60), .B1(\REGISTERS[5][0] ), 
        .B2(n62), .ZN(n934) );
  NAND4_X1 U1043 ( .A1(n937), .A2(n936), .A3(n935), .A4(n934), .ZN(n938) );
  NOR4_X1 U1044 ( .A1(n941), .A2(n940), .A3(n939), .A4(n938), .ZN(n942) );
  AOI22_X1 U1045 ( .A1(n69), .A2(n136), .B1(n942), .B2(n72), .ZN(N379) );
  AOI22_X1 U1046 ( .A1(\REGISTERS[3][1] ), .A2(n1591), .B1(\REGISTERS[28][1] ), 
        .B2(n60), .ZN(n946) );
  AOI22_X1 U1047 ( .A1(\REGISTERS[20][1] ), .A2(n1615), .B1(\REGISTERS[13][1] ), .B2(n45), .ZN(n945) );
  AOI22_X1 U1048 ( .A1(\REGISTERS[1][1] ), .A2(n1576), .B1(\REGISTERS[17][1] ), 
        .B2(n52), .ZN(n944) );
  AOI22_X1 U1049 ( .A1(\REGISTERS[18][1] ), .A2(n1604), .B1(\REGISTERS[6][1] ), 
        .B2(n67), .ZN(n943) );
  NAND4_X1 U1050 ( .A1(n946), .A2(n945), .A3(n944), .A4(n943), .ZN(n962) );
  AOI22_X1 U1051 ( .A1(\REGISTERS[12][1] ), .A2(n56), .B1(\REGISTERS[5][1] ), 
        .B2(n62), .ZN(n950) );
  AOI22_X1 U1052 ( .A1(\REGISTERS[24][1] ), .A2(n1588), .B1(\REGISTERS[30][1] ), .B2(n65), .ZN(n949) );
  AOI22_X1 U1053 ( .A1(\REGISTERS[4][1] ), .A2(n37), .B1(\REGISTERS[16][1] ), 
        .B2(n63), .ZN(n948) );
  AOI22_X1 U1054 ( .A1(\REGISTERS[27][1] ), .A2(n1577), .B1(\REGISTERS[0][1] ), 
        .B2(n64), .ZN(n947) );
  NAND4_X1 U1055 ( .A1(n950), .A2(n949), .A3(n948), .A4(n947), .ZN(n961) );
  AOI22_X1 U1056 ( .A1(\REGISTERS[26][1] ), .A2(n57), .B1(\REGISTERS[21][1] ), 
        .B2(n53), .ZN(n954) );
  AOI22_X1 U1057 ( .A1(\REGISTERS[14][1] ), .A2(n1581), .B1(\REGISTERS[11][1] ), .B2(n49), .ZN(n953) );
  AOI22_X1 U1058 ( .A1(\REGISTERS[8][1] ), .A2(n1575), .B1(\REGISTERS[15][1] ), 
        .B2(n55), .ZN(n952) );
  AOI22_X1 U1059 ( .A1(\REGISTERS[25][1] ), .A2(n1610), .B1(\REGISTERS[7][1] ), 
        .B2(n1580), .ZN(n951) );
  NAND4_X1 U1060 ( .A1(n954), .A2(n953), .A3(n952), .A4(n951), .ZN(n960) );
  AOI22_X1 U1061 ( .A1(\REGISTERS[23][1] ), .A2(n1589), .B1(\REGISTERS[19][1] ), .B2(n58), .ZN(n958) );
  AOI22_X1 U1062 ( .A1(\REGISTERS[22][1] ), .A2(n51), .B1(\REGISTERS[2][1] ), 
        .B2(n46), .ZN(n957) );
  AOI22_X1 U1063 ( .A1(\REGISTERS[10][1] ), .A2(n1578), .B1(\REGISTERS[29][1] ), .B2(n68), .ZN(n956) );
  AOI22_X1 U1064 ( .A1(\REGISTERS[9][1] ), .A2(n1579), .B1(\REGISTERS[31][1] ), 
        .B2(n54), .ZN(n955) );
  NAND4_X1 U1065 ( .A1(n958), .A2(n957), .A3(n956), .A4(n955), .ZN(n959) );
  NOR4_X1 U1066 ( .A1(n962), .A2(n961), .A3(n960), .A4(n959), .ZN(n963) );
  AOI22_X1 U1067 ( .A1(n70), .A2(n1778), .B1(n963), .B2(n71), .ZN(N380) );
  AOI22_X1 U1068 ( .A1(\REGISTERS[9][2] ), .A2(n42), .B1(\REGISTERS[10][2] ), 
        .B2(n41), .ZN(n967) );
  AOI22_X1 U1069 ( .A1(\REGISTERS[30][2] ), .A2(n65), .B1(\REGISTERS[3][2] ), 
        .B2(n50), .ZN(n966) );
  AOI22_X1 U1070 ( .A1(\REGISTERS[12][2] ), .A2(n1601), .B1(\REGISTERS[6][2] ), 
        .B2(n67), .ZN(n965) );
  AOI22_X1 U1071 ( .A1(\REGISTERS[22][2] ), .A2(n1592), .B1(\REGISTERS[15][2] ), .B2(n55), .ZN(n964) );
  NAND4_X1 U1072 ( .A1(n967), .A2(n966), .A3(n965), .A4(n964), .ZN(n983) );
  AOI22_X1 U1073 ( .A1(\REGISTERS[19][2] ), .A2(n1603), .B1(\REGISTERS[18][2] ), .B2(n59), .ZN(n971) );
  AOI22_X1 U1074 ( .A1(\REGISTERS[21][2] ), .A2(n1598), .B1(\REGISTERS[26][2] ), .B2(n57), .ZN(n970) );
  AOI22_X1 U1075 ( .A1(\REGISTERS[5][2] ), .A2(n62), .B1(\REGISTERS[8][2] ), 
        .B2(n38), .ZN(n969) );
  AOI22_X1 U1076 ( .A1(\REGISTERS[17][2] ), .A2(n1593), .B1(\REGISTERS[14][2] ), .B2(n44), .ZN(n968) );
  NAND4_X1 U1077 ( .A1(n971), .A2(n970), .A3(n969), .A4(n968), .ZN(n982) );
  AOI22_X1 U1078 ( .A1(\REGISTERS[28][2] ), .A2(n1605), .B1(\REGISTERS[7][2] ), 
        .B2(n1580), .ZN(n975) );
  AOI22_X1 U1079 ( .A1(\REGISTERS[16][2] ), .A2(n1612), .B1(\REGISTERS[31][2] ), .B2(n54), .ZN(n974) );
  AOI22_X1 U1080 ( .A1(\REGISTERS[24][2] ), .A2(n47), .B1(\REGISTERS[11][2] ), 
        .B2(n49), .ZN(n973) );
  AOI22_X1 U1081 ( .A1(\REGISTERS[0][2] ), .A2(n1613), .B1(\REGISTERS[2][2] ), 
        .B2(n46), .ZN(n972) );
  NAND4_X1 U1082 ( .A1(n975), .A2(n974), .A3(n973), .A4(n972), .ZN(n981) );
  AOI22_X1 U1083 ( .A1(\REGISTERS[25][2] ), .A2(n1610), .B1(\REGISTERS[4][2] ), 
        .B2(n37), .ZN(n979) );
  AOI22_X1 U1084 ( .A1(\REGISTERS[20][2] ), .A2(n1615), .B1(\REGISTERS[29][2] ), .B2(n68), .ZN(n978) );
  AOI22_X1 U1085 ( .A1(\REGISTERS[1][2] ), .A2(n1576), .B1(\REGISTERS[27][2] ), 
        .B2(n40), .ZN(n977) );
  AOI22_X1 U1086 ( .A1(\REGISTERS[23][2] ), .A2(n48), .B1(\REGISTERS[13][2] ), 
        .B2(n45), .ZN(n976) );
  NAND4_X1 U1087 ( .A1(n979), .A2(n978), .A3(n977), .A4(n976), .ZN(n980) );
  NOR4_X1 U1088 ( .A1(n983), .A2(n982), .A3(n981), .A4(n980), .ZN(n984) );
  AOI22_X1 U1089 ( .A1(n70), .A2(n132), .B1(n984), .B2(n72), .ZN(N381) );
  AOI22_X1 U1090 ( .A1(\REGISTERS[2][3] ), .A2(n46), .B1(\REGISTERS[12][3] ), 
        .B2(n56), .ZN(n988) );
  AOI22_X1 U1091 ( .A1(\REGISTERS[3][3] ), .A2(n50), .B1(\REGISTERS[8][3] ), 
        .B2(n38), .ZN(n987) );
  AOI22_X1 U1092 ( .A1(\REGISTERS[16][3] ), .A2(n63), .B1(\REGISTERS[31][3] ), 
        .B2(n54), .ZN(n986) );
  AOI22_X1 U1093 ( .A1(\REGISTERS[18][3] ), .A2(n1604), .B1(\REGISTERS[25][3] ), .B2(n61), .ZN(n985) );
  NAND4_X1 U1094 ( .A1(n988), .A2(n987), .A3(n986), .A4(n985), .ZN(n1004) );
  AOI22_X1 U1095 ( .A1(\REGISTERS[20][3] ), .A2(n66), .B1(\REGISTERS[26][3] ), 
        .B2(n57), .ZN(n992) );
  AOI22_X1 U1096 ( .A1(\REGISTERS[27][3] ), .A2(n1577), .B1(\REGISTERS[17][3] ), .B2(n52), .ZN(n991) );
  AOI22_X1 U1097 ( .A1(\REGISTERS[14][3] ), .A2(n44), .B1(\REGISTERS[23][3] ), 
        .B2(n48), .ZN(n990) );
  AOI22_X1 U1098 ( .A1(\REGISTERS[9][3] ), .A2(n1579), .B1(\REGISTERS[28][3] ), 
        .B2(n60), .ZN(n989) );
  NAND4_X1 U1099 ( .A1(n992), .A2(n991), .A3(n990), .A4(n989), .ZN(n1003) );
  AOI22_X1 U1100 ( .A1(\REGISTERS[30][3] ), .A2(n1614), .B1(\REGISTERS[5][3] ), 
        .B2(n62), .ZN(n996) );
  AOI22_X1 U1101 ( .A1(\REGISTERS[0][3] ), .A2(n1613), .B1(\REGISTERS[22][3] ), 
        .B2(n51), .ZN(n995) );
  AOI22_X1 U1102 ( .A1(\REGISTERS[15][3] ), .A2(n55), .B1(\REGISTERS[1][3] ), 
        .B2(n39), .ZN(n994) );
  AOI22_X1 U1103 ( .A1(\REGISTERS[21][3] ), .A2(n53), .B1(\REGISTERS[19][3] ), 
        .B2(n58), .ZN(n993) );
  NAND4_X1 U1104 ( .A1(n996), .A2(n995), .A3(n994), .A4(n993), .ZN(n1002) );
  AOI22_X1 U1105 ( .A1(\REGISTERS[4][3] ), .A2(n1574), .B1(\REGISTERS[7][3] ), 
        .B2(n43), .ZN(n1000) );
  AOI22_X1 U1106 ( .A1(\REGISTERS[10][3] ), .A2(n1578), .B1(\REGISTERS[24][3] ), .B2(n47), .ZN(n999) );
  AOI22_X1 U1107 ( .A1(\REGISTERS[29][3] ), .A2(n1617), .B1(\REGISTERS[13][3] ), .B2(n45), .ZN(n998) );
  AOI22_X1 U1108 ( .A1(\REGISTERS[11][3] ), .A2(n49), .B1(\REGISTERS[6][3] ), 
        .B2(n67), .ZN(n997) );
  NAND4_X1 U1109 ( .A1(n1000), .A2(n999), .A3(n998), .A4(n997), .ZN(n1001) );
  NOR4_X1 U1110 ( .A1(n1004), .A2(n1003), .A3(n1002), .A4(n1001), .ZN(n1005)
         );
  AOI22_X1 U1111 ( .A1(n70), .A2(n130), .B1(n1005), .B2(n71), .ZN(N382) );
  AOI22_X1 U1112 ( .A1(\REGISTERS[0][4] ), .A2(n64), .B1(\REGISTERS[30][4] ), 
        .B2(n65), .ZN(n1009) );
  AOI22_X1 U1113 ( .A1(\REGISTERS[18][4] ), .A2(n1604), .B1(\REGISTERS[9][4] ), 
        .B2(n42), .ZN(n1008) );
  AOI22_X1 U1114 ( .A1(\REGISTERS[3][4] ), .A2(n1591), .B1(\REGISTERS[7][4] ), 
        .B2(n43), .ZN(n1007) );
  AOI22_X1 U1115 ( .A1(\REGISTERS[26][4] ), .A2(n1602), .B1(\REGISTERS[19][4] ), .B2(n58), .ZN(n1006) );
  NAND4_X1 U1116 ( .A1(n1009), .A2(n1008), .A3(n1007), .A4(n1006), .ZN(n1026)
         );
  AOI22_X1 U1117 ( .A1(\REGISTERS[27][4] ), .A2(n40), .B1(\REGISTERS[8][4] ), 
        .B2(n38), .ZN(n1013) );
  AOI22_X1 U1118 ( .A1(\REGISTERS[1][4] ), .A2(n1576), .B1(\REGISTERS[10][4] ), 
        .B2(n41), .ZN(n1012) );
  AOI22_X1 U1119 ( .A1(\REGISTERS[25][4] ), .A2(n61), .B1(\REGISTERS[22][4] ), 
        .B2(n51), .ZN(n1011) );
  AOI22_X1 U1120 ( .A1(\REGISTERS[4][4] ), .A2(n37), .B1(\REGISTERS[20][4] ), 
        .B2(n66), .ZN(n1010) );
  NAND4_X1 U1121 ( .A1(n1013), .A2(n1012), .A3(n1011), .A4(n1010), .ZN(n1025)
         );
  AOI22_X1 U1122 ( .A1(\REGISTERS[28][4] ), .A2(n60), .B1(\REGISTERS[23][4] ), 
        .B2(n48), .ZN(n1017) );
  AOI22_X1 U1123 ( .A1(\REGISTERS[14][4] ), .A2(n1581), .B1(\REGISTERS[5][4] ), 
        .B2(n62), .ZN(n1016) );
  AOI22_X1 U1124 ( .A1(\REGISTERS[16][4] ), .A2(n1612), .B1(\REGISTERS[2][4] ), 
        .B2(n46), .ZN(n1015) );
  AOI22_X1 U1125 ( .A1(\REGISTERS[21][4] ), .A2(n1598), .B1(\REGISTERS[31][4] ), .B2(n54), .ZN(n1014) );
  NAND4_X1 U1126 ( .A1(n1017), .A2(n1016), .A3(n1015), .A4(n1014), .ZN(n1023)
         );
  AOI22_X1 U1127 ( .A1(\REGISTERS[29][4] ), .A2(n1617), .B1(\REGISTERS[24][4] ), .B2(n47), .ZN(n1021) );
  AOI22_X1 U1128 ( .A1(\REGISTERS[13][4] ), .A2(n1586), .B1(\REGISTERS[6][4] ), 
        .B2(n67), .ZN(n1020) );
  AOI22_X1 U1129 ( .A1(\REGISTERS[15][4] ), .A2(n1600), .B1(\REGISTERS[12][4] ), .B2(n56), .ZN(n1019) );
  AOI22_X1 U1130 ( .A1(\REGISTERS[11][4] ), .A2(n49), .B1(\REGISTERS[17][4] ), 
        .B2(n52), .ZN(n1018) );
  NAND4_X1 U1131 ( .A1(n1021), .A2(n1020), .A3(n1019), .A4(n1018), .ZN(n1022)
         );
  NOR4_X1 U1132 ( .A1(n1026), .A2(n1025), .A3(n1023), .A4(n1022), .ZN(n1027)
         );
  AOI22_X1 U1133 ( .A1(n70), .A2(n128), .B1(n1027), .B2(n72), .ZN(N383) );
  AOI22_X1 U1134 ( .A1(\REGISTERS[25][5] ), .A2(n61), .B1(\REGISTERS[16][5] ), 
        .B2(n63), .ZN(n1031) );
  AOI22_X1 U1135 ( .A1(\REGISTERS[14][5] ), .A2(n1581), .B1(\REGISTERS[12][5] ), .B2(n56), .ZN(n1030) );
  AOI22_X1 U1136 ( .A1(\REGISTERS[30][5] ), .A2(n1614), .B1(\REGISTERS[8][5] ), 
        .B2(n38), .ZN(n1029) );
  AOI22_X1 U1137 ( .A1(\REGISTERS[3][5] ), .A2(n50), .B1(\REGISTERS[0][5] ), 
        .B2(n64), .ZN(n1028) );
  NAND4_X1 U1138 ( .A1(n1031), .A2(n1030), .A3(n1029), .A4(n1028), .ZN(n1047)
         );
  AOI22_X1 U1139 ( .A1(\REGISTERS[20][5] ), .A2(n66), .B1(\REGISTERS[10][5] ), 
        .B2(n41), .ZN(n1035) );
  AOI22_X1 U1140 ( .A1(\REGISTERS[28][5] ), .A2(n1605), .B1(\REGISTERS[18][5] ), .B2(n59), .ZN(n1034) );
  AOI22_X1 U1141 ( .A1(\REGISTERS[17][5] ), .A2(n1593), .B1(\REGISTERS[5][5] ), 
        .B2(n62), .ZN(n1033) );
  AOI22_X1 U1142 ( .A1(\REGISTERS[13][5] ), .A2(n45), .B1(\REGISTERS[31][5] ), 
        .B2(n54), .ZN(n1032) );
  NAND4_X1 U1143 ( .A1(n1035), .A2(n1034), .A3(n1033), .A4(n1032), .ZN(n1046)
         );
  AOI22_X1 U1144 ( .A1(\REGISTERS[26][5] ), .A2(n1602), .B1(\REGISTERS[15][5] ), .B2(n55), .ZN(n1039) );
  AOI22_X1 U1145 ( .A1(\REGISTERS[11][5] ), .A2(n49), .B1(\REGISTERS[19][5] ), 
        .B2(n58), .ZN(n1038) );
  AOI22_X1 U1146 ( .A1(\REGISTERS[21][5] ), .A2(n53), .B1(\REGISTERS[6][5] ), 
        .B2(n67), .ZN(n1037) );
  AOI22_X1 U1147 ( .A1(\REGISTERS[22][5] ), .A2(n51), .B1(\REGISTERS[4][5] ), 
        .B2(n37), .ZN(n1036) );
  NAND4_X1 U1148 ( .A1(n1039), .A2(n1038), .A3(n1037), .A4(n1036), .ZN(n1045)
         );
  AOI22_X1 U1149 ( .A1(\REGISTERS[29][5] ), .A2(n68), .B1(\REGISTERS[7][5] ), 
        .B2(n43), .ZN(n1043) );
  AOI22_X1 U1150 ( .A1(\REGISTERS[1][5] ), .A2(n1576), .B1(\REGISTERS[2][5] ), 
        .B2(n46), .ZN(n1042) );
  AOI22_X1 U1151 ( .A1(\REGISTERS[23][5] ), .A2(n48), .B1(\REGISTERS[27][5] ), 
        .B2(n40), .ZN(n1041) );
  AOI22_X1 U1152 ( .A1(\REGISTERS[24][5] ), .A2(n47), .B1(\REGISTERS[9][5] ), 
        .B2(n42), .ZN(n1040) );
  NAND4_X1 U1153 ( .A1(n1043), .A2(n1042), .A3(n1041), .A4(n1040), .ZN(n1044)
         );
  NOR4_X1 U1154 ( .A1(n1047), .A2(n1046), .A3(n1045), .A4(n1044), .ZN(n1048)
         );
  AOI22_X1 U1155 ( .A1(n70), .A2(n126), .B1(n1048), .B2(n71), .ZN(N384) );
  AOI22_X1 U1156 ( .A1(\REGISTERS[21][6] ), .A2(n1598), .B1(\REGISTERS[28][6] ), .B2(n60), .ZN(n1052) );
  AOI22_X1 U1157 ( .A1(\REGISTERS[18][6] ), .A2(n59), .B1(\REGISTERS[22][6] ), 
        .B2(n51), .ZN(n1051) );
  AOI22_X1 U1158 ( .A1(\REGISTERS[11][6] ), .A2(n1590), .B1(\REGISTERS[9][6] ), 
        .B2(n42), .ZN(n1050) );
  AOI22_X1 U1159 ( .A1(\REGISTERS[16][6] ), .A2(n1612), .B1(\REGISTERS[20][6] ), .B2(n66), .ZN(n1049) );
  NAND4_X1 U1160 ( .A1(n1052), .A2(n1051), .A3(n1050), .A4(n1049), .ZN(n1068)
         );
  AOI22_X1 U1161 ( .A1(\REGISTERS[6][6] ), .A2(n1616), .B1(\REGISTERS[26][6] ), 
        .B2(n57), .ZN(n1056) );
  AOI22_X1 U1162 ( .A1(\REGISTERS[25][6] ), .A2(n61), .B1(\REGISTERS[10][6] ), 
        .B2(n41), .ZN(n1055) );
  AOI22_X1 U1163 ( .A1(\REGISTERS[5][6] ), .A2(n1611), .B1(\REGISTERS[30][6] ), 
        .B2(n65), .ZN(n1054) );
  AOI22_X1 U1164 ( .A1(\REGISTERS[3][6] ), .A2(n50), .B1(\REGISTERS[12][6] ), 
        .B2(n56), .ZN(n1053) );
  NAND4_X1 U1165 ( .A1(n1056), .A2(n1055), .A3(n1054), .A4(n1053), .ZN(n1067)
         );
  AOI22_X1 U1166 ( .A1(\REGISTERS[13][6] ), .A2(n1586), .B1(\REGISTERS[8][6] ), 
        .B2(n38), .ZN(n1060) );
  AOI22_X1 U1167 ( .A1(\REGISTERS[15][6] ), .A2(n1600), .B1(\REGISTERS[29][6] ), .B2(n68), .ZN(n1059) );
  AOI22_X1 U1168 ( .A1(\REGISTERS[27][6] ), .A2(n40), .B1(\REGISTERS[24][6] ), 
        .B2(n47), .ZN(n1058) );
  AOI22_X1 U1169 ( .A1(\REGISTERS[14][6] ), .A2(n44), .B1(\REGISTERS[2][6] ), 
        .B2(n46), .ZN(n1057) );
  NAND4_X1 U1170 ( .A1(n1060), .A2(n1059), .A3(n1058), .A4(n1057), .ZN(n1066)
         );
  AOI22_X1 U1171 ( .A1(\REGISTERS[31][6] ), .A2(n1599), .B1(\REGISTERS[1][6] ), 
        .B2(n39), .ZN(n1064) );
  AOI22_X1 U1172 ( .A1(\REGISTERS[7][6] ), .A2(n1580), .B1(\REGISTERS[4][6] ), 
        .B2(n37), .ZN(n1063) );
  AOI22_X1 U1173 ( .A1(\REGISTERS[19][6] ), .A2(n1603), .B1(\REGISTERS[17][6] ), .B2(n52), .ZN(n1062) );
  AOI22_X1 U1174 ( .A1(\REGISTERS[0][6] ), .A2(n64), .B1(\REGISTERS[23][6] ), 
        .B2(n48), .ZN(n1061) );
  NAND4_X1 U1175 ( .A1(n1064), .A2(n1063), .A3(n1062), .A4(n1061), .ZN(n1065)
         );
  NOR4_X1 U1176 ( .A1(n1068), .A2(n1067), .A3(n1066), .A4(n1065), .ZN(n1069)
         );
  AOI22_X1 U1177 ( .A1(n1627), .A2(n124), .B1(n1069), .B2(n71), .ZN(N385) );
  AOI22_X1 U1178 ( .A1(\REGISTERS[27][7] ), .A2(n40), .B1(\REGISTERS[1][7] ), 
        .B2(n39), .ZN(n1073) );
  AOI22_X1 U1179 ( .A1(\REGISTERS[29][7] ), .A2(n68), .B1(\REGISTERS[15][7] ), 
        .B2(n55), .ZN(n1072) );
  AOI22_X1 U1180 ( .A1(\REGISTERS[5][7] ), .A2(n62), .B1(\REGISTERS[30][7] ), 
        .B2(n65), .ZN(n1071) );
  AOI22_X1 U1181 ( .A1(\REGISTERS[28][7] ), .A2(n1605), .B1(\REGISTERS[17][7] ), .B2(n52), .ZN(n1070) );
  NAND4_X1 U1182 ( .A1(n1073), .A2(n1072), .A3(n1071), .A4(n1070), .ZN(n1089)
         );
  AOI22_X1 U1183 ( .A1(\REGISTERS[2][7] ), .A2(n1587), .B1(\REGISTERS[20][7] ), 
        .B2(n66), .ZN(n1077) );
  AOI22_X1 U1184 ( .A1(\REGISTERS[25][7] ), .A2(n1610), .B1(\REGISTERS[21][7] ), .B2(n53), .ZN(n1076) );
  AOI22_X1 U1185 ( .A1(\REGISTERS[12][7] ), .A2(n1601), .B1(\REGISTERS[26][7] ), .B2(n57), .ZN(n1075) );
  AOI22_X1 U1186 ( .A1(\REGISTERS[24][7] ), .A2(n1588), .B1(\REGISTERS[4][7] ), 
        .B2(n37), .ZN(n1074) );
  NAND4_X1 U1187 ( .A1(n1077), .A2(n1076), .A3(n1075), .A4(n1074), .ZN(n1088)
         );
  AOI22_X1 U1188 ( .A1(\REGISTERS[10][7] ), .A2(n1578), .B1(\REGISTERS[11][7] ), .B2(n49), .ZN(n1081) );
  AOI22_X1 U1189 ( .A1(\REGISTERS[16][7] ), .A2(n1612), .B1(\REGISTERS[18][7] ), .B2(n59), .ZN(n1080) );
  AOI22_X1 U1190 ( .A1(\REGISTERS[31][7] ), .A2(n1599), .B1(\REGISTERS[14][7] ), .B2(n44), .ZN(n1079) );
  AOI22_X1 U1191 ( .A1(\REGISTERS[9][7] ), .A2(n42), .B1(\REGISTERS[22][7] ), 
        .B2(n51), .ZN(n1078) );
  NAND4_X1 U1192 ( .A1(n1081), .A2(n1080), .A3(n1079), .A4(n1078), .ZN(n1087)
         );
  AOI22_X1 U1193 ( .A1(\REGISTERS[6][7] ), .A2(n67), .B1(\REGISTERS[13][7] ), 
        .B2(n45), .ZN(n1085) );
  AOI22_X1 U1194 ( .A1(\REGISTERS[7][7] ), .A2(n1580), .B1(\REGISTERS[3][7] ), 
        .B2(n50), .ZN(n1084) );
  AOI22_X1 U1195 ( .A1(\REGISTERS[19][7] ), .A2(n58), .B1(\REGISTERS[8][7] ), 
        .B2(n38), .ZN(n1083) );
  AOI22_X1 U1196 ( .A1(\REGISTERS[23][7] ), .A2(n1589), .B1(\REGISTERS[0][7] ), 
        .B2(n64), .ZN(n1082) );
  NAND4_X1 U1197 ( .A1(n1085), .A2(n1084), .A3(n1083), .A4(n1082), .ZN(n1086)
         );
  NOR4_X1 U1198 ( .A1(n1089), .A2(n1088), .A3(n1087), .A4(n1086), .ZN(n1090)
         );
  AOI22_X1 U1199 ( .A1(n1627), .A2(n122), .B1(n1090), .B2(n72), .ZN(N386) );
  AOI22_X1 U1200 ( .A1(\REGISTERS[30][8] ), .A2(n1614), .B1(\REGISTERS[24][8] ), .B2(n47), .ZN(n1094) );
  AOI22_X1 U1201 ( .A1(\REGISTERS[0][8] ), .A2(n1613), .B1(\REGISTERS[16][8] ), 
        .B2(n63), .ZN(n1093) );
  AOI22_X1 U1202 ( .A1(\REGISTERS[13][8] ), .A2(n1586), .B1(\REGISTERS[20][8] ), .B2(n66), .ZN(n1092) );
  AOI22_X1 U1203 ( .A1(\REGISTERS[14][8] ), .A2(n44), .B1(\REGISTERS[2][8] ), 
        .B2(n46), .ZN(n1091) );
  NAND4_X1 U1204 ( .A1(n1094), .A2(n1093), .A3(n1092), .A4(n1091), .ZN(n1110)
         );
  AOI22_X1 U1205 ( .A1(\REGISTERS[31][8] ), .A2(n54), .B1(\REGISTERS[15][8] ), 
        .B2(n55), .ZN(n1098) );
  AOI22_X1 U1206 ( .A1(\REGISTERS[27][8] ), .A2(n40), .B1(\REGISTERS[12][8] ), 
        .B2(n56), .ZN(n1097) );
  AOI22_X1 U1207 ( .A1(\REGISTERS[7][8] ), .A2(n1580), .B1(\REGISTERS[22][8] ), 
        .B2(n51), .ZN(n1096) );
  AOI22_X1 U1208 ( .A1(\REGISTERS[21][8] ), .A2(n1598), .B1(\REGISTERS[9][8] ), 
        .B2(n42), .ZN(n1095) );
  NAND4_X1 U1209 ( .A1(n1098), .A2(n1097), .A3(n1096), .A4(n1095), .ZN(n1109)
         );
  AOI22_X1 U1210 ( .A1(\REGISTERS[29][8] ), .A2(n1617), .B1(\REGISTERS[6][8] ), 
        .B2(n67), .ZN(n1102) );
  AOI22_X1 U1211 ( .A1(\REGISTERS[25][8] ), .A2(n1610), .B1(\REGISTERS[5][8] ), 
        .B2(n62), .ZN(n1101) );
  AOI22_X1 U1212 ( .A1(\REGISTERS[26][8] ), .A2(n57), .B1(\REGISTERS[17][8] ), 
        .B2(n52), .ZN(n1100) );
  AOI22_X1 U1213 ( .A1(\REGISTERS[8][8] ), .A2(n1575), .B1(\REGISTERS[11][8] ), 
        .B2(n49), .ZN(n1099) );
  NAND4_X1 U1214 ( .A1(n1102), .A2(n1101), .A3(n1100), .A4(n1099), .ZN(n1108)
         );
  AOI22_X1 U1215 ( .A1(\REGISTERS[19][8] ), .A2(n58), .B1(\REGISTERS[1][8] ), 
        .B2(n39), .ZN(n1106) );
  AOI22_X1 U1216 ( .A1(\REGISTERS[3][8] ), .A2(n50), .B1(\REGISTERS[18][8] ), 
        .B2(n59), .ZN(n1105) );
  AOI22_X1 U1217 ( .A1(\REGISTERS[28][8] ), .A2(n1605), .B1(\REGISTERS[10][8] ), .B2(n41), .ZN(n1104) );
  AOI22_X1 U1218 ( .A1(\REGISTERS[4][8] ), .A2(n1574), .B1(\REGISTERS[23][8] ), 
        .B2(n48), .ZN(n1103) );
  NAND4_X1 U1219 ( .A1(n1106), .A2(n1105), .A3(n1104), .A4(n1103), .ZN(n1107)
         );
  NOR4_X1 U1220 ( .A1(n1110), .A2(n1109), .A3(n1108), .A4(n1107), .ZN(n1111)
         );
  AOI22_X1 U1221 ( .A1(n1627), .A2(n120), .B1(n1111), .B2(n72), .ZN(N387) );
  AOI22_X1 U1222 ( .A1(\REGISTERS[15][9] ), .A2(n1600), .B1(\REGISTERS[26][9] ), .B2(n57), .ZN(n1115) );
  AOI22_X1 U1223 ( .A1(\REGISTERS[2][9] ), .A2(n1587), .B1(\REGISTERS[25][9] ), 
        .B2(n61), .ZN(n1114) );
  AOI22_X1 U1224 ( .A1(\REGISTERS[19][9] ), .A2(n58), .B1(\REGISTERS[24][9] ), 
        .B2(n47), .ZN(n1113) );
  AOI22_X1 U1225 ( .A1(\REGISTERS[3][9] ), .A2(n50), .B1(\REGISTERS[16][9] ), 
        .B2(n63), .ZN(n1112) );
  NAND4_X1 U1226 ( .A1(n1115), .A2(n1114), .A3(n1113), .A4(n1112), .ZN(n1131)
         );
  AOI22_X1 U1227 ( .A1(\REGISTERS[21][9] ), .A2(n1598), .B1(\REGISTERS[6][9] ), 
        .B2(n67), .ZN(n1119) );
  AOI22_X1 U1228 ( .A1(\REGISTERS[5][9] ), .A2(n1611), .B1(\REGISTERS[9][9] ), 
        .B2(n42), .ZN(n1118) );
  AOI22_X1 U1229 ( .A1(\REGISTERS[31][9] ), .A2(n54), .B1(\REGISTERS[11][9] ), 
        .B2(n49), .ZN(n1117) );
  AOI22_X1 U1230 ( .A1(\REGISTERS[27][9] ), .A2(n40), .B1(\REGISTERS[13][9] ), 
        .B2(n45), .ZN(n1116) );
  NAND4_X1 U1231 ( .A1(n1119), .A2(n1118), .A3(n1117), .A4(n1116), .ZN(n1130)
         );
  AOI22_X1 U1232 ( .A1(\REGISTERS[22][9] ), .A2(n1592), .B1(\REGISTERS[7][9] ), 
        .B2(n43), .ZN(n1123) );
  AOI22_X1 U1233 ( .A1(\REGISTERS[8][9] ), .A2(n1575), .B1(\REGISTERS[20][9] ), 
        .B2(n66), .ZN(n1122) );
  AOI22_X1 U1234 ( .A1(\REGISTERS[14][9] ), .A2(n44), .B1(\REGISTERS[1][9] ), 
        .B2(n39), .ZN(n1121) );
  AOI22_X1 U1235 ( .A1(\REGISTERS[17][9] ), .A2(n52), .B1(\REGISTERS[28][9] ), 
        .B2(n60), .ZN(n1120) );
  NAND4_X1 U1236 ( .A1(n1123), .A2(n1122), .A3(n1121), .A4(n1120), .ZN(n1129)
         );
  AOI22_X1 U1237 ( .A1(\REGISTERS[30][9] ), .A2(n1614), .B1(\REGISTERS[12][9] ), .B2(n56), .ZN(n1127) );
  AOI22_X1 U1238 ( .A1(\REGISTERS[29][9] ), .A2(n1617), .B1(\REGISTERS[4][9] ), 
        .B2(n37), .ZN(n1126) );
  AOI22_X1 U1239 ( .A1(\REGISTERS[10][9] ), .A2(n1578), .B1(\REGISTERS[0][9] ), 
        .B2(n64), .ZN(n1125) );
  AOI22_X1 U1240 ( .A1(\REGISTERS[18][9] ), .A2(n59), .B1(\REGISTERS[23][9] ), 
        .B2(n48), .ZN(n1124) );
  NAND4_X1 U1241 ( .A1(n1127), .A2(n1126), .A3(n1125), .A4(n1124), .ZN(n1128)
         );
  NOR4_X1 U1242 ( .A1(n1131), .A2(n1130), .A3(n1129), .A4(n1128), .ZN(n1132)
         );
  AOI22_X1 U1243 ( .A1(n1627), .A2(n118), .B1(n1132), .B2(n71), .ZN(N388) );
  AOI22_X1 U1244 ( .A1(\REGISTERS[3][10] ), .A2(n50), .B1(\REGISTERS[9][10] ), 
        .B2(n42), .ZN(n1136) );
  AOI22_X1 U1245 ( .A1(\REGISTERS[27][10] ), .A2(n1577), .B1(
        \REGISTERS[17][10] ), .B2(n52), .ZN(n1135) );
  AOI22_X1 U1246 ( .A1(\REGISTERS[2][10] ), .A2(n1587), .B1(
        \REGISTERS[18][10] ), .B2(n59), .ZN(n1134) );
  AOI22_X1 U1247 ( .A1(\REGISTERS[4][10] ), .A2(n1574), .B1(
        \REGISTERS[19][10] ), .B2(n58), .ZN(n1133) );
  NAND4_X1 U1248 ( .A1(n1136), .A2(n1135), .A3(n1134), .A4(n1133), .ZN(n1152)
         );
  AOI22_X1 U1249 ( .A1(\REGISTERS[23][10] ), .A2(n1589), .B1(
        \REGISTERS[8][10] ), .B2(n38), .ZN(n1140) );
  AOI22_X1 U1250 ( .A1(\REGISTERS[1][10] ), .A2(n1576), .B1(
        \REGISTERS[16][10] ), .B2(n63), .ZN(n1139) );
  AOI22_X1 U1251 ( .A1(\REGISTERS[24][10] ), .A2(n1588), .B1(
        \REGISTERS[26][10] ), .B2(n57), .ZN(n1138) );
  AOI22_X1 U1252 ( .A1(\REGISTERS[31][10] ), .A2(n54), .B1(\REGISTERS[11][10] ), .B2(n49), .ZN(n1137) );
  NAND4_X1 U1253 ( .A1(n1140), .A2(n1139), .A3(n1138), .A4(n1137), .ZN(n1151)
         );
  AOI22_X1 U1254 ( .A1(\REGISTERS[22][10] ), .A2(n1592), .B1(
        \REGISTERS[29][10] ), .B2(n68), .ZN(n1144) );
  AOI22_X1 U1255 ( .A1(\REGISTERS[15][10] ), .A2(n1600), .B1(
        \REGISTERS[0][10] ), .B2(n64), .ZN(n1143) );
  AOI22_X1 U1256 ( .A1(\REGISTERS[10][10] ), .A2(n1578), .B1(
        \REGISTERS[25][10] ), .B2(n61), .ZN(n1142) );
  AOI22_X1 U1257 ( .A1(\REGISTERS[14][10] ), .A2(n1581), .B1(
        \REGISTERS[6][10] ), .B2(n67), .ZN(n1141) );
  NAND4_X1 U1258 ( .A1(n1144), .A2(n1143), .A3(n1142), .A4(n1141), .ZN(n1150)
         );
  AOI22_X1 U1259 ( .A1(\REGISTERS[20][10] ), .A2(n66), .B1(\REGISTERS[7][10] ), 
        .B2(n43), .ZN(n1148) );
  AOI22_X1 U1260 ( .A1(\REGISTERS[12][10] ), .A2(n56), .B1(\REGISTERS[28][10] ), .B2(n60), .ZN(n1147) );
  AOI22_X1 U1261 ( .A1(\REGISTERS[21][10] ), .A2(n1598), .B1(
        \REGISTERS[30][10] ), .B2(n65), .ZN(n1146) );
  AOI22_X1 U1262 ( .A1(\REGISTERS[5][10] ), .A2(n1611), .B1(
        \REGISTERS[13][10] ), .B2(n45), .ZN(n1145) );
  NAND4_X1 U1263 ( .A1(n1148), .A2(n1147), .A3(n1146), .A4(n1145), .ZN(n1149)
         );
  NOR4_X1 U1264 ( .A1(n1152), .A2(n1151), .A3(n1150), .A4(n1149), .ZN(n1153)
         );
  AOI22_X1 U1265 ( .A1(n1627), .A2(n116), .B1(n1153), .B2(n72), .ZN(N389) );
  AOI22_X1 U1266 ( .A1(\REGISTERS[23][11] ), .A2(n1589), .B1(
        \REGISTERS[21][11] ), .B2(n53), .ZN(n1157) );
  AOI22_X1 U1267 ( .A1(\REGISTERS[10][11] ), .A2(n1578), .B1(
        \REGISTERS[6][11] ), .B2(n67), .ZN(n1156) );
  AOI22_X1 U1268 ( .A1(\REGISTERS[2][11] ), .A2(n1587), .B1(
        \REGISTERS[14][11] ), .B2(n44), .ZN(n1155) );
  AOI22_X1 U1269 ( .A1(\REGISTERS[9][11] ), .A2(n42), .B1(\REGISTERS[7][11] ), 
        .B2(n43), .ZN(n1154) );
  NAND4_X1 U1270 ( .A1(n1157), .A2(n1156), .A3(n1155), .A4(n1154), .ZN(n1173)
         );
  AOI22_X1 U1271 ( .A1(\REGISTERS[1][11] ), .A2(n1576), .B1(
        \REGISTERS[27][11] ), .B2(n40), .ZN(n1161) );
  AOI22_X1 U1272 ( .A1(\REGISTERS[13][11] ), .A2(n1586), .B1(
        \REGISTERS[11][11] ), .B2(n49), .ZN(n1160) );
  AOI22_X1 U1273 ( .A1(\REGISTERS[18][11] ), .A2(n1604), .B1(
        \REGISTERS[24][11] ), .B2(n47), .ZN(n1159) );
  AOI22_X1 U1274 ( .A1(\REGISTERS[3][11] ), .A2(n1591), .B1(
        \REGISTERS[20][11] ), .B2(n66), .ZN(n1158) );
  NAND4_X1 U1275 ( .A1(n1161), .A2(n1160), .A3(n1159), .A4(n1158), .ZN(n1172)
         );
  AOI22_X1 U1276 ( .A1(\REGISTERS[29][11] ), .A2(n1617), .B1(
        \REGISTERS[4][11] ), .B2(n37), .ZN(n1165) );
  AOI22_X1 U1277 ( .A1(\REGISTERS[25][11] ), .A2(n1610), .B1(
        \REGISTERS[30][11] ), .B2(n65), .ZN(n1164) );
  AOI22_X1 U1278 ( .A1(\REGISTERS[8][11] ), .A2(n1575), .B1(
        \REGISTERS[22][11] ), .B2(n51), .ZN(n1163) );
  AOI22_X1 U1279 ( .A1(\REGISTERS[19][11] ), .A2(n58), .B1(\REGISTERS[5][11] ), 
        .B2(n62), .ZN(n1162) );
  NAND4_X1 U1280 ( .A1(n1165), .A2(n1164), .A3(n1163), .A4(n1162), .ZN(n1171)
         );
  AOI22_X1 U1281 ( .A1(\REGISTERS[26][11] ), .A2(n1602), .B1(
        \REGISTERS[15][11] ), .B2(n55), .ZN(n1169) );
  AOI22_X1 U1282 ( .A1(\REGISTERS[31][11] ), .A2(n1599), .B1(
        \REGISTERS[0][11] ), .B2(n64), .ZN(n1168) );
  AOI22_X1 U1283 ( .A1(\REGISTERS[17][11] ), .A2(n52), .B1(\REGISTERS[28][11] ), .B2(n60), .ZN(n1167) );
  AOI22_X1 U1284 ( .A1(\REGISTERS[12][11] ), .A2(n56), .B1(\REGISTERS[16][11] ), .B2(n63), .ZN(n1166) );
  NAND4_X1 U1285 ( .A1(n1169), .A2(n1168), .A3(n1167), .A4(n1166), .ZN(n1170)
         );
  NOR4_X1 U1286 ( .A1(n1173), .A2(n1172), .A3(n1171), .A4(n1170), .ZN(n1174)
         );
  AOI22_X1 U1287 ( .A1(n1627), .A2(n114), .B1(n1174), .B2(n71), .ZN(N390) );
  AOI22_X1 U1288 ( .A1(\REGISTERS[25][12] ), .A2(n1610), .B1(
        \REGISTERS[8][12] ), .B2(n38), .ZN(n1178) );
  AOI22_X1 U1289 ( .A1(\REGISTERS[21][12] ), .A2(n1598), .B1(
        \REGISTERS[30][12] ), .B2(n65), .ZN(n1177) );
  AOI22_X1 U1290 ( .A1(\REGISTERS[26][12] ), .A2(n1602), .B1(
        \REGISTERS[18][12] ), .B2(n59), .ZN(n1176) );
  AOI22_X1 U1291 ( .A1(\REGISTERS[19][12] ), .A2(n58), .B1(\REGISTERS[22][12] ), .B2(n51), .ZN(n1175) );
  NAND4_X1 U1292 ( .A1(n1178), .A2(n1177), .A3(n1176), .A4(n1175), .ZN(n1194)
         );
  AOI22_X1 U1293 ( .A1(\REGISTERS[3][12] ), .A2(n1591), .B1(
        \REGISTERS[10][12] ), .B2(n41), .ZN(n1182) );
  AOI22_X1 U1294 ( .A1(\REGISTERS[11][12] ), .A2(n1590), .B1(
        \REGISTERS[5][12] ), .B2(n62), .ZN(n1181) );
  AOI22_X1 U1295 ( .A1(\REGISTERS[4][12] ), .A2(n1574), .B1(
        \REGISTERS[23][12] ), .B2(n48), .ZN(n1180) );
  AOI22_X1 U1296 ( .A1(\REGISTERS[20][12] ), .A2(n1615), .B1(
        \REGISTERS[0][12] ), .B2(n64), .ZN(n1179) );
  NAND4_X1 U1297 ( .A1(n1182), .A2(n1181), .A3(n1180), .A4(n1179), .ZN(n1193)
         );
  AOI22_X1 U1298 ( .A1(\REGISTERS[6][12] ), .A2(n1616), .B1(
        \REGISTERS[28][12] ), .B2(n60), .ZN(n1186) );
  AOI22_X1 U1299 ( .A1(\REGISTERS[9][12] ), .A2(n1579), .B1(
        \REGISTERS[15][12] ), .B2(n55), .ZN(n1185) );
  AOI22_X1 U1300 ( .A1(\REGISTERS[2][12] ), .A2(n1587), .B1(
        \REGISTERS[27][12] ), .B2(n40), .ZN(n1184) );
  AOI22_X1 U1301 ( .A1(\REGISTERS[31][12] ), .A2(n1599), .B1(
        \REGISTERS[1][12] ), .B2(n39), .ZN(n1183) );
  NAND4_X1 U1302 ( .A1(n1186), .A2(n1185), .A3(n1184), .A4(n1183), .ZN(n1192)
         );
  AOI22_X1 U1303 ( .A1(\REGISTERS[17][12] ), .A2(n52), .B1(\REGISTERS[13][12] ), .B2(n45), .ZN(n1190) );
  AOI22_X1 U1304 ( .A1(\REGISTERS[16][12] ), .A2(n1612), .B1(
        \REGISTERS[12][12] ), .B2(n56), .ZN(n1189) );
  AOI22_X1 U1305 ( .A1(\REGISTERS[14][12] ), .A2(n1581), .B1(
        \REGISTERS[7][12] ), .B2(n43), .ZN(n1188) );
  AOI22_X1 U1306 ( .A1(\REGISTERS[24][12] ), .A2(n1588), .B1(
        \REGISTERS[29][12] ), .B2(n68), .ZN(n1187) );
  NAND4_X1 U1307 ( .A1(n1190), .A2(n1189), .A3(n1188), .A4(n1187), .ZN(n1191)
         );
  NOR4_X1 U1308 ( .A1(n1194), .A2(n1193), .A3(n1192), .A4(n1191), .ZN(n1195)
         );
  AOI22_X1 U1309 ( .A1(n69), .A2(n112), .B1(n1195), .B2(n72), .ZN(N391) );
  AOI22_X1 U1310 ( .A1(\REGISTERS[31][13] ), .A2(n1599), .B1(
        \REGISTERS[27][13] ), .B2(n40), .ZN(n1199) );
  AOI22_X1 U1311 ( .A1(\REGISTERS[22][13] ), .A2(n1592), .B1(
        \REGISTERS[8][13] ), .B2(n38), .ZN(n1198) );
  AOI22_X1 U1312 ( .A1(\REGISTERS[14][13] ), .A2(n1581), .B1(
        \REGISTERS[21][13] ), .B2(n53), .ZN(n1197) );
  AOI22_X1 U1313 ( .A1(\REGISTERS[5][13] ), .A2(n1611), .B1(\REGISTERS[6][13] ), .B2(n1616), .ZN(n1196) );
  NAND4_X1 U1314 ( .A1(n1199), .A2(n1198), .A3(n1197), .A4(n1196), .ZN(n1215)
         );
  AOI22_X1 U1315 ( .A1(\REGISTERS[12][13] ), .A2(n56), .B1(\REGISTERS[4][13] ), 
        .B2(n37), .ZN(n1203) );
  AOI22_X1 U1316 ( .A1(\REGISTERS[13][13] ), .A2(n1586), .B1(
        \REGISTERS[30][13] ), .B2(n65), .ZN(n1202) );
  AOI22_X1 U1317 ( .A1(\REGISTERS[17][13] ), .A2(n1593), .B1(
        \REGISTERS[3][13] ), .B2(n50), .ZN(n1201) );
  AOI22_X1 U1318 ( .A1(\REGISTERS[11][13] ), .A2(n1590), .B1(
        \REGISTERS[20][13] ), .B2(n66), .ZN(n1200) );
  NAND4_X1 U1319 ( .A1(n1203), .A2(n1202), .A3(n1201), .A4(n1200), .ZN(n1214)
         );
  AOI22_X1 U1320 ( .A1(\REGISTERS[23][13] ), .A2(n1589), .B1(
        \REGISTERS[18][13] ), .B2(n59), .ZN(n1207) );
  AOI22_X1 U1321 ( .A1(\REGISTERS[0][13] ), .A2(n1613), .B1(
        \REGISTERS[29][13] ), .B2(n68), .ZN(n1206) );
  AOI22_X1 U1322 ( .A1(\REGISTERS[9][13] ), .A2(n1579), .B1(
        \REGISTERS[26][13] ), .B2(n57), .ZN(n1205) );
  AOI22_X1 U1323 ( .A1(\REGISTERS[28][13] ), .A2(n1605), .B1(
        \REGISTERS[7][13] ), .B2(n43), .ZN(n1204) );
  NAND4_X1 U1324 ( .A1(n1207), .A2(n1206), .A3(n1205), .A4(n1204), .ZN(n1213)
         );
  AOI22_X1 U1325 ( .A1(\REGISTERS[24][13] ), .A2(n1588), .B1(
        \REGISTERS[16][13] ), .B2(n63), .ZN(n1211) );
  AOI22_X1 U1326 ( .A1(\REGISTERS[19][13] ), .A2(n58), .B1(\REGISTERS[1][13] ), 
        .B2(n39), .ZN(n1210) );
  AOI22_X1 U1327 ( .A1(\REGISTERS[10][13] ), .A2(n1578), .B1(
        \REGISTERS[25][13] ), .B2(n61), .ZN(n1209) );
  AOI22_X1 U1328 ( .A1(\REGISTERS[2][13] ), .A2(n1587), .B1(
        \REGISTERS[15][13] ), .B2(n55), .ZN(n1208) );
  NAND4_X1 U1329 ( .A1(n1211), .A2(n1210), .A3(n1209), .A4(n1208), .ZN(n1212)
         );
  NOR4_X1 U1330 ( .A1(n1215), .A2(n1214), .A3(n1213), .A4(n1212), .ZN(n1216)
         );
  AOI22_X1 U1331 ( .A1(n69), .A2(n110), .B1(n1216), .B2(n71), .ZN(N392) );
  AOI22_X1 U1332 ( .A1(\REGISTERS[22][14] ), .A2(n1592), .B1(
        \REGISTERS[13][14] ), .B2(n45), .ZN(n1220) );
  AOI22_X1 U1333 ( .A1(\REGISTERS[7][14] ), .A2(n1580), .B1(\REGISTERS[5][14] ), .B2(n62), .ZN(n1219) );
  AOI22_X1 U1334 ( .A1(\REGISTERS[26][14] ), .A2(n1602), .B1(
        \REGISTERS[27][14] ), .B2(n40), .ZN(n1218) );
  AOI22_X1 U1335 ( .A1(\REGISTERS[20][14] ), .A2(n1615), .B1(
        \REGISTERS[25][14] ), .B2(n61), .ZN(n1217) );
  NAND4_X1 U1336 ( .A1(n1220), .A2(n1219), .A3(n1218), .A4(n1217), .ZN(n1236)
         );
  AOI22_X1 U1337 ( .A1(\REGISTERS[4][14] ), .A2(n1574), .B1(
        \REGISTERS[18][14] ), .B2(n59), .ZN(n1224) );
  AOI22_X1 U1338 ( .A1(\REGISTERS[12][14] ), .A2(n1601), .B1(
        \REGISTERS[1][14] ), .B2(n39), .ZN(n1223) );
  AOI22_X1 U1339 ( .A1(\REGISTERS[24][14] ), .A2(n47), .B1(\REGISTERS[14][14] ), .B2(n44), .ZN(n1222) );
  AOI22_X1 U1340 ( .A1(\REGISTERS[19][14] ), .A2(n58), .B1(\REGISTERS[9][14] ), 
        .B2(n42), .ZN(n1221) );
  NAND4_X1 U1341 ( .A1(n1224), .A2(n1223), .A3(n1222), .A4(n1221), .ZN(n1235)
         );
  AOI22_X1 U1342 ( .A1(\REGISTERS[17][14] ), .A2(n1593), .B1(
        \REGISTERS[11][14] ), .B2(n49), .ZN(n1228) );
  AOI22_X1 U1343 ( .A1(\REGISTERS[31][14] ), .A2(n1599), .B1(
        \REGISTERS[30][14] ), .B2(n65), .ZN(n1227) );
  AOI22_X1 U1344 ( .A1(\REGISTERS[28][14] ), .A2(n1605), .B1(
        \REGISTERS[10][14] ), .B2(n41), .ZN(n1226) );
  AOI22_X1 U1345 ( .A1(\REGISTERS[2][14] ), .A2(n1587), .B1(
        \REGISTERS[21][14] ), .B2(n53), .ZN(n1225) );
  NAND4_X1 U1346 ( .A1(n1228), .A2(n1227), .A3(n1226), .A4(n1225), .ZN(n1234)
         );
  AOI22_X1 U1347 ( .A1(\REGISTERS[29][14] ), .A2(n1617), .B1(
        \REGISTERS[23][14] ), .B2(n48), .ZN(n1232) );
  AOI22_X1 U1348 ( .A1(\REGISTERS[0][14] ), .A2(n1613), .B1(
        \REGISTERS[15][14] ), .B2(n55), .ZN(n1231) );
  AOI22_X1 U1349 ( .A1(\REGISTERS[16][14] ), .A2(n1612), .B1(
        \REGISTERS[6][14] ), .B2(n67), .ZN(n1230) );
  AOI22_X1 U1350 ( .A1(\REGISTERS[8][14] ), .A2(n1575), .B1(\REGISTERS[3][14] ), .B2(n50), .ZN(n1229) );
  NAND4_X1 U1351 ( .A1(n1232), .A2(n1231), .A3(n1230), .A4(n1229), .ZN(n1233)
         );
  NOR4_X1 U1352 ( .A1(n1236), .A2(n1235), .A3(n1234), .A4(n1233), .ZN(n1237)
         );
  AOI22_X1 U1353 ( .A1(n69), .A2(n108), .B1(n1237), .B2(n72), .ZN(N393) );
  AOI22_X1 U1354 ( .A1(\REGISTERS[16][15] ), .A2(n63), .B1(\REGISTERS[30][15] ), .B2(n1614), .ZN(n1241) );
  AOI22_X1 U1355 ( .A1(\REGISTERS[29][15] ), .A2(n1617), .B1(
        \REGISTERS[12][15] ), .B2(n56), .ZN(n1240) );
  AOI22_X1 U1356 ( .A1(\REGISTERS[24][15] ), .A2(n47), .B1(\REGISTERS[10][15] ), .B2(n41), .ZN(n1239) );
  AOI22_X1 U1357 ( .A1(\REGISTERS[18][15] ), .A2(n1604), .B1(
        \REGISTERS[14][15] ), .B2(n44), .ZN(n1238) );
  NAND4_X1 U1358 ( .A1(n1241), .A2(n1240), .A3(n1239), .A4(n1238), .ZN(n1257)
         );
  AOI22_X1 U1359 ( .A1(\REGISTERS[20][15] ), .A2(n66), .B1(\REGISTERS[26][15] ), .B2(n57), .ZN(n1245) );
  AOI22_X1 U1360 ( .A1(\REGISTERS[6][15] ), .A2(n1616), .B1(\REGISTERS[4][15] ), .B2(n37), .ZN(n1244) );
  AOI22_X1 U1361 ( .A1(\REGISTERS[7][15] ), .A2(n1580), .B1(\REGISTERS[8][15] ), .B2(n38), .ZN(n1243) );
  AOI22_X1 U1362 ( .A1(\REGISTERS[19][15] ), .A2(n58), .B1(\REGISTERS[2][15] ), 
        .B2(n46), .ZN(n1242) );
  NAND4_X1 U1363 ( .A1(n1245), .A2(n1244), .A3(n1243), .A4(n1242), .ZN(n1256)
         );
  AOI22_X1 U1364 ( .A1(\REGISTERS[17][15] ), .A2(n1593), .B1(
        \REGISTERS[23][15] ), .B2(n48), .ZN(n1249) );
  AOI22_X1 U1365 ( .A1(\REGISTERS[27][15] ), .A2(n1577), .B1(
        \REGISTERS[28][15] ), .B2(n60), .ZN(n1248) );
  AOI22_X1 U1366 ( .A1(\REGISTERS[25][15] ), .A2(n1610), .B1(
        \REGISTERS[15][15] ), .B2(n1600), .ZN(n1247) );
  AOI22_X1 U1367 ( .A1(\REGISTERS[3][15] ), .A2(n1591), .B1(\REGISTERS[9][15] ), .B2(n42), .ZN(n1246) );
  NAND4_X1 U1368 ( .A1(n1249), .A2(n1248), .A3(n1247), .A4(n1246), .ZN(n1255)
         );
  AOI22_X1 U1369 ( .A1(\REGISTERS[22][15] ), .A2(n51), .B1(\REGISTERS[5][15] ), 
        .B2(n62), .ZN(n1253) );
  AOI22_X1 U1370 ( .A1(\REGISTERS[0][15] ), .A2(n1613), .B1(\REGISTERS[1][15] ), .B2(n39), .ZN(n1252) );
  AOI22_X1 U1371 ( .A1(\REGISTERS[31][15] ), .A2(n1599), .B1(
        \REGISTERS[11][15] ), .B2(n1590), .ZN(n1251) );
  AOI22_X1 U1372 ( .A1(\REGISTERS[13][15] ), .A2(n1586), .B1(
        \REGISTERS[21][15] ), .B2(n53), .ZN(n1250) );
  NAND4_X1 U1373 ( .A1(n1253), .A2(n1252), .A3(n1251), .A4(n1250), .ZN(n1254)
         );
  NOR4_X1 U1374 ( .A1(n1257), .A2(n1256), .A3(n1255), .A4(n1254), .ZN(n1258)
         );
  AOI22_X1 U1375 ( .A1(n69), .A2(n106), .B1(n1258), .B2(n71), .ZN(N394) );
  AOI22_X1 U1376 ( .A1(\REGISTERS[11][16] ), .A2(n1590), .B1(
        \REGISTERS[3][16] ), .B2(n50), .ZN(n1262) );
  AOI22_X1 U1377 ( .A1(\REGISTERS[12][16] ), .A2(n1601), .B1(
        \REGISTERS[20][16] ), .B2(n66), .ZN(n1261) );
  AOI22_X1 U1378 ( .A1(\REGISTERS[29][16] ), .A2(n1617), .B1(
        \REGISTERS[23][16] ), .B2(n48), .ZN(n1260) );
  AOI22_X1 U1379 ( .A1(\REGISTERS[6][16] ), .A2(n1616), .B1(\REGISTERS[0][16] ), .B2(n64), .ZN(n1259) );
  NAND4_X1 U1380 ( .A1(n1262), .A2(n1261), .A3(n1260), .A4(n1259), .ZN(n1278)
         );
  AOI22_X1 U1381 ( .A1(\REGISTERS[17][16] ), .A2(n1593), .B1(
        \REGISTERS[2][16] ), .B2(n46), .ZN(n1266) );
  AOI22_X1 U1382 ( .A1(\REGISTERS[18][16] ), .A2(n1604), .B1(
        \REGISTERS[24][16] ), .B2(n47), .ZN(n1265) );
  AOI22_X1 U1383 ( .A1(\REGISTERS[22][16] ), .A2(n51), .B1(\REGISTERS[5][16] ), 
        .B2(n62), .ZN(n1264) );
  AOI22_X1 U1384 ( .A1(\REGISTERS[4][16] ), .A2(n1574), .B1(
        \REGISTERS[28][16] ), .B2(n60), .ZN(n1263) );
  NAND4_X1 U1385 ( .A1(n1266), .A2(n1265), .A3(n1264), .A4(n1263), .ZN(n1277)
         );
  AOI22_X1 U1386 ( .A1(\REGISTERS[27][16] ), .A2(n1577), .B1(
        \REGISTERS[26][16] ), .B2(n57), .ZN(n1270) );
  AOI22_X1 U1387 ( .A1(\REGISTERS[9][16] ), .A2(n1579), .B1(
        \REGISTERS[14][16] ), .B2(n44), .ZN(n1269) );
  AOI22_X1 U1388 ( .A1(\REGISTERS[16][16] ), .A2(n1612), .B1(
        \REGISTERS[1][16] ), .B2(n39), .ZN(n1268) );
  AOI22_X1 U1389 ( .A1(\REGISTERS[19][16] ), .A2(n58), .B1(\REGISTERS[30][16] ), .B2(n1614), .ZN(n1267) );
  NAND4_X1 U1390 ( .A1(n1270), .A2(n1269), .A3(n1268), .A4(n1267), .ZN(n1276)
         );
  AOI22_X1 U1391 ( .A1(\REGISTERS[25][16] ), .A2(n1610), .B1(
        \REGISTERS[15][16] ), .B2(n1600), .ZN(n1274) );
  AOI22_X1 U1392 ( .A1(\REGISTERS[7][16] ), .A2(n1580), .B1(
        \REGISTERS[31][16] ), .B2(n54), .ZN(n1273) );
  AOI22_X1 U1393 ( .A1(\REGISTERS[13][16] ), .A2(n1586), .B1(
        \REGISTERS[21][16] ), .B2(n53), .ZN(n1272) );
  AOI22_X1 U1394 ( .A1(\REGISTERS[10][16] ), .A2(n41), .B1(\REGISTERS[8][16] ), 
        .B2(n38), .ZN(n1271) );
  NAND4_X1 U1395 ( .A1(n1274), .A2(n1273), .A3(n1272), .A4(n1271), .ZN(n1275)
         );
  NOR4_X1 U1396 ( .A1(n1278), .A2(n1277), .A3(n1276), .A4(n1275), .ZN(n1279)
         );
  AOI22_X1 U1397 ( .A1(n69), .A2(n104), .B1(n1279), .B2(n72), .ZN(N395) );
  AOI22_X1 U1398 ( .A1(\REGISTERS[24][17] ), .A2(n1588), .B1(
        \REGISTERS[0][17] ), .B2(n64), .ZN(n1283) );
  AOI22_X1 U1399 ( .A1(\REGISTERS[6][17] ), .A2(n1616), .B1(
        \REGISTERS[29][17] ), .B2(n68), .ZN(n1282) );
  AOI22_X1 U1400 ( .A1(\REGISTERS[5][17] ), .A2(n1611), .B1(
        \REGISTERS[21][17] ), .B2(n53), .ZN(n1281) );
  AOI22_X1 U1401 ( .A1(\REGISTERS[28][17] ), .A2(n1605), .B1(
        \REGISTERS[1][17] ), .B2(n39), .ZN(n1280) );
  NAND4_X1 U1402 ( .A1(n1283), .A2(n1282), .A3(n1281), .A4(n1280), .ZN(n1299)
         );
  AOI22_X1 U1403 ( .A1(\REGISTERS[14][17] ), .A2(n1581), .B1(
        \REGISTERS[16][17] ), .B2(n63), .ZN(n1287) );
  AOI22_X1 U1404 ( .A1(\REGISTERS[27][17] ), .A2(n1577), .B1(
        \REGISTERS[25][17] ), .B2(n61), .ZN(n1286) );
  AOI22_X1 U1405 ( .A1(\REGISTERS[3][17] ), .A2(n1591), .B1(
        \REGISTERS[10][17] ), .B2(n41), .ZN(n1285) );
  AOI22_X1 U1406 ( .A1(\REGISTERS[19][17] ), .A2(n1603), .B1(
        \REGISTERS[8][17] ), .B2(n38), .ZN(n1284) );
  NAND4_X1 U1407 ( .A1(n1287), .A2(n1286), .A3(n1285), .A4(n1284), .ZN(n1298)
         );
  AOI22_X1 U1408 ( .A1(\REGISTERS[17][17] ), .A2(n1593), .B1(
        \REGISTERS[9][17] ), .B2(n42), .ZN(n1291) );
  AOI22_X1 U1409 ( .A1(\REGISTERS[2][17] ), .A2(n1587), .B1(
        \REGISTERS[23][17] ), .B2(n48), .ZN(n1290) );
  AOI22_X1 U1410 ( .A1(\REGISTERS[18][17] ), .A2(n1604), .B1(
        \REGISTERS[7][17] ), .B2(n43), .ZN(n1289) );
  AOI22_X1 U1411 ( .A1(\REGISTERS[15][17] ), .A2(n1600), .B1(
        \REGISTERS[13][17] ), .B2(n45), .ZN(n1288) );
  NAND4_X1 U1412 ( .A1(n1291), .A2(n1290), .A3(n1289), .A4(n1288), .ZN(n1297)
         );
  AOI22_X1 U1413 ( .A1(\REGISTERS[26][17] ), .A2(n1602), .B1(
        \REGISTERS[11][17] ), .B2(n49), .ZN(n1295) );
  AOI22_X1 U1414 ( .A1(\REGISTERS[22][17] ), .A2(n51), .B1(\REGISTERS[4][17] ), 
        .B2(n37), .ZN(n1294) );
  AOI22_X1 U1415 ( .A1(\REGISTERS[20][17] ), .A2(n1615), .B1(
        \REGISTERS[12][17] ), .B2(n56), .ZN(n1293) );
  AOI22_X1 U1416 ( .A1(\REGISTERS[31][17] ), .A2(n1599), .B1(
        \REGISTERS[30][17] ), .B2(n65), .ZN(n1292) );
  NAND4_X1 U1417 ( .A1(n1295), .A2(n1294), .A3(n1293), .A4(n1292), .ZN(n1296)
         );
  NOR4_X1 U1418 ( .A1(n1299), .A2(n1298), .A3(n1297), .A4(n1296), .ZN(n1300)
         );
  AOI22_X1 U1419 ( .A1(n69), .A2(n102), .B1(n1300), .B2(n71), .ZN(N396) );
  AOI22_X1 U1420 ( .A1(\REGISTERS[30][18] ), .A2(n1614), .B1(
        \REGISTERS[20][18] ), .B2(n66), .ZN(n1304) );
  AOI22_X1 U1421 ( .A1(\REGISTERS[21][18] ), .A2(n1598), .B1(
        \REGISTERS[4][18] ), .B2(n1574), .ZN(n1303) );
  AOI22_X1 U1422 ( .A1(\REGISTERS[17][18] ), .A2(n1593), .B1(
        \REGISTERS[18][18] ), .B2(n59), .ZN(n1302) );
  AOI22_X1 U1423 ( .A1(\REGISTERS[11][18] ), .A2(n1590), .B1(
        \REGISTERS[3][18] ), .B2(n50), .ZN(n1301) );
  NAND4_X1 U1424 ( .A1(n1304), .A2(n1303), .A3(n1302), .A4(n1301), .ZN(n1320)
         );
  AOI22_X1 U1425 ( .A1(\REGISTERS[14][18] ), .A2(n1581), .B1(
        \REGISTERS[16][18] ), .B2(n63), .ZN(n1308) );
  AOI22_X1 U1426 ( .A1(\REGISTERS[12][18] ), .A2(n1601), .B1(
        \REGISTERS[15][18] ), .B2(n55), .ZN(n1307) );
  AOI22_X1 U1427 ( .A1(\REGISTERS[24][18] ), .A2(n1588), .B1(
        \REGISTERS[25][18] ), .B2(n61), .ZN(n1306) );
  AOI22_X1 U1428 ( .A1(\REGISTERS[22][18] ), .A2(n51), .B1(\REGISTERS[23][18] ), .B2(n48), .ZN(n1305) );
  NAND4_X1 U1429 ( .A1(n1308), .A2(n1307), .A3(n1306), .A4(n1305), .ZN(n1319)
         );
  AOI22_X1 U1430 ( .A1(\REGISTERS[9][18] ), .A2(n1579), .B1(\REGISTERS[7][18] ), .B2(n43), .ZN(n1312) );
  AOI22_X1 U1431 ( .A1(\REGISTERS[0][18] ), .A2(n1613), .B1(
        \REGISTERS[27][18] ), .B2(n40), .ZN(n1311) );
  AOI22_X1 U1432 ( .A1(\REGISTERS[13][18] ), .A2(n1586), .B1(
        \REGISTERS[31][18] ), .B2(n54), .ZN(n1310) );
  AOI22_X1 U1433 ( .A1(\REGISTERS[28][18] ), .A2(n1605), .B1(
        \REGISTERS[2][18] ), .B2(n46), .ZN(n1309) );
  NAND4_X1 U1434 ( .A1(n1312), .A2(n1311), .A3(n1310), .A4(n1309), .ZN(n1318)
         );
  AOI22_X1 U1435 ( .A1(\REGISTERS[19][18] ), .A2(n1603), .B1(
        \REGISTERS[26][18] ), .B2(n57), .ZN(n1316) );
  AOI22_X1 U1436 ( .A1(\REGISTERS[29][18] ), .A2(n68), .B1(\REGISTERS[8][18] ), 
        .B2(n38), .ZN(n1315) );
  AOI22_X1 U1437 ( .A1(\REGISTERS[6][18] ), .A2(n1616), .B1(\REGISTERS[5][18] ), .B2(n62), .ZN(n1314) );
  AOI22_X1 U1438 ( .A1(\REGISTERS[10][18] ), .A2(n1578), .B1(
        \REGISTERS[1][18] ), .B2(n39), .ZN(n1313) );
  NAND4_X1 U1439 ( .A1(n1316), .A2(n1315), .A3(n1314), .A4(n1313), .ZN(n1317)
         );
  NOR4_X1 U1440 ( .A1(n1320), .A2(n1319), .A3(n1318), .A4(n1317), .ZN(n1321)
         );
  AOI22_X1 U1441 ( .A1(n69), .A2(n100), .B1(n1321), .B2(n72), .ZN(N397) );
  AOI22_X1 U1442 ( .A1(\REGISTERS[25][19] ), .A2(n61), .B1(\REGISTERS[10][19] ), .B2(n41), .ZN(n1325) );
  AOI22_X1 U1443 ( .A1(\REGISTERS[8][19] ), .A2(n1575), .B1(
        \REGISTERS[29][19] ), .B2(n68), .ZN(n1324) );
  AOI22_X1 U1444 ( .A1(\REGISTERS[20][19] ), .A2(n1615), .B1(
        \REGISTERS[2][19] ), .B2(n46), .ZN(n1323) );
  AOI22_X1 U1445 ( .A1(\REGISTERS[19][19] ), .A2(n1603), .B1(
        \REGISTERS[17][19] ), .B2(n52), .ZN(n1322) );
  NAND4_X1 U1446 ( .A1(n1325), .A2(n1324), .A3(n1323), .A4(n1322), .ZN(n1341)
         );
  AOI22_X1 U1447 ( .A1(\REGISTERS[9][19] ), .A2(n1579), .B1(\REGISTERS[0][19] ), .B2(n64), .ZN(n1329) );
  AOI22_X1 U1448 ( .A1(\REGISTERS[5][19] ), .A2(n1611), .B1(
        \REGISTERS[28][19] ), .B2(n60), .ZN(n1328) );
  AOI22_X1 U1449 ( .A1(\REGISTERS[21][19] ), .A2(n53), .B1(\REGISTERS[6][19] ), 
        .B2(n67), .ZN(n1327) );
  AOI22_X1 U1450 ( .A1(\REGISTERS[12][19] ), .A2(n56), .B1(\REGISTERS[16][19] ), .B2(n63), .ZN(n1326) );
  NAND4_X1 U1451 ( .A1(n1329), .A2(n1328), .A3(n1327), .A4(n1326), .ZN(n1340)
         );
  AOI22_X1 U1452 ( .A1(\REGISTERS[7][19] ), .A2(n43), .B1(\REGISTERS[24][19] ), 
        .B2(n47), .ZN(n1333) );
  AOI22_X1 U1453 ( .A1(\REGISTERS[14][19] ), .A2(n44), .B1(\REGISTERS[15][19] ), .B2(n55), .ZN(n1332) );
  AOI22_X1 U1454 ( .A1(\REGISTERS[18][19] ), .A2(n1604), .B1(
        \REGISTERS[3][19] ), .B2(n50), .ZN(n1331) );
  AOI22_X1 U1455 ( .A1(\REGISTERS[1][19] ), .A2(n1576), .B1(
        \REGISTERS[13][19] ), .B2(n45), .ZN(n1330) );
  NAND4_X1 U1456 ( .A1(n1333), .A2(n1332), .A3(n1331), .A4(n1330), .ZN(n1339)
         );
  AOI22_X1 U1457 ( .A1(\REGISTERS[30][19] ), .A2(n1614), .B1(
        \REGISTERS[4][19] ), .B2(n1574), .ZN(n1337) );
  AOI22_X1 U1458 ( .A1(\REGISTERS[22][19] ), .A2(n51), .B1(\REGISTERS[23][19] ), .B2(n48), .ZN(n1336) );
  AOI22_X1 U1459 ( .A1(\REGISTERS[11][19] ), .A2(n1590), .B1(
        \REGISTERS[31][19] ), .B2(n54), .ZN(n1335) );
  AOI22_X1 U1460 ( .A1(\REGISTERS[27][19] ), .A2(n1577), .B1(
        \REGISTERS[26][19] ), .B2(n57), .ZN(n1334) );
  NAND4_X1 U1461 ( .A1(n1337), .A2(n1336), .A3(n1335), .A4(n1334), .ZN(n1338)
         );
  NOR4_X1 U1462 ( .A1(n1341), .A2(n1340), .A3(n1339), .A4(n1338), .ZN(n1342)
         );
  AOI22_X1 U1463 ( .A1(n69), .A2(n98), .B1(n1342), .B2(n72), .ZN(N398) );
  AOI22_X1 U1464 ( .A1(\REGISTERS[29][20] ), .A2(n1617), .B1(
        \REGISTERS[3][20] ), .B2(n50), .ZN(n1346) );
  AOI22_X1 U1465 ( .A1(\REGISTERS[20][20] ), .A2(n1615), .B1(
        \REGISTERS[31][20] ), .B2(n54), .ZN(n1345) );
  AOI22_X1 U1466 ( .A1(\REGISTERS[6][20] ), .A2(n1616), .B1(\REGISTERS[4][20] ), .B2(n37), .ZN(n1344) );
  AOI22_X1 U1467 ( .A1(\REGISTERS[2][20] ), .A2(n1587), .B1(
        \REGISTERS[16][20] ), .B2(n63), .ZN(n1343) );
  NAND4_X1 U1468 ( .A1(n1346), .A2(n1345), .A3(n1344), .A4(n1343), .ZN(n1362)
         );
  AOI22_X1 U1469 ( .A1(\REGISTERS[21][20] ), .A2(n1598), .B1(
        \REGISTERS[28][20] ), .B2(n60), .ZN(n1350) );
  AOI22_X1 U1470 ( .A1(\REGISTERS[10][20] ), .A2(n1578), .B1(
        \REGISTERS[8][20] ), .B2(n38), .ZN(n1349) );
  AOI22_X1 U1471 ( .A1(\REGISTERS[23][20] ), .A2(n1589), .B1(
        \REGISTERS[13][20] ), .B2(n45), .ZN(n1348) );
  AOI22_X1 U1472 ( .A1(\REGISTERS[26][20] ), .A2(n1602), .B1(
        \REGISTERS[25][20] ), .B2(n61), .ZN(n1347) );
  NAND4_X1 U1473 ( .A1(n1350), .A2(n1349), .A3(n1348), .A4(n1347), .ZN(n1361)
         );
  AOI22_X1 U1474 ( .A1(\REGISTERS[27][20] ), .A2(n1577), .B1(
        \REGISTERS[7][20] ), .B2(n43), .ZN(n1354) );
  AOI22_X1 U1475 ( .A1(\REGISTERS[19][20] ), .A2(n1603), .B1(
        \REGISTERS[9][20] ), .B2(n42), .ZN(n1353) );
  AOI22_X1 U1476 ( .A1(\REGISTERS[18][20] ), .A2(n1604), .B1(
        \REGISTERS[24][20] ), .B2(n47), .ZN(n1352) );
  AOI22_X1 U1477 ( .A1(\REGISTERS[30][20] ), .A2(n1614), .B1(
        \REGISTERS[12][20] ), .B2(n56), .ZN(n1351) );
  NAND4_X1 U1478 ( .A1(n1354), .A2(n1353), .A3(n1352), .A4(n1351), .ZN(n1360)
         );
  AOI22_X1 U1479 ( .A1(\REGISTERS[11][20] ), .A2(n1590), .B1(
        \REGISTERS[15][20] ), .B2(n55), .ZN(n1358) );
  AOI22_X1 U1480 ( .A1(\REGISTERS[17][20] ), .A2(n1593), .B1(
        \REGISTERS[5][20] ), .B2(n62), .ZN(n1357) );
  AOI22_X1 U1481 ( .A1(\REGISTERS[1][20] ), .A2(n1576), .B1(
        \REGISTERS[14][20] ), .B2(n44), .ZN(n1356) );
  AOI22_X1 U1482 ( .A1(\REGISTERS[22][20] ), .A2(n51), .B1(\REGISTERS[0][20] ), 
        .B2(n64), .ZN(n1355) );
  NAND4_X1 U1483 ( .A1(n1358), .A2(n1357), .A3(n1356), .A4(n1355), .ZN(n1359)
         );
  NOR4_X1 U1484 ( .A1(n1362), .A2(n1361), .A3(n1360), .A4(n1359), .ZN(n1363)
         );
  AOI22_X1 U1485 ( .A1(n69), .A2(n96), .B1(n1363), .B2(n71), .ZN(N399) );
  AOI22_X1 U1486 ( .A1(\REGISTERS[12][21] ), .A2(n1601), .B1(
        \REGISTERS[26][21] ), .B2(n57), .ZN(n1367) );
  AOI22_X1 U1487 ( .A1(\REGISTERS[22][21] ), .A2(n1592), .B1(
        \REGISTERS[20][21] ), .B2(n66), .ZN(n1366) );
  AOI22_X1 U1488 ( .A1(\REGISTERS[5][21] ), .A2(n1611), .B1(
        \REGISTERS[16][21] ), .B2(n63), .ZN(n1365) );
  AOI22_X1 U1489 ( .A1(\REGISTERS[28][21] ), .A2(n60), .B1(\REGISTERS[27][21] ), .B2(n40), .ZN(n1364) );
  NAND4_X1 U1490 ( .A1(n1367), .A2(n1366), .A3(n1365), .A4(n1364), .ZN(n1383)
         );
  AOI22_X1 U1491 ( .A1(\REGISTERS[0][21] ), .A2(n1613), .B1(\REGISTERS[6][21] ), .B2(n67), .ZN(n1371) );
  AOI22_X1 U1492 ( .A1(\REGISTERS[9][21] ), .A2(n1579), .B1(\REGISTERS[8][21] ), .B2(n1575), .ZN(n1370) );
  AOI22_X1 U1493 ( .A1(\REGISTERS[3][21] ), .A2(n1591), .B1(
        \REGISTERS[30][21] ), .B2(n65), .ZN(n1369) );
  AOI22_X1 U1494 ( .A1(\REGISTERS[2][21] ), .A2(n46), .B1(\REGISTERS[24][21] ), 
        .B2(n47), .ZN(n1368) );
  NAND4_X1 U1495 ( .A1(n1371), .A2(n1370), .A3(n1369), .A4(n1368), .ZN(n1382)
         );
  AOI22_X1 U1496 ( .A1(\REGISTERS[29][21] ), .A2(n68), .B1(\REGISTERS[15][21] ), .B2(n55), .ZN(n1375) );
  AOI22_X1 U1497 ( .A1(\REGISTERS[19][21] ), .A2(n1603), .B1(
        \REGISTERS[11][21] ), .B2(n49), .ZN(n1374) );
  AOI22_X1 U1498 ( .A1(\REGISTERS[1][21] ), .A2(n1576), .B1(
        \REGISTERS[13][21] ), .B2(n45), .ZN(n1373) );
  AOI22_X1 U1499 ( .A1(\REGISTERS[10][21] ), .A2(n1578), .B1(
        \REGISTERS[18][21] ), .B2(n59), .ZN(n1372) );
  NAND4_X1 U1500 ( .A1(n1375), .A2(n1374), .A3(n1373), .A4(n1372), .ZN(n1381)
         );
  AOI22_X1 U1501 ( .A1(\REGISTERS[21][21] ), .A2(n1598), .B1(
        \REGISTERS[4][21] ), .B2(n37), .ZN(n1379) );
  AOI22_X1 U1502 ( .A1(\REGISTERS[14][21] ), .A2(n1581), .B1(
        \REGISTERS[17][21] ), .B2(n52), .ZN(n1378) );
  AOI22_X1 U1503 ( .A1(\REGISTERS[7][21] ), .A2(n1580), .B1(
        \REGISTERS[25][21] ), .B2(n61), .ZN(n1377) );
  AOI22_X1 U1504 ( .A1(\REGISTERS[31][21] ), .A2(n54), .B1(\REGISTERS[23][21] ), .B2(n48), .ZN(n1376) );
  NAND4_X1 U1505 ( .A1(n1379), .A2(n1378), .A3(n1377), .A4(n1376), .ZN(n1380)
         );
  NOR4_X1 U1506 ( .A1(n1383), .A2(n1382), .A3(n1381), .A4(n1380), .ZN(n1384)
         );
  AOI22_X1 U1507 ( .A1(n69), .A2(n1781), .B1(n1384), .B2(n72), .ZN(N400) );
  AOI22_X1 U1508 ( .A1(\REGISTERS[13][22] ), .A2(n45), .B1(\REGISTERS[22][22] ), .B2(n51), .ZN(n1388) );
  AOI22_X1 U1509 ( .A1(\REGISTERS[9][22] ), .A2(n42), .B1(\REGISTERS[1][22] ), 
        .B2(n39), .ZN(n1387) );
  AOI22_X1 U1510 ( .A1(\REGISTERS[31][22] ), .A2(n1599), .B1(
        \REGISTERS[4][22] ), .B2(n37), .ZN(n1386) );
  AOI22_X1 U1511 ( .A1(\REGISTERS[27][22] ), .A2(n40), .B1(\REGISTERS[20][22] ), .B2(n66), .ZN(n1385) );
  NAND4_X1 U1512 ( .A1(n1388), .A2(n1387), .A3(n1386), .A4(n1385), .ZN(n1404)
         );
  AOI22_X1 U1513 ( .A1(\REGISTERS[23][22] ), .A2(n1589), .B1(
        \REGISTERS[25][22] ), .B2(n61), .ZN(n1392) );
  AOI22_X1 U1514 ( .A1(\REGISTERS[21][22] ), .A2(n53), .B1(\REGISTERS[11][22] ), .B2(n49), .ZN(n1391) );
  AOI22_X1 U1515 ( .A1(\REGISTERS[3][22] ), .A2(n1591), .B1(
        \REGISTERS[28][22] ), .B2(n60), .ZN(n1390) );
  AOI22_X1 U1516 ( .A1(\REGISTERS[12][22] ), .A2(n1601), .B1(
        \REGISTERS[29][22] ), .B2(n68), .ZN(n1389) );
  NAND4_X1 U1517 ( .A1(n1392), .A2(n1391), .A3(n1390), .A4(n1389), .ZN(n1403)
         );
  AOI22_X1 U1518 ( .A1(\REGISTERS[24][22] ), .A2(n1588), .B1(
        \REGISTERS[14][22] ), .B2(n44), .ZN(n1396) );
  AOI22_X1 U1519 ( .A1(\REGISTERS[18][22] ), .A2(n59), .B1(\REGISTERS[8][22] ), 
        .B2(n1575), .ZN(n1395) );
  AOI22_X1 U1520 ( .A1(\REGISTERS[6][22] ), .A2(n1616), .B1(
        \REGISTERS[19][22] ), .B2(n58), .ZN(n1394) );
  AOI22_X1 U1521 ( .A1(\REGISTERS[5][22] ), .A2(n62), .B1(\REGISTERS[16][22] ), 
        .B2(n63), .ZN(n1393) );
  NAND4_X1 U1522 ( .A1(n1396), .A2(n1395), .A3(n1394), .A4(n1393), .ZN(n1402)
         );
  AOI22_X1 U1523 ( .A1(\REGISTERS[2][22] ), .A2(n1587), .B1(
        \REGISTERS[15][22] ), .B2(n55), .ZN(n1400) );
  AOI22_X1 U1524 ( .A1(\REGISTERS[10][22] ), .A2(n41), .B1(\REGISTERS[30][22] ), .B2(n65), .ZN(n1399) );
  AOI22_X1 U1525 ( .A1(\REGISTERS[7][22] ), .A2(n43), .B1(\REGISTERS[17][22] ), 
        .B2(n52), .ZN(n1398) );
  AOI22_X1 U1526 ( .A1(\REGISTERS[26][22] ), .A2(n1602), .B1(
        \REGISTERS[0][22] ), .B2(n64), .ZN(n1397) );
  NAND4_X1 U1527 ( .A1(n1400), .A2(n1399), .A3(n1398), .A4(n1397), .ZN(n1401)
         );
  NOR4_X1 U1528 ( .A1(n1404), .A2(n1403), .A3(n1402), .A4(n1401), .ZN(n1405)
         );
  AOI22_X1 U1529 ( .A1(n69), .A2(n92), .B1(n1405), .B2(n72), .ZN(N401) );
  AOI22_X1 U1530 ( .A1(\REGISTERS[14][23] ), .A2(n44), .B1(\REGISTERS[4][23] ), 
        .B2(n37), .ZN(n1409) );
  AOI22_X1 U1531 ( .A1(\REGISTERS[2][23] ), .A2(n46), .B1(\REGISTERS[10][23] ), 
        .B2(n41), .ZN(n1408) );
  AOI22_X1 U1532 ( .A1(\REGISTERS[20][23] ), .A2(n1615), .B1(
        \REGISTERS[1][23] ), .B2(n39), .ZN(n1407) );
  AOI22_X1 U1533 ( .A1(\REGISTERS[6][23] ), .A2(n1616), .B1(
        \REGISTERS[17][23] ), .B2(n52), .ZN(n1406) );
  NAND4_X1 U1534 ( .A1(n1409), .A2(n1408), .A3(n1407), .A4(n1406), .ZN(n1425)
         );
  AOI22_X1 U1535 ( .A1(\REGISTERS[18][23] ), .A2(n1604), .B1(
        \REGISTERS[3][23] ), .B2(n50), .ZN(n1413) );
  AOI22_X1 U1536 ( .A1(\REGISTERS[19][23] ), .A2(n1603), .B1(
        \REGISTERS[29][23] ), .B2(n68), .ZN(n1412) );
  AOI22_X1 U1537 ( .A1(\REGISTERS[16][23] ), .A2(n1612), .B1(
        \REGISTERS[30][23] ), .B2(n65), .ZN(n1411) );
  AOI22_X1 U1538 ( .A1(\REGISTERS[27][23] ), .A2(n1577), .B1(
        \REGISTERS[21][23] ), .B2(n53), .ZN(n1410) );
  NAND4_X1 U1539 ( .A1(n1413), .A2(n1412), .A3(n1411), .A4(n1410), .ZN(n1424)
         );
  AOI22_X1 U1540 ( .A1(\REGISTERS[9][23] ), .A2(n1579), .B1(
        \REGISTERS[31][23] ), .B2(n54), .ZN(n1417) );
  AOI22_X1 U1541 ( .A1(\REGISTERS[22][23] ), .A2(n1592), .B1(
        \REGISTERS[12][23] ), .B2(n56), .ZN(n1416) );
  AOI22_X1 U1542 ( .A1(\REGISTERS[0][23] ), .A2(n64), .B1(\REGISTERS[24][23] ), 
        .B2(n47), .ZN(n1415) );
  AOI22_X1 U1543 ( .A1(\REGISTERS[5][23] ), .A2(n62), .B1(\REGISTERS[11][23] ), 
        .B2(n49), .ZN(n1414) );
  NAND4_X1 U1544 ( .A1(n1417), .A2(n1416), .A3(n1415), .A4(n1414), .ZN(n1423)
         );
  AOI22_X1 U1545 ( .A1(\REGISTERS[28][23] ), .A2(n1605), .B1(
        \REGISTERS[15][23] ), .B2(n55), .ZN(n1421) );
  AOI22_X1 U1546 ( .A1(\REGISTERS[8][23] ), .A2(n38), .B1(\REGISTERS[23][23] ), 
        .B2(n48), .ZN(n1420) );
  AOI22_X1 U1547 ( .A1(\REGISTERS[26][23] ), .A2(n1602), .B1(
        \REGISTERS[13][23] ), .B2(n45), .ZN(n1419) );
  AOI22_X1 U1548 ( .A1(\REGISTERS[7][23] ), .A2(n1580), .B1(
        \REGISTERS[25][23] ), .B2(n61), .ZN(n1418) );
  NAND4_X1 U1549 ( .A1(n1421), .A2(n1420), .A3(n1419), .A4(n1418), .ZN(n1422)
         );
  NOR4_X1 U1550 ( .A1(n1425), .A2(n1424), .A3(n1423), .A4(n1422), .ZN(n1426)
         );
  AOI22_X1 U1551 ( .A1(n69), .A2(n90), .B1(n1426), .B2(n72), .ZN(N402) );
  AOI22_X1 U1552 ( .A1(\REGISTERS[8][24] ), .A2(n1575), .B1(\REGISTERS[4][24] ), .B2(n37), .ZN(n1430) );
  AOI22_X1 U1553 ( .A1(\REGISTERS[5][24] ), .A2(n62), .B1(\REGISTERS[1][24] ), 
        .B2(n39), .ZN(n1429) );
  AOI22_X1 U1554 ( .A1(\REGISTERS[25][24] ), .A2(n1610), .B1(
        \REGISTERS[20][24] ), .B2(n66), .ZN(n1428) );
  AOI22_X1 U1555 ( .A1(\REGISTERS[22][24] ), .A2(n1592), .B1(
        \REGISTERS[24][24] ), .B2(n47), .ZN(n1427) );
  NAND4_X1 U1556 ( .A1(n1430), .A2(n1429), .A3(n1428), .A4(n1427), .ZN(n1446)
         );
  AOI22_X1 U1557 ( .A1(\REGISTERS[0][24] ), .A2(n1613), .B1(
        \REGISTERS[28][24] ), .B2(n60), .ZN(n1434) );
  AOI22_X1 U1558 ( .A1(\REGISTERS[19][24] ), .A2(n1603), .B1(
        \REGISTERS[11][24] ), .B2(n49), .ZN(n1433) );
  AOI22_X1 U1559 ( .A1(\REGISTERS[12][24] ), .A2(n1601), .B1(
        \REGISTERS[9][24] ), .B2(n42), .ZN(n1432) );
  AOI22_X1 U1560 ( .A1(\REGISTERS[17][24] ), .A2(n52), .B1(\REGISTERS[21][24] ), .B2(n53), .ZN(n1431) );
  NAND4_X1 U1561 ( .A1(n1434), .A2(n1433), .A3(n1432), .A4(n1431), .ZN(n1445)
         );
  AOI22_X1 U1562 ( .A1(\REGISTERS[27][24] ), .A2(n40), .B1(\REGISTERS[3][24] ), 
        .B2(n50), .ZN(n1438) );
  AOI22_X1 U1563 ( .A1(\REGISTERS[16][24] ), .A2(n1612), .B1(
        \REGISTERS[15][24] ), .B2(n55), .ZN(n1437) );
  AOI22_X1 U1564 ( .A1(\REGISTERS[29][24] ), .A2(n1617), .B1(
        \REGISTERS[6][24] ), .B2(n67), .ZN(n1436) );
  AOI22_X1 U1565 ( .A1(\REGISTERS[30][24] ), .A2(n65), .B1(\REGISTERS[18][24] ), .B2(n59), .ZN(n1435) );
  NAND4_X1 U1566 ( .A1(n1438), .A2(n1437), .A3(n1436), .A4(n1435), .ZN(n1444)
         );
  AOI22_X1 U1567 ( .A1(\REGISTERS[14][24] ), .A2(n1581), .B1(
        \REGISTERS[7][24] ), .B2(n43), .ZN(n1442) );
  AOI22_X1 U1568 ( .A1(\REGISTERS[26][24] ), .A2(n57), .B1(\REGISTERS[13][24] ), .B2(n45), .ZN(n1441) );
  AOI22_X1 U1569 ( .A1(\REGISTERS[2][24] ), .A2(n46), .B1(\REGISTERS[31][24] ), 
        .B2(n54), .ZN(n1440) );
  AOI22_X1 U1570 ( .A1(\REGISTERS[10][24] ), .A2(n41), .B1(\REGISTERS[23][24] ), .B2(n48), .ZN(n1439) );
  NAND4_X1 U1571 ( .A1(n1442), .A2(n1441), .A3(n1440), .A4(n1439), .ZN(n1443)
         );
  NOR4_X1 U1572 ( .A1(n1446), .A2(n1445), .A3(n1444), .A4(n1443), .ZN(n1447)
         );
  AOI22_X1 U1573 ( .A1(n70), .A2(n1780), .B1(n1447), .B2(n72), .ZN(N403) );
  AOI22_X1 U1574 ( .A1(\REGISTERS[14][25] ), .A2(n44), .B1(\REGISTERS[22][25] ), .B2(n51), .ZN(n1451) );
  AOI22_X1 U1575 ( .A1(\REGISTERS[23][25] ), .A2(n1589), .B1(
        \REGISTERS[29][25] ), .B2(n68), .ZN(n1450) );
  AOI22_X1 U1576 ( .A1(\REGISTERS[27][25] ), .A2(n1577), .B1(
        \REGISTERS[4][25] ), .B2(n37), .ZN(n1449) );
  AOI22_X1 U1577 ( .A1(\REGISTERS[24][25] ), .A2(n1588), .B1(
        \REGISTERS[10][25] ), .B2(n41), .ZN(n1448) );
  NAND4_X1 U1578 ( .A1(n1451), .A2(n1450), .A3(n1449), .A4(n1448), .ZN(n1467)
         );
  AOI22_X1 U1579 ( .A1(\REGISTERS[25][25] ), .A2(n61), .B1(\REGISTERS[1][25] ), 
        .B2(n39), .ZN(n1455) );
  AOI22_X1 U1580 ( .A1(\REGISTERS[26][25] ), .A2(n1602), .B1(
        \REGISTERS[0][25] ), .B2(n64), .ZN(n1454) );
  AOI22_X1 U1581 ( .A1(\REGISTERS[18][25] ), .A2(n59), .B1(\REGISTERS[9][25] ), 
        .B2(n42), .ZN(n1453) );
  AOI22_X1 U1582 ( .A1(\REGISTERS[3][25] ), .A2(n50), .B1(\REGISTERS[6][25] ), 
        .B2(n67), .ZN(n1452) );
  NAND4_X1 U1583 ( .A1(n1455), .A2(n1454), .A3(n1453), .A4(n1452), .ZN(n1466)
         );
  AOI22_X1 U1584 ( .A1(\REGISTERS[8][25] ), .A2(n38), .B1(\REGISTERS[12][25] ), 
        .B2(n56), .ZN(n1459) );
  AOI22_X1 U1585 ( .A1(\REGISTERS[17][25] ), .A2(n1593), .B1(
        \REGISTERS[16][25] ), .B2(n63), .ZN(n1458) );
  AOI22_X1 U1586 ( .A1(\REGISTERS[11][25] ), .A2(n1590), .B1(
        \REGISTERS[31][25] ), .B2(n54), .ZN(n1457) );
  AOI22_X1 U1587 ( .A1(\REGISTERS[2][25] ), .A2(n46), .B1(\REGISTERS[13][25] ), 
        .B2(n45), .ZN(n1456) );
  NAND4_X1 U1588 ( .A1(n1459), .A2(n1458), .A3(n1457), .A4(n1456), .ZN(n1465)
         );
  AOI22_X1 U1589 ( .A1(\REGISTERS[19][25] ), .A2(n58), .B1(\REGISTERS[7][25] ), 
        .B2(n43), .ZN(n1463) );
  AOI22_X1 U1590 ( .A1(\REGISTERS[5][25] ), .A2(n1611), .B1(
        \REGISTERS[28][25] ), .B2(n60), .ZN(n1462) );
  AOI22_X1 U1591 ( .A1(\REGISTERS[30][25] ), .A2(n1614), .B1(
        \REGISTERS[15][25] ), .B2(n55), .ZN(n1461) );
  AOI22_X1 U1592 ( .A1(\REGISTERS[20][25] ), .A2(n66), .B1(\REGISTERS[21][25] ), .B2(n53), .ZN(n1460) );
  NAND4_X1 U1593 ( .A1(n1463), .A2(n1462), .A3(n1461), .A4(n1460), .ZN(n1464)
         );
  NOR4_X1 U1594 ( .A1(n1467), .A2(n1466), .A3(n1465), .A4(n1464), .ZN(n1468)
         );
  AOI22_X1 U1595 ( .A1(n70), .A2(n86), .B1(n1468), .B2(n71), .ZN(N404) );
  AOI22_X1 U1596 ( .A1(\REGISTERS[12][26] ), .A2(n56), .B1(\REGISTERS[10][26] ), .B2(n41), .ZN(n1472) );
  AOI22_X1 U1597 ( .A1(\REGISTERS[15][26] ), .A2(n1600), .B1(
        \REGISTERS[0][26] ), .B2(n64), .ZN(n1471) );
  AOI22_X1 U1598 ( .A1(\REGISTERS[1][26] ), .A2(n39), .B1(\REGISTERS[4][26] ), 
        .B2(n37), .ZN(n1470) );
  AOI22_X1 U1599 ( .A1(\REGISTERS[28][26] ), .A2(n60), .B1(\REGISTERS[23][26] ), .B2(n48), .ZN(n1469) );
  NAND4_X1 U1600 ( .A1(n1472), .A2(n1471), .A3(n1470), .A4(n1469), .ZN(n1488)
         );
  AOI22_X1 U1601 ( .A1(\REGISTERS[22][26] ), .A2(n1592), .B1(
        \REGISTERS[6][26] ), .B2(n67), .ZN(n1476) );
  AOI22_X1 U1602 ( .A1(\REGISTERS[25][26] ), .A2(n1610), .B1(
        \REGISTERS[27][26] ), .B2(n40), .ZN(n1475) );
  AOI22_X1 U1603 ( .A1(\REGISTERS[19][26] ), .A2(n1603), .B1(
        \REGISTERS[17][26] ), .B2(n52), .ZN(n1474) );
  AOI22_X1 U1604 ( .A1(\REGISTERS[24][26] ), .A2(n1588), .B1(
        \REGISTERS[30][26] ), .B2(n65), .ZN(n1473) );
  NAND4_X1 U1605 ( .A1(n1476), .A2(n1475), .A3(n1474), .A4(n1473), .ZN(n1487)
         );
  AOI22_X1 U1606 ( .A1(\REGISTERS[16][26] ), .A2(n1612), .B1(
        \REGISTERS[11][26] ), .B2(n49), .ZN(n1480) );
  AOI22_X1 U1607 ( .A1(\REGISTERS[3][26] ), .A2(n1591), .B1(
        \REGISTERS[18][26] ), .B2(n59), .ZN(n1479) );
  AOI22_X1 U1608 ( .A1(\REGISTERS[9][26] ), .A2(n42), .B1(\REGISTERS[7][26] ), 
        .B2(n43), .ZN(n1478) );
  AOI22_X1 U1609 ( .A1(\REGISTERS[31][26] ), .A2(n54), .B1(\REGISTERS[14][26] ), .B2(n44), .ZN(n1477) );
  NAND4_X1 U1610 ( .A1(n1480), .A2(n1479), .A3(n1478), .A4(n1477), .ZN(n1486)
         );
  AOI22_X1 U1611 ( .A1(\REGISTERS[21][26] ), .A2(n53), .B1(\REGISTERS[8][26] ), 
        .B2(n38), .ZN(n1484) );
  AOI22_X1 U1612 ( .A1(\REGISTERS[20][26] ), .A2(n1615), .B1(
        \REGISTERS[2][26] ), .B2(n46), .ZN(n1483) );
  AOI22_X1 U1613 ( .A1(\REGISTERS[13][26] ), .A2(n1586), .B1(
        \REGISTERS[5][26] ), .B2(n62), .ZN(n1482) );
  AOI22_X1 U1614 ( .A1(\REGISTERS[29][26] ), .A2(n68), .B1(\REGISTERS[26][26] ), .B2(n57), .ZN(n1481) );
  NAND4_X1 U1615 ( .A1(n1484), .A2(n1483), .A3(n1482), .A4(n1481), .ZN(n1485)
         );
  NOR4_X1 U1616 ( .A1(n1488), .A2(n1487), .A3(n1486), .A4(n1485), .ZN(n1489)
         );
  AOI22_X1 U1617 ( .A1(n70), .A2(n84), .B1(n1489), .B2(n71), .ZN(N405) );
  AOI22_X1 U1618 ( .A1(\REGISTERS[26][27] ), .A2(n57), .B1(\REGISTERS[7][27] ), 
        .B2(n43), .ZN(n1493) );
  AOI22_X1 U1619 ( .A1(\REGISTERS[9][27] ), .A2(n1579), .B1(
        \REGISTERS[20][27] ), .B2(n66), .ZN(n1492) );
  AOI22_X1 U1620 ( .A1(\REGISTERS[18][27] ), .A2(n1604), .B1(
        \REGISTERS[27][27] ), .B2(n40), .ZN(n1491) );
  AOI22_X1 U1621 ( .A1(\REGISTERS[31][27] ), .A2(n1599), .B1(
        \REGISTERS[0][27] ), .B2(n64), .ZN(n1490) );
  NAND4_X1 U1622 ( .A1(n1493), .A2(n1492), .A3(n1491), .A4(n1490), .ZN(n1509)
         );
  AOI22_X1 U1623 ( .A1(\REGISTERS[2][27] ), .A2(n46), .B1(\REGISTERS[29][27] ), 
        .B2(n68), .ZN(n1497) );
  AOI22_X1 U1624 ( .A1(\REGISTERS[1][27] ), .A2(n1576), .B1(
        \REGISTERS[19][27] ), .B2(n58), .ZN(n1496) );
  AOI22_X1 U1625 ( .A1(\REGISTERS[5][27] ), .A2(n1611), .B1(
        \REGISTERS[22][27] ), .B2(n51), .ZN(n1495) );
  AOI22_X1 U1626 ( .A1(\REGISTERS[15][27] ), .A2(n1600), .B1(
        \REGISTERS[14][27] ), .B2(n44), .ZN(n1494) );
  NAND4_X1 U1627 ( .A1(n1497), .A2(n1496), .A3(n1495), .A4(n1494), .ZN(n1508)
         );
  AOI22_X1 U1628 ( .A1(\REGISTERS[10][27] ), .A2(n1578), .B1(
        \REGISTERS[6][27] ), .B2(n67), .ZN(n1501) );
  AOI22_X1 U1629 ( .A1(\REGISTERS[11][27] ), .A2(n1590), .B1(
        \REGISTERS[30][27] ), .B2(n65), .ZN(n1500) );
  AOI22_X1 U1630 ( .A1(\REGISTERS[3][27] ), .A2(n1591), .B1(
        \REGISTERS[25][27] ), .B2(n61), .ZN(n1499) );
  AOI22_X1 U1631 ( .A1(\REGISTERS[16][27] ), .A2(n1612), .B1(
        \REGISTERS[8][27] ), .B2(n38), .ZN(n1498) );
  NAND4_X1 U1632 ( .A1(n1501), .A2(n1500), .A3(n1499), .A4(n1498), .ZN(n1507)
         );
  AOI22_X1 U1633 ( .A1(\REGISTERS[17][27] ), .A2(n52), .B1(\REGISTERS[28][27] ), .B2(n60), .ZN(n1505) );
  AOI22_X1 U1634 ( .A1(\REGISTERS[12][27] ), .A2(n1601), .B1(
        \REGISTERS[24][27] ), .B2(n47), .ZN(n1504) );
  AOI22_X1 U1635 ( .A1(\REGISTERS[13][27] ), .A2(n45), .B1(\REGISTERS[4][27] ), 
        .B2(n37), .ZN(n1503) );
  AOI22_X1 U1636 ( .A1(\REGISTERS[23][27] ), .A2(n1589), .B1(
        \REGISTERS[21][27] ), .B2(n53), .ZN(n1502) );
  NAND4_X1 U1637 ( .A1(n1505), .A2(n1504), .A3(n1503), .A4(n1502), .ZN(n1506)
         );
  NOR4_X1 U1638 ( .A1(n1509), .A2(n1508), .A3(n1507), .A4(n1506), .ZN(n1510)
         );
  AOI22_X1 U1639 ( .A1(n70), .A2(n1779), .B1(n1510), .B2(n71), .ZN(N406) );
  AOI22_X1 U1640 ( .A1(\REGISTERS[20][28] ), .A2(n66), .B1(\REGISTERS[19][28] ), .B2(n58), .ZN(n1514) );
  AOI22_X1 U1641 ( .A1(\REGISTERS[4][28] ), .A2(n1574), .B1(
        \REGISTERS[28][28] ), .B2(n60), .ZN(n1513) );
  AOI22_X1 U1642 ( .A1(\REGISTERS[6][28] ), .A2(n1616), .B1(
        \REGISTERS[29][28] ), .B2(n68), .ZN(n1512) );
  AOI22_X1 U1643 ( .A1(\REGISTERS[21][28] ), .A2(n1598), .B1(
        \REGISTERS[30][28] ), .B2(n65), .ZN(n1511) );
  NAND4_X1 U1644 ( .A1(n1514), .A2(n1513), .A3(n1512), .A4(n1511), .ZN(n1530)
         );
  AOI22_X1 U1645 ( .A1(\REGISTERS[13][28] ), .A2(n1586), .B1(
        \REGISTERS[16][28] ), .B2(n63), .ZN(n1518) );
  AOI22_X1 U1646 ( .A1(\REGISTERS[24][28] ), .A2(n1588), .B1(
        \REGISTERS[14][28] ), .B2(n44), .ZN(n1517) );
  AOI22_X1 U1647 ( .A1(\REGISTERS[12][28] ), .A2(n56), .B1(\REGISTERS[23][28] ), .B2(n48), .ZN(n1516) );
  AOI22_X1 U1648 ( .A1(\REGISTERS[9][28] ), .A2(n42), .B1(\REGISTERS[7][28] ), 
        .B2(n43), .ZN(n1515) );
  NAND4_X1 U1649 ( .A1(n1518), .A2(n1517), .A3(n1516), .A4(n1515), .ZN(n1529)
         );
  AOI22_X1 U1650 ( .A1(\REGISTERS[18][28] ), .A2(n59), .B1(\REGISTERS[17][28] ), .B2(n52), .ZN(n1522) );
  AOI22_X1 U1651 ( .A1(\REGISTERS[8][28] ), .A2(n1575), .B1(\REGISTERS[5][28] ), .B2(n62), .ZN(n1521) );
  AOI22_X1 U1652 ( .A1(\REGISTERS[11][28] ), .A2(n1590), .B1(
        \REGISTERS[26][28] ), .B2(n57), .ZN(n1520) );
  AOI22_X1 U1653 ( .A1(\REGISTERS[15][28] ), .A2(n1600), .B1(
        \REGISTERS[3][28] ), .B2(n50), .ZN(n1519) );
  NAND4_X1 U1654 ( .A1(n1522), .A2(n1521), .A3(n1520), .A4(n1519), .ZN(n1528)
         );
  AOI22_X1 U1655 ( .A1(\REGISTERS[0][28] ), .A2(n64), .B1(\REGISTERS[10][28] ), 
        .B2(n41), .ZN(n1526) );
  AOI22_X1 U1656 ( .A1(\REGISTERS[2][28] ), .A2(n1587), .B1(\REGISTERS[1][28] ), .B2(n39), .ZN(n1525) );
  AOI22_X1 U1657 ( .A1(\REGISTERS[22][28] ), .A2(n1592), .B1(
        \REGISTERS[25][28] ), .B2(n61), .ZN(n1524) );
  AOI22_X1 U1658 ( .A1(\REGISTERS[27][28] ), .A2(n40), .B1(\REGISTERS[31][28] ), .B2(n54), .ZN(n1523) );
  NAND4_X1 U1659 ( .A1(n1526), .A2(n1525), .A3(n1524), .A4(n1523), .ZN(n1527)
         );
  NOR4_X1 U1660 ( .A1(n1530), .A2(n1529), .A3(n1528), .A4(n1527), .ZN(n1531)
         );
  AOI22_X1 U1661 ( .A1(n70), .A2(n80), .B1(n1531), .B2(n71), .ZN(N407) );
  AOI22_X1 U1662 ( .A1(\REGISTERS[24][29] ), .A2(n47), .B1(\REGISTERS[9][29] ), 
        .B2(n42), .ZN(n1535) );
  AOI22_X1 U1663 ( .A1(\REGISTERS[10][29] ), .A2(n41), .B1(\REGISTERS[26][29] ), .B2(n57), .ZN(n1534) );
  AOI22_X1 U1664 ( .A1(\REGISTERS[20][29] ), .A2(n1615), .B1(
        \REGISTERS[23][29] ), .B2(n48), .ZN(n1533) );
  AOI22_X1 U1665 ( .A1(\REGISTERS[8][29] ), .A2(n38), .B1(\REGISTERS[12][29] ), 
        .B2(n56), .ZN(n1532) );
  NAND4_X1 U1666 ( .A1(n1535), .A2(n1534), .A3(n1533), .A4(n1532), .ZN(n1551)
         );
  AOI22_X1 U1667 ( .A1(\REGISTERS[17][29] ), .A2(n1593), .B1(
        \REGISTERS[30][29] ), .B2(n65), .ZN(n1539) );
  AOI22_X1 U1668 ( .A1(\REGISTERS[19][29] ), .A2(n58), .B1(\REGISTERS[2][29] ), 
        .B2(n46), .ZN(n1538) );
  AOI22_X1 U1669 ( .A1(\REGISTERS[16][29] ), .A2(n63), .B1(\REGISTERS[6][29] ), 
        .B2(n67), .ZN(n1537) );
  AOI22_X1 U1670 ( .A1(\REGISTERS[3][29] ), .A2(n1591), .B1(
        \REGISTERS[14][29] ), .B2(n44), .ZN(n1536) );
  NAND4_X1 U1671 ( .A1(n1539), .A2(n1538), .A3(n1537), .A4(n1536), .ZN(n1550)
         );
  AOI22_X1 U1672 ( .A1(\REGISTERS[0][29] ), .A2(n1613), .B1(
        \REGISTERS[31][29] ), .B2(n54), .ZN(n1543) );
  AOI22_X1 U1673 ( .A1(\REGISTERS[28][29] ), .A2(n1605), .B1(
        \REGISTERS[13][29] ), .B2(n45), .ZN(n1542) );
  AOI22_X1 U1674 ( .A1(\REGISTERS[15][29] ), .A2(n55), .B1(\REGISTERS[11][29] ), .B2(n49), .ZN(n1541) );
  AOI22_X1 U1675 ( .A1(\REGISTERS[4][29] ), .A2(n1574), .B1(
        \REGISTERS[27][29] ), .B2(n40), .ZN(n1540) );
  NAND4_X1 U1676 ( .A1(n1543), .A2(n1542), .A3(n1541), .A4(n1540), .ZN(n1549)
         );
  AOI22_X1 U1677 ( .A1(\REGISTERS[25][29] ), .A2(n61), .B1(\REGISTERS[18][29] ), .B2(n59), .ZN(n1547) );
  AOI22_X1 U1678 ( .A1(\REGISTERS[22][29] ), .A2(n1592), .B1(
        \REGISTERS[29][29] ), .B2(n68), .ZN(n1546) );
  AOI22_X1 U1679 ( .A1(\REGISTERS[5][29] ), .A2(n1611), .B1(\REGISTERS[7][29] ), .B2(n43), .ZN(n1545) );
  AOI22_X1 U1680 ( .A1(\REGISTERS[1][29] ), .A2(n39), .B1(\REGISTERS[21][29] ), 
        .B2(n53), .ZN(n1544) );
  NAND4_X1 U1681 ( .A1(n1547), .A2(n1546), .A3(n1545), .A4(n1544), .ZN(n1548)
         );
  NOR4_X1 U1682 ( .A1(n1551), .A2(n1550), .A3(n1549), .A4(n1548), .ZN(n1552)
         );
  AOI22_X1 U1683 ( .A1(n70), .A2(n1777), .B1(n1552), .B2(n71), .ZN(N408) );
  AOI22_X1 U1684 ( .A1(\REGISTERS[16][30] ), .A2(n63), .B1(\REGISTERS[17][30] ), .B2(n52), .ZN(n1556) );
  AOI22_X1 U1685 ( .A1(\REGISTERS[30][30] ), .A2(n1614), .B1(
        \REGISTERS[4][30] ), .B2(n37), .ZN(n1555) );
  AOI22_X1 U1686 ( .A1(\REGISTERS[22][30] ), .A2(n51), .B1(\REGISTERS[27][30] ), .B2(n40), .ZN(n1554) );
  AOI22_X1 U1687 ( .A1(\REGISTERS[23][30] ), .A2(n1589), .B1(
        \REGISTERS[8][30] ), .B2(n38), .ZN(n1553) );
  NAND4_X1 U1688 ( .A1(n1556), .A2(n1555), .A3(n1554), .A4(n1553), .ZN(n1572)
         );
  AOI22_X1 U1689 ( .A1(\REGISTERS[3][30] ), .A2(n50), .B1(\REGISTERS[28][30] ), 
        .B2(n60), .ZN(n1560) );
  AOI22_X1 U1690 ( .A1(\REGISTERS[20][30] ), .A2(n66), .B1(\REGISTERS[14][30] ), .B2(n44), .ZN(n1559) );
  AOI22_X1 U1691 ( .A1(\REGISTERS[6][30] ), .A2(n67), .B1(\REGISTERS[11][30] ), 
        .B2(n49), .ZN(n1558) );
  AOI22_X1 U1692 ( .A1(\REGISTERS[13][30] ), .A2(n45), .B1(\REGISTERS[18][30] ), .B2(n59), .ZN(n1557) );
  NAND4_X1 U1693 ( .A1(n1560), .A2(n1559), .A3(n1558), .A4(n1557), .ZN(n1571)
         );
  AOI22_X1 U1694 ( .A1(\REGISTERS[15][30] ), .A2(n1600), .B1(
        \REGISTERS[21][30] ), .B2(n53), .ZN(n1564) );
  AOI22_X1 U1695 ( .A1(\REGISTERS[5][30] ), .A2(n1611), .B1(\REGISTERS[9][30] ), .B2(n42), .ZN(n1563) );
  AOI22_X1 U1696 ( .A1(\REGISTERS[31][30] ), .A2(n54), .B1(\REGISTERS[25][30] ), .B2(n61), .ZN(n1562) );
  AOI22_X1 U1697 ( .A1(\REGISTERS[12][30] ), .A2(n1601), .B1(
        \REGISTERS[0][30] ), .B2(n64), .ZN(n1561) );
  NAND4_X1 U1698 ( .A1(n1564), .A2(n1563), .A3(n1562), .A4(n1561), .ZN(n1570)
         );
  AOI22_X1 U1699 ( .A1(\REGISTERS[1][30] ), .A2(n1576), .B1(
        \REGISTERS[24][30] ), .B2(n47), .ZN(n1568) );
  AOI22_X1 U1700 ( .A1(\REGISTERS[26][30] ), .A2(n1602), .B1(
        \REGISTERS[2][30] ), .B2(n46), .ZN(n1567) );
  AOI22_X1 U1701 ( .A1(\REGISTERS[19][30] ), .A2(n1603), .B1(
        \REGISTERS[29][30] ), .B2(n68), .ZN(n1566) );
  AOI22_X1 U1702 ( .A1(\REGISTERS[10][30] ), .A2(n41), .B1(\REGISTERS[7][30] ), 
        .B2(n43), .ZN(n1565) );
  NAND4_X1 U1703 ( .A1(n1568), .A2(n1567), .A3(n1566), .A4(n1565), .ZN(n1569)
         );
  NOR4_X1 U1704 ( .A1(n1572), .A2(n1571), .A3(n1570), .A4(n1569), .ZN(n1573)
         );
  AOI22_X1 U1705 ( .A1(n70), .A2(n76), .B1(n1573), .B2(n71), .ZN(N409) );
  AOI22_X1 U1706 ( .A1(\REGISTERS[8][31] ), .A2(n1575), .B1(\REGISTERS[4][31] ), .B2(n37), .ZN(n1585) );
  AOI22_X1 U1707 ( .A1(\REGISTERS[27][31] ), .A2(n1577), .B1(
        \REGISTERS[1][31] ), .B2(n39), .ZN(n1584) );
  AOI22_X1 U1708 ( .A1(\REGISTERS[9][31] ), .A2(n1579), .B1(
        \REGISTERS[10][31] ), .B2(n41), .ZN(n1583) );
  AOI22_X1 U1709 ( .A1(\REGISTERS[14][31] ), .A2(n1581), .B1(
        \REGISTERS[7][31] ), .B2(n43), .ZN(n1582) );
  NAND4_X1 U1710 ( .A1(n1585), .A2(n1584), .A3(n1583), .A4(n1582), .ZN(n1625)
         );
  AOI22_X1 U1711 ( .A1(\REGISTERS[2][31] ), .A2(n46), .B1(\REGISTERS[13][31] ), 
        .B2(n45), .ZN(n1597) );
  AOI22_X1 U1712 ( .A1(\REGISTERS[23][31] ), .A2(n1589), .B1(
        \REGISTERS[24][31] ), .B2(n47), .ZN(n1596) );
  AOI22_X1 U1713 ( .A1(\REGISTERS[3][31] ), .A2(n50), .B1(\REGISTERS[11][31] ), 
        .B2(n49), .ZN(n1595) );
  AOI22_X1 U1714 ( .A1(\REGISTERS[17][31] ), .A2(n52), .B1(\REGISTERS[22][31] ), .B2(n51), .ZN(n1594) );
  NAND4_X1 U1715 ( .A1(n1597), .A2(n1596), .A3(n1595), .A4(n1594), .ZN(n1624)
         );
  AOI22_X1 U1716 ( .A1(\REGISTERS[31][31] ), .A2(n1599), .B1(
        \REGISTERS[21][31] ), .B2(n53), .ZN(n1609) );
  AOI22_X1 U1717 ( .A1(\REGISTERS[12][31] ), .A2(n1601), .B1(
        \REGISTERS[15][31] ), .B2(n55), .ZN(n1608) );
  AOI22_X1 U1718 ( .A1(\REGISTERS[19][31] ), .A2(n58), .B1(\REGISTERS[26][31] ), .B2(n57), .ZN(n1607) );
  AOI22_X1 U1719 ( .A1(\REGISTERS[28][31] ), .A2(n1605), .B1(
        \REGISTERS[18][31] ), .B2(n59), .ZN(n1606) );
  NAND4_X1 U1720 ( .A1(n1609), .A2(n1608), .A3(n1607), .A4(n1606), .ZN(n1623)
         );
  AOI22_X1 U1721 ( .A1(\REGISTERS[5][31] ), .A2(n62), .B1(\REGISTERS[25][31] ), 
        .B2(n61), .ZN(n1621) );
  AOI22_X1 U1722 ( .A1(\REGISTERS[0][31] ), .A2(n1613), .B1(
        \REGISTERS[16][31] ), .B2(n63), .ZN(n1620) );
  AOI22_X1 U1723 ( .A1(\REGISTERS[20][31] ), .A2(n1615), .B1(
        \REGISTERS[30][31] ), .B2(n65), .ZN(n1619) );
  AOI22_X1 U1724 ( .A1(\REGISTERS[29][31] ), .A2(n1617), .B1(
        \REGISTERS[6][31] ), .B2(n67), .ZN(n1618) );
  NAND4_X1 U1725 ( .A1(n1621), .A2(n1620), .A3(n1619), .A4(n1618), .ZN(n1622)
         );
  NOR4_X1 U1726 ( .A1(n1625), .A2(n1624), .A3(n1623), .A4(n1622), .ZN(n1626)
         );
  AOI22_X1 U1727 ( .A1(n70), .A2(n74), .B1(n1626), .B2(n71), .ZN(N410) );
  OAI21_X1 U1728 ( .B1(n1629), .B2(n1628), .A(RST), .ZN(N81) );
  INV_X2 U53 ( .A(n126), .ZN(n125) );
  BUF_X2 U9 ( .A(RST), .Z(n145) );
  BUF_X2 U6 ( .A(RST), .Z(n155) );
  BUF_X2 U8 ( .A(n150), .Z(n152) );
  BUF_X2 U4 ( .A(RST), .Z(n137) );
  BUF_X2 U11 ( .A(RST), .Z(n138) );
  BUF_X2 U7 ( .A(RST), .Z(n151) );
  BUF_X2 U15 ( .A(n153), .Z(n148) );
  BUF_X2 U10 ( .A(n153), .Z(n143) );
  BUF_X2 U17 ( .A(RST), .Z(n141) );
  BUF_X2 U3 ( .A(RST), .Z(n142) );
  BUF_X2 U12 ( .A(RST), .Z(n154) );
  BUF_X2 U5 ( .A(RST), .Z(n140) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n1776), .CK(net7260), .Q(
        \REGISTERS[31][0] ) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n1775), .CK(net7250), .Q(
        \REGISTERS[29][0] ) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n1774), .CK(net7240), .Q(
        \REGISTERS[27][0] ) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n1773), .CK(net7230), .Q(
        \REGISTERS[25][0] ) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n1772), .CK(net7220), .Q(
        \REGISTERS[23][0] ) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n1771), .CK(net7210), .Q(
        \REGISTERS[21][0] ) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n1770), .CK(net7205), .Q(
        \REGISTERS[20][0] ) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n1769), .CK(net7195), .Q(
        \REGISTERS[18][0] ) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n1768), .CK(net7185), .Q(
        \REGISTERS[16][0] ) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n1767), .CK(net7175), .Q(
        \REGISTERS[14][0] ) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n1766), .CK(net7170), .Q(
        \REGISTERS[13][0] ) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n1765), .CK(net7165), .Q(
        \REGISTERS[12][0] ) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n1764), .CK(net7160), .Q(
        \REGISTERS[11][0] ) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n1763), .CK(net7155), .Q(
        \REGISTERS[10][0] ) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n1762), .CK(net7150), .Q(\REGISTERS[9][0] ) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n1761), .CK(net7145), .Q(\REGISTERS[8][0] ) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n1760), .CK(net7260), .Q(
        \REGISTERS[31][7] ) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n1759), .CK(net7250), .Q(
        \REGISTERS[29][7] ) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n1758), .CK(net7240), .Q(
        \REGISTERS[27][7] ) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n1757), .CK(net7230), .Q(
        \REGISTERS[25][7] ) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n1756), .CK(net7220), .Q(
        \REGISTERS[23][7] ) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n1755), .CK(net7210), .Q(
        \REGISTERS[21][7] ) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n1754), .CK(net7205), .Q(
        \REGISTERS[20][7] ) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n1753), .CK(net7195), .Q(
        \REGISTERS[18][7] ) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n1752), .CK(net7185), .Q(
        \REGISTERS[16][7] ) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n1751), .CK(net7175), .Q(
        \REGISTERS[14][7] ) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n1750), .CK(net7170), .Q(
        \REGISTERS[13][7] ) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n1749), .CK(net7165), .Q(
        \REGISTERS[12][7] ) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n1748), .CK(net7160), .Q(
        \REGISTERS[11][7] ) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n1747), .CK(net7155), .Q(
        \REGISTERS[10][7] ) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n1746), .CK(net7150), .Q(\REGISTERS[9][7] ) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n1745), .CK(net7145), .Q(\REGISTERS[8][7] ) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n1744), .CK(net7260), .Q(
        \REGISTERS[31][15] ) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n1743), .CK(net7250), .Q(
        \REGISTERS[29][15] ) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n1742), .CK(net7240), .Q(
        \REGISTERS[27][15] ) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n1741), .CK(net7230), .Q(
        \REGISTERS[25][15] ) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n1740), .CK(net7220), .Q(
        \REGISTERS[23][15] ) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n1739), .CK(net7210), .Q(
        \REGISTERS[21][15] ) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n1738), .CK(net7205), .Q(
        \REGISTERS[20][15] ) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n1737), .CK(net7195), .Q(
        \REGISTERS[18][15] ) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n1736), .CK(net7185), .Q(
        \REGISTERS[16][15] ) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n1735), .CK(net7175), .Q(
        \REGISTERS[14][15] ) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n1734), .CK(net7170), .Q(
        \REGISTERS[13][15] ) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n1733), .CK(net7165), .Q(
        \REGISTERS[12][15] ) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n1732), .CK(net7160), .Q(
        \REGISTERS[11][15] ) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n1731), .CK(net7155), .Q(
        \REGISTERS[10][15] ) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n1730), .CK(net7150), .Q(
        \REGISTERS[9][15] ) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n1729), .CK(net7145), .Q(
        \REGISTERS[8][15] ) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n1728), .CK(net7205), .Q(
        \REGISTERS[20][16] ) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n1727), .CK(net7205), .Q(
        \REGISTERS[20][13] ) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n1726), .CK(net7205), .Q(
        \REGISTERS[20][11] ) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n1725), .CK(net7205), .Q(
        \REGISTERS[20][4] ) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n1724), .CK(net7195), .Q(
        \REGISTERS[18][16] ) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n1723), .CK(net7195), .Q(
        \REGISTERS[18][13] ) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n1722), .CK(net7195), .Q(
        \REGISTERS[18][11] ) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n1721), .CK(net7195), .Q(
        \REGISTERS[18][4] ) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n1720), .CK(net7185), .Q(
        \REGISTERS[16][16] ) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n1719), .CK(net7185), .Q(
        \REGISTERS[16][13] ) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n1718), .CK(net7185), .Q(
        \REGISTERS[16][11] ) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n1717), .CK(net7185), .Q(
        \REGISTERS[16][4] ) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n1716), .CK(net7175), .Q(
        \REGISTERS[14][16] ) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n1715), .CK(net7175), .Q(
        \REGISTERS[14][13] ) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n1714), .CK(net7175), .Q(
        \REGISTERS[14][11] ) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n1713), .CK(net7175), .Q(
        \REGISTERS[14][4] ) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n1712), .CK(net7170), .Q(
        \REGISTERS[13][16] ) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n1782), .CK(net7195), .Q(
        \REGISTERS[18][30] ) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n1784), .CK(net7195), .Q(
        \REGISTERS[18][23] ) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n1783), .CK(net7195), .Q(
        \REGISTERS[18][29] ) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n1788), .CK(net7195), .Q(
        \REGISTERS[18][21] ) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n1787), .CK(net7195), .Q(
        \REGISTERS[18][24] ) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n1786), .CK(net7195), .Q(
        \REGISTERS[18][27] ) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n1711), .CK(net7205), .Q(
        \REGISTERS[20][6] ) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n1785), .CK(net7195), .Q(
        \REGISTERS[18][1] ) );
  DFF_X2 \REGISTERS_reg[31][12]  ( .D(n1710), .CK(net7260), .Q(
        \REGISTERS[31][12] ) );
  DFF_X2 \REGISTERS_reg[30][12]  ( .D(n1709), .CK(net7255), .Q(
        \REGISTERS[30][12] ) );
  DFF_X2 \REGISTERS_reg[29][12]  ( .D(n1708), .CK(net7250), .Q(
        \REGISTERS[29][12] ) );
  DFF_X2 \REGISTERS_reg[28][12]  ( .D(n1707), .CK(net7245), .Q(
        \REGISTERS[28][12] ) );
  DFF_X2 \REGISTERS_reg[27][12]  ( .D(n1706), .CK(net7240), .Q(
        \REGISTERS[27][12] ) );
  DFF_X2 \REGISTERS_reg[26][12]  ( .D(n1705), .CK(net7235), .Q(
        \REGISTERS[26][12] ) );
  DFF_X2 \REGISTERS_reg[25][12]  ( .D(n1704), .CK(net7230), .Q(
        \REGISTERS[25][12] ) );
  DFF_X2 \REGISTERS_reg[24][12]  ( .D(n1703), .CK(net7225), .Q(
        \REGISTERS[24][12] ) );
  DFF_X2 \REGISTERS_reg[23][12]  ( .D(n1702), .CK(net7220), .Q(
        \REGISTERS[23][12] ) );
  DFF_X2 \REGISTERS_reg[22][12]  ( .D(n1701), .CK(net7215), .Q(
        \REGISTERS[22][12] ) );
  DFF_X2 \REGISTERS_reg[21][12]  ( .D(n1700), .CK(net7210), .Q(
        \REGISTERS[21][12] ) );
  DFF_X2 \REGISTERS_reg[19][12]  ( .D(n1699), .CK(net7200), .Q(
        \REGISTERS[19][12] ) );
  DFF_X2 \REGISTERS_reg[17][12]  ( .D(n1698), .CK(net7190), .Q(
        \REGISTERS[17][12] ) );
  DFF_X2 \REGISTERS_reg[15][12]  ( .D(n1697), .CK(net7180), .Q(
        \REGISTERS[15][12] ) );
  DFF_X2 \REGISTERS_reg[7][12]  ( .D(n1696), .CK(net7140), .Q(
        \REGISTERS[7][12] ) );
  DFF_X2 \REGISTERS_reg[6][12]  ( .D(n1695), .CK(net7135), .Q(
        \REGISTERS[6][12] ) );
  DFF_X2 \REGISTERS_reg[5][12]  ( .D(n1694), .CK(net7130), .Q(
        \REGISTERS[5][12] ) );
  DFF_X2 \REGISTERS_reg[4][12]  ( .D(n1693), .CK(net7125), .Q(
        \REGISTERS[4][12] ) );
  DFF_X2 \REGISTERS_reg[3][12]  ( .D(n1692), .CK(net7120), .Q(
        \REGISTERS[3][12] ) );
  DFF_X2 \REGISTERS_reg[2][12]  ( .D(n1691), .CK(net7115), .Q(
        \REGISTERS[2][12] ) );
  DFF_X2 \REGISTERS_reg[1][12]  ( .D(n1690), .CK(net7110), .Q(
        \REGISTERS[1][12] ) );
  DFF_X2 \REGISTERS_reg[0][12]  ( .D(n1689), .CK(net7104), .Q(
        \REGISTERS[0][12] ) );
  DFF_X2 \REGISTERS_reg[31][9]  ( .D(n1688), .CK(net7260), .Q(
        \REGISTERS[31][9] ) );
  DFF_X2 \REGISTERS_reg[30][9]  ( .D(n1687), .CK(net7255), .Q(
        \REGISTERS[30][9] ) );
  DFF_X2 \REGISTERS_reg[29][9]  ( .D(n1686), .CK(net7250), .Q(
        \REGISTERS[29][9] ) );
  DFF_X2 \REGISTERS_reg[28][9]  ( .D(n1685), .CK(net7245), .Q(
        \REGISTERS[28][9] ) );
  DFF_X2 \REGISTERS_reg[27][9]  ( .D(n1684), .CK(net7240), .Q(
        \REGISTERS[27][9] ) );
  DFF_X2 \REGISTERS_reg[26][9]  ( .D(n1683), .CK(net7235), .Q(
        \REGISTERS[26][9] ) );
  DFF_X2 \REGISTERS_reg[25][9]  ( .D(n1682), .CK(net7230), .Q(
        \REGISTERS[25][9] ) );
  DFF_X2 \REGISTERS_reg[24][9]  ( .D(n1681), .CK(net7225), .Q(
        \REGISTERS[24][9] ) );
  DFF_X2 \REGISTERS_reg[23][9]  ( .D(n1680), .CK(net7220), .Q(
        \REGISTERS[23][9] ) );
  DFF_X2 \REGISTERS_reg[22][9]  ( .D(n1679), .CK(net7215), .Q(
        \REGISTERS[22][9] ) );
  DFF_X2 \REGISTERS_reg[21][9]  ( .D(n1678), .CK(net7210), .Q(
        \REGISTERS[21][9] ) );
  DFF_X2 \REGISTERS_reg[19][9]  ( .D(n1677), .CK(net7200), .Q(
        \REGISTERS[19][9] ) );
  DFF_X2 \REGISTERS_reg[17][9]  ( .D(n1676), .CK(net7190), .Q(
        \REGISTERS[17][9] ) );
  DFF_X2 \REGISTERS_reg[15][9]  ( .D(n1675), .CK(net7180), .Q(
        \REGISTERS[15][9] ) );
  DFF_X2 \REGISTERS_reg[7][9]  ( .D(n1674), .CK(net7140), .Q(\REGISTERS[7][9] ) );
  DFF_X2 \REGISTERS_reg[6][9]  ( .D(n1673), .CK(net7135), .Q(\REGISTERS[6][9] ) );
  DFF_X2 \REGISTERS_reg[5][9]  ( .D(n1672), .CK(net7130), .Q(\REGISTERS[5][9] ) );
  DFF_X2 \REGISTERS_reg[4][9]  ( .D(n1671), .CK(net7125), .Q(\REGISTERS[4][9] ) );
  DFF_X2 \REGISTERS_reg[3][9]  ( .D(n1670), .CK(net7120), .Q(\REGISTERS[3][9] ) );
  DFF_X2 \REGISTERS_reg[2][9]  ( .D(n1669), .CK(net7115), .Q(\REGISTERS[2][9] ) );
  DFF_X2 \REGISTERS_reg[1][9]  ( .D(n1668), .CK(net7110), .Q(\REGISTERS[1][9] ) );
  DFF_X2 \REGISTERS_reg[0][9]  ( .D(n1667), .CK(net7104), .Q(\REGISTERS[0][9] ) );
  DFF_X2 \REGISTERS_reg[31][18]  ( .D(n1666), .CK(net7260), .Q(
        \REGISTERS[31][18] ) );
  DFF_X2 \REGISTERS_reg[30][18]  ( .D(n1665), .CK(net7255), .Q(
        \REGISTERS[30][18] ) );
  DFF_X2 \REGISTERS_reg[29][18]  ( .D(n1664), .CK(net7250), .Q(
        \REGISTERS[29][18] ) );
  DFF_X2 \REGISTERS_reg[28][18]  ( .D(n1663), .CK(net7245), .Q(
        \REGISTERS[28][18] ) );
  DFF_X2 \REGISTERS_reg[27][18]  ( .D(n1662), .CK(net7240), .Q(
        \REGISTERS[27][18] ) );
  DFF_X2 \REGISTERS_reg[26][18]  ( .D(n1661), .CK(net7235), .Q(
        \REGISTERS[26][18] ) );
  DFF_X2 \REGISTERS_reg[25][18]  ( .D(n1660), .CK(net7230), .Q(
        \REGISTERS[25][18] ) );
  DFF_X2 \REGISTERS_reg[24][18]  ( .D(n1659), .CK(net7225), .Q(
        \REGISTERS[24][18] ) );
  DFF_X2 \REGISTERS_reg[23][18]  ( .D(n1658), .CK(net7220), .Q(
        \REGISTERS[23][18] ) );
  DFF_X2 \REGISTERS_reg[22][18]  ( .D(n1657), .CK(net7215), .Q(
        \REGISTERS[22][18] ) );
  DFF_X2 \REGISTERS_reg[21][18]  ( .D(n1656), .CK(net7210), .Q(
        \REGISTERS[21][18] ) );
  DFF_X2 \REGISTERS_reg[19][18]  ( .D(n1655), .CK(net7200), .Q(
        \REGISTERS[19][18] ) );
  DFF_X2 \REGISTERS_reg[17][18]  ( .D(n1654), .CK(net7190), .Q(
        \REGISTERS[17][18] ) );
  DFF_X2 \REGISTERS_reg[15][18]  ( .D(n1653), .CK(net7180), .Q(
        \REGISTERS[15][18] ) );
  DFF_X2 \REGISTERS_reg[7][18]  ( .D(n1652), .CK(net7140), .Q(
        \REGISTERS[7][18] ) );
  DFF_X2 \REGISTERS_reg[6][18]  ( .D(n1651), .CK(net7135), .Q(
        \REGISTERS[6][18] ) );
  DFF_X2 \REGISTERS_reg[5][18]  ( .D(n1650), .CK(net7130), .Q(
        \REGISTERS[5][18] ) );
  DFF_X2 \REGISTERS_reg[4][18]  ( .D(n1649), .CK(net7125), .Q(
        \REGISTERS[4][18] ) );
  DFF_X2 \REGISTERS_reg[3][18]  ( .D(n1648), .CK(net7120), .Q(
        \REGISTERS[3][18] ) );
  DFF_X2 \REGISTERS_reg[2][18]  ( .D(n1647), .CK(net7115), .Q(
        \REGISTERS[2][18] ) );
  DFF_X2 \REGISTERS_reg[1][18]  ( .D(n1646), .CK(net7110), .Q(
        \REGISTERS[1][18] ) );
  BUF_X2 U14 ( .A(RST), .Z(n147) );
  CLKBUF_X3 U16 ( .A(DATAIN[14]), .Z(n1630) );
  CLKBUF_X3 U20 ( .A(DATAIN[3]), .Z(n1631) );
  INV_X4 U22 ( .A(n90), .ZN(n89) );
  INV_X4 U23 ( .A(n108), .ZN(n107) );
  CLKBUF_X3 U24 ( .A(DATAIN[5]), .Z(n1632) );
  INV_X4 U25 ( .A(n130), .ZN(n129) );
  INV_X2 U26 ( .A(n106), .ZN(n105) );
  INV_X1 U27 ( .A(n104), .ZN(n1633) );
  INV_X1 U28 ( .A(n110), .ZN(n1634) );
  INV_X1 U29 ( .A(n114), .ZN(n1635) );
  BUF_X4 U30 ( .A(DATAIN[10]), .Z(n1636) );
  NAND2_X1 U31 ( .A1(EN), .A2(n1795), .ZN(n164) );
  BUF_X1 U32 ( .A(DATAIN[29]), .Z(n1637) );
  CLKBUF_X3 U33 ( .A(DATAIN[29]), .Z(n1638) );
  BUF_X1 U34 ( .A(DATAIN[1]), .Z(n1639) );
  CLKBUF_X3 U35 ( .A(DATAIN[1]), .Z(n1640) );
  BUF_X2 U36 ( .A(DATAIN[27]), .Z(n1641) );
  BUF_X2 U37 ( .A(DATAIN[24]), .Z(n1642) );
  BUF_X2 U38 ( .A(DATAIN[21]), .Z(n1643) );
  BUF_X2 U39 ( .A(DATAIN[17]), .Z(n1644) );
  BUF_X2 U41 ( .A(DATAIN[19]), .Z(n1645) );
  CLKBUF_X2 U43 ( .A(RST), .Z(n150) );
  CLKBUF_X2 U44 ( .A(RST), .Z(n153) );
  AND2_X1 U46 ( .A1(n99), .A2(RST), .ZN(n1646) );
  AND2_X1 U47 ( .A1(n99), .A2(n154), .ZN(n1647) );
  AND2_X1 U48 ( .A1(n99), .A2(RST), .ZN(n1648) );
  AND2_X1 U49 ( .A1(n99), .A2(RST), .ZN(n1649) );
  AND2_X1 U50 ( .A1(n99), .A2(n155), .ZN(n1650) );
  AND2_X1 U51 ( .A1(n99), .A2(n151), .ZN(n1651) );
  AND2_X1 U52 ( .A1(n99), .A2(RST), .ZN(n1652) );
  AND2_X1 U168 ( .A1(n99), .A2(n143), .ZN(n1653) );
  AND2_X1 U184 ( .A1(n99), .A2(n150), .ZN(n1654) );
  AND2_X1 U193 ( .A1(n99), .A2(n137), .ZN(n1655) );
  AND2_X1 U202 ( .A1(n99), .A2(RST), .ZN(n1656) );
  AND2_X1 U1730 ( .A1(n99), .A2(n141), .ZN(n1657) );
  AND2_X1 U1731 ( .A1(n99), .A2(n140), .ZN(n1658) );
  AND2_X1 U1732 ( .A1(n99), .A2(n143), .ZN(n1659) );
  AND2_X1 U1733 ( .A1(n99), .A2(n148), .ZN(n1660) );
  AND2_X1 U1734 ( .A1(n99), .A2(RST), .ZN(n1661) );
  AND2_X1 U1735 ( .A1(n99), .A2(n141), .ZN(n1662) );
  AND2_X1 U1736 ( .A1(n99), .A2(n139), .ZN(n1663) );
  AND2_X1 U1737 ( .A1(n99), .A2(n137), .ZN(n1664) );
  AND2_X1 U1738 ( .A1(n99), .A2(n146), .ZN(n1665) );
  AND2_X1 U1739 ( .A1(n99), .A2(RST), .ZN(n1666) );
  AND2_X1 U1740 ( .A1(n117), .A2(n155), .ZN(n1667) );
  AND2_X1 U1741 ( .A1(n117), .A2(RST), .ZN(n1668) );
  AND2_X1 U1742 ( .A1(n117), .A2(n154), .ZN(n1669) );
  AND2_X1 U1743 ( .A1(n117), .A2(RST), .ZN(n1670) );
  AND2_X1 U1744 ( .A1(n117), .A2(RST), .ZN(n1671) );
  AND2_X1 U1745 ( .A1(n117), .A2(RST), .ZN(n1672) );
  AND2_X1 U1746 ( .A1(n117), .A2(n151), .ZN(n1673) );
  AND2_X1 U1747 ( .A1(n117), .A2(n143), .ZN(n1674) );
  AND2_X1 U1748 ( .A1(n117), .A2(n154), .ZN(n1675) );
  AND2_X1 U1749 ( .A1(n117), .A2(RST), .ZN(n1676) );
  AND2_X1 U1750 ( .A1(n117), .A2(n137), .ZN(n1677) );
  AND2_X1 U1751 ( .A1(n117), .A2(RST), .ZN(n1678) );
  AND2_X1 U1752 ( .A1(n117), .A2(n137), .ZN(n1679) );
  AND2_X1 U1753 ( .A1(n117), .A2(n138), .ZN(n1680) );
  AND2_X1 U1754 ( .A1(n117), .A2(n144), .ZN(n1681) );
  AND2_X1 U1755 ( .A1(n117), .A2(n140), .ZN(n1682) );
  AND2_X1 U1756 ( .A1(n117), .A2(RST), .ZN(n1683) );
  AND2_X1 U1757 ( .A1(n117), .A2(n141), .ZN(n1684) );
  AND2_X1 U1758 ( .A1(n117), .A2(n139), .ZN(n1685) );
  AND2_X1 U1759 ( .A1(n117), .A2(n137), .ZN(n1686) );
  AND2_X1 U1760 ( .A1(n117), .A2(RST), .ZN(n1687) );
  AND2_X1 U1761 ( .A1(n117), .A2(RST), .ZN(n1688) );
  AND2_X1 U1762 ( .A1(n111), .A2(n155), .ZN(n1689) );
  AND2_X1 U1763 ( .A1(n111), .A2(RST), .ZN(n1690) );
  AND2_X1 U1764 ( .A1(n111), .A2(n154), .ZN(n1691) );
  AND2_X1 U1765 ( .A1(n111), .A2(RST), .ZN(n1692) );
  AND2_X1 U1766 ( .A1(n111), .A2(RST), .ZN(n1693) );
  AND2_X1 U1767 ( .A1(n111), .A2(n144), .ZN(n1694) );
  AND2_X1 U1768 ( .A1(n111), .A2(n151), .ZN(n1695) );
  AND2_X1 U1769 ( .A1(n111), .A2(RST), .ZN(n1696) );
  AND2_X1 U1770 ( .A1(n111), .A2(RST), .ZN(n1697) );
  AND2_X1 U1771 ( .A1(n111), .A2(n152), .ZN(n1698) );
  AND2_X1 U1772 ( .A1(n111), .A2(RST), .ZN(n1699) );
  AND2_X1 U1773 ( .A1(n111), .A2(RST), .ZN(n1700) );
  AND2_X1 U1774 ( .A1(n111), .A2(RST), .ZN(n1701) );
  AND2_X1 U1775 ( .A1(n111), .A2(n139), .ZN(n1702) );
  AND2_X1 U1776 ( .A1(n111), .A2(n146), .ZN(n1703) );
  AND2_X1 U1777 ( .A1(n111), .A2(n142), .ZN(n1704) );
  AND2_X1 U1778 ( .A1(n111), .A2(n148), .ZN(n1705) );
  AND2_X1 U1779 ( .A1(n111), .A2(n141), .ZN(n1706) );
  AND2_X1 U1780 ( .A1(n111), .A2(n139), .ZN(n1707) );
  AND2_X1 U1781 ( .A1(n111), .A2(n137), .ZN(n1708) );
  AND2_X1 U1782 ( .A1(n111), .A2(RST), .ZN(n1709) );
  AND2_X1 U1783 ( .A1(n111), .A2(n146), .ZN(n1710) );
  AND2_X1 U1784 ( .A1(DATAIN[6]), .A2(n150), .ZN(n1711) );
  AND2_X1 U1785 ( .A1(n1633), .A2(n146), .ZN(n1712) );
  AND2_X1 U1786 ( .A1(DATAIN[4]), .A2(n144), .ZN(n1713) );
  AND2_X1 U1787 ( .A1(n1635), .A2(RST), .ZN(n1714) );
  AND2_X1 U1788 ( .A1(n1634), .A2(RST), .ZN(n1715) );
  AND2_X1 U1789 ( .A1(n1633), .A2(n148), .ZN(n1716) );
  AND2_X1 U1790 ( .A1(DATAIN[4]), .A2(n143), .ZN(n1717) );
  AND2_X1 U1791 ( .A1(n1635), .A2(n154), .ZN(n1718) );
  AND2_X1 U1792 ( .A1(n1634), .A2(RST), .ZN(n1719) );
  AND2_X1 U1793 ( .A1(n1633), .A2(n150), .ZN(n1720) );
  AND2_X1 U1794 ( .A1(DATAIN[4]), .A2(RST), .ZN(n1721) );
  AND2_X1 U1795 ( .A1(n1635), .A2(RST), .ZN(n1722) );
  AND2_X1 U1796 ( .A1(n1634), .A2(n138), .ZN(n1723) );
  AND2_X1 U1797 ( .A1(n1633), .A2(RST), .ZN(n1724) );
  AND2_X1 U1798 ( .A1(DATAIN[4]), .A2(RST), .ZN(n1725) );
  AND2_X1 U1799 ( .A1(n1635), .A2(RST), .ZN(n1726) );
  AND2_X1 U1800 ( .A1(n1634), .A2(RST), .ZN(n1727) );
  AND2_X1 U1801 ( .A1(n1633), .A2(n146), .ZN(n1728) );
  AND2_X1 U1802 ( .A1(DATAIN[15]), .A2(RST), .ZN(n1729) );
  AND2_X1 U1803 ( .A1(DATAIN[15]), .A2(n149), .ZN(n1730) );
  AND2_X1 U1804 ( .A1(DATAIN[15]), .A2(n147), .ZN(n1731) );
  AND2_X1 U1805 ( .A1(DATAIN[15]), .A2(RST), .ZN(n1732) );
  AND2_X1 U1806 ( .A1(DATAIN[15]), .A2(n154), .ZN(n1733) );
  AND2_X1 U1807 ( .A1(DATAIN[15]), .A2(n146), .ZN(n1734) );
  AND2_X1 U1808 ( .A1(DATAIN[15]), .A2(n149), .ZN(n1735) );
  AND2_X1 U1809 ( .A1(DATAIN[15]), .A2(RST), .ZN(n1736) );
  AND2_X1 U1810 ( .A1(DATAIN[15]), .A2(n148), .ZN(n1737) );
  AND2_X1 U1811 ( .A1(DATAIN[15]), .A2(RST), .ZN(n1738) );
  AND2_X1 U1812 ( .A1(DATAIN[15]), .A2(RST), .ZN(n1739) );
  AND2_X1 U1813 ( .A1(DATAIN[15]), .A2(RST), .ZN(n1740) );
  AND2_X1 U1814 ( .A1(DATAIN[15]), .A2(n138), .ZN(n1741) );
  AND2_X1 U1815 ( .A1(DATAIN[15]), .A2(n141), .ZN(n1742) );
  AND2_X1 U1816 ( .A1(DATAIN[15]), .A2(n137), .ZN(n1743) );
  AND2_X1 U1817 ( .A1(DATAIN[15]), .A2(RST), .ZN(n1744) );
  AND2_X1 U1818 ( .A1(DATAIN[7]), .A2(n147), .ZN(n1745) );
  AND2_X1 U1819 ( .A1(DATAIN[7]), .A2(n149), .ZN(n1746) );
  AND2_X1 U1820 ( .A1(DATAIN[7]), .A2(n147), .ZN(n1747) );
  AND2_X1 U1821 ( .A1(DATAIN[7]), .A2(RST), .ZN(n1748) );
  AND2_X1 U1822 ( .A1(DATAIN[7]), .A2(n150), .ZN(n1749) );
  AND2_X1 U1823 ( .A1(DATAIN[7]), .A2(n146), .ZN(n1750) );
  AND2_X1 U1824 ( .A1(DATAIN[7]), .A2(n147), .ZN(n1751) );
  AND2_X1 U1825 ( .A1(DATAIN[7]), .A2(n145), .ZN(n1752) );
  AND2_X1 U1826 ( .A1(DATAIN[7]), .A2(n144), .ZN(n1753) );
  AND2_X1 U1827 ( .A1(DATAIN[7]), .A2(RST), .ZN(n1754) );
  AND2_X1 U1828 ( .A1(DATAIN[7]), .A2(n142), .ZN(n1755) );
  AND2_X1 U1829 ( .A1(DATAIN[7]), .A2(n140), .ZN(n1756) );
  AND2_X1 U1830 ( .A1(DATAIN[7]), .A2(n141), .ZN(n1757) );
  AND2_X1 U1831 ( .A1(DATAIN[7]), .A2(n141), .ZN(n1758) );
  AND2_X1 U1832 ( .A1(DATAIN[7]), .A2(n137), .ZN(n1759) );
  AND2_X1 U1833 ( .A1(DATAIN[7]), .A2(n139), .ZN(n1760) );
  AND2_X1 U1834 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1761) );
  AND2_X1 U1835 ( .A1(DATAIN[0]), .A2(n148), .ZN(n1762) );
  AND2_X1 U1836 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1763) );
  AND2_X1 U1837 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1764) );
  AND2_X1 U1838 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1765) );
  AND2_X1 U1839 ( .A1(DATAIN[0]), .A2(n145), .ZN(n1766) );
  AND2_X1 U1840 ( .A1(DATAIN[0]), .A2(n144), .ZN(n1767) );
  AND2_X1 U1841 ( .A1(DATAIN[0]), .A2(n143), .ZN(n1768) );
  AND2_X1 U1842 ( .A1(DATAIN[0]), .A2(n145), .ZN(n1769) );
  AND2_X1 U1843 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1770) );
  AND2_X1 U1844 ( .A1(DATAIN[0]), .A2(n141), .ZN(n1771) );
  AND2_X1 U1845 ( .A1(DATAIN[0]), .A2(n149), .ZN(n1772) );
  AND2_X1 U1846 ( .A1(DATAIN[0]), .A2(n148), .ZN(n1773) );
  AND2_X1 U1847 ( .A1(DATAIN[0]), .A2(n140), .ZN(n1774) );
  AND2_X1 U1848 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1775) );
  AND2_X1 U1849 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1776) );
  BUF_X2 U1850 ( .A(n78), .Z(n1777) );
  BUF_X2 U1851 ( .A(n134), .Z(n1778) );
  BUF_X2 U1852 ( .A(n82), .Z(n1779) );
  BUF_X2 U1853 ( .A(n88), .Z(n1780) );
  BUF_X2 U1854 ( .A(n94), .Z(n1781) );
  AND2_X1 U1855 ( .A1(DATAIN[30]), .A2(RST), .ZN(n1782) );
  AND2_X1 U1856 ( .A1(n1638), .A2(RST), .ZN(n1783) );
  AND2_X1 U1857 ( .A1(DATAIN[23]), .A2(n141), .ZN(n1784) );
  AND2_X1 U1858 ( .A1(n1640), .A2(RST), .ZN(n1785) );
  AND2_X1 U1859 ( .A1(n1641), .A2(n137), .ZN(n1786) );
  AND2_X1 U1860 ( .A1(n1642), .A2(n140), .ZN(n1787) );
  AND2_X1 U1861 ( .A1(n1643), .A2(RST), .ZN(n1788) );
  BUF_X2 U1862 ( .A(DATAIN[8]), .Z(n1789) );
  BUF_X2 U1863 ( .A(DATAIN[9]), .Z(n1790) );
  BUF_X2 U1864 ( .A(DATAIN[18]), .Z(n1791) );
  BUF_X2 U1865 ( .A(DATAIN[26]), .Z(n1792) );
  BUF_X2 U1866 ( .A(DATAIN[22]), .Z(n1793) );
  BUF_X2 U1867 ( .A(DATAIN[12]), .Z(n1794) );
  NOR2_X2 U1868 ( .A1(n1797), .A2(n1796), .ZN(n1795) );
  NAND2_X2 U1869 ( .A1(n897), .A2(WR), .ZN(n1796) );
  INV_X2 U1870 ( .A(n894), .ZN(n1797) );
  NAND2_X1 U1871 ( .A1(EN), .A2(n1798), .ZN(n156) );
  NOR2_X2 U1872 ( .A1(n1800), .A2(n1799), .ZN(n1798) );
  NAND2_X2 U1873 ( .A1(ADD_WR[4]), .A2(WR), .ZN(n1799) );
  INV_X2 U1874 ( .A(n897), .ZN(n1800) );
  NAND2_X1 U1875 ( .A1(EN), .A2(n1801), .ZN(n157) );
  NOR2_X2 U1876 ( .A1(n1803), .A2(n1802), .ZN(n1801) );
  NAND2_X2 U1877 ( .A1(ADD_WR[3]), .A2(WR), .ZN(n1802) );
  INV_X2 U1878 ( .A(n894), .ZN(n1803) );
  INV_X2 U1879 ( .A(n76), .ZN(n75) );
  INV_X2 U1880 ( .A(n88), .ZN(n87) );
  INV_X2 U1881 ( .A(n94), .ZN(n93) );
  INV_X2 U1882 ( .A(n134), .ZN(n133) );
  INV_X2 U1883 ( .A(n78), .ZN(n77) );
  INV_X2 U1884 ( .A(n82), .ZN(n81) );
  INV_X2 U1885 ( .A(n110), .ZN(n109) );
  INV_X2 U1886 ( .A(n114), .ZN(n113) );
  INV_X2 U1887 ( .A(n98), .ZN(n97) );
  INV_X2 U1888 ( .A(n102), .ZN(n101) );
  INV_X2 U1889 ( .A(n104), .ZN(n103) );
  INV_X2 U1890 ( .A(n118), .ZN(n117) );
  INV_X2 U1891 ( .A(n84), .ZN(n83) );
  INV_X2 U1892 ( .A(n92), .ZN(n91) );
  INV_X2 U1893 ( .A(n100), .ZN(n99) );
  INV_X2 U1894 ( .A(n112), .ZN(n111) );
  INV_X2 U1895 ( .A(n128), .ZN(n127) );
  NAND2_X1 U1896 ( .A1(EN), .A2(n1804), .ZN(n1629) );
  INV_X2 U1897 ( .A(n1805), .ZN(n1804) );
  NAND3_X1 U1898 ( .A1(ADD_WR[4]), .A2(ADD_WR[3]), .A3(WR), .ZN(n1805) );
  CLKBUF_X1 U1899 ( .A(EN), .Z(n1806) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n1808), .CK(net7260), .Q(
        \REGISTERS[31][28] ) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n1807), .CK(net7260), .Q(
        \REGISTERS[31][31] ) );
  INV_X2 U45 ( .A(n136), .ZN(n135) );
  AND2_X1 U1900 ( .A1(DATAIN[31]), .A2(n153), .ZN(n1807) );
  AND2_X1 U1901 ( .A1(DATAIN[28]), .A2(RST), .ZN(n1808) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n1810), .CK(net7170), .Q(
        \REGISTERS[13][11] ) );
  AND2_X1 U1903 ( .A1(DATAIN[11]), .A2(n146), .ZN(n1810) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n1811), .CK(net7165), .Q(
        \REGISTERS[12][16] ) );
  AND2_X1 U1904 ( .A1(DATAIN[16]), .A2(n154), .ZN(n1811) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n2694), .CK(net7170), .Q(
        \REGISTERS[13][4] ) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n2693), .CK(net7165), .Q(
        \REGISTERS[12][4] ) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n2692), .CK(net7160), .Q(
        \REGISTERS[11][4] ) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n2691), .CK(net7155), .Q(
        \REGISTERS[10][4] ) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n2690), .CK(net7150), .Q(\REGISTERS[9][4] ) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n2689), .CK(net7145), .Q(\REGISTERS[8][4] ) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n2688), .CK(net7205), .Q(
        \REGISTERS[20][30] ) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n2687), .CK(net7185), .Q(
        \REGISTERS[16][30] ) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n2686), .CK(net7175), .Q(
        \REGISTERS[14][30] ) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n2685), .CK(net7170), .Q(
        \REGISTERS[13][30] ) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n2684), .CK(net7165), .Q(
        \REGISTERS[12][30] ) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n2683), .CK(net7160), .Q(
        \REGISTERS[11][30] ) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n2682), .CK(net7155), .Q(
        \REGISTERS[10][30] ) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n2681), .CK(net7150), .Q(
        \REGISTERS[9][30] ) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n2680), .CK(net7145), .Q(
        \REGISTERS[8][30] ) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n2679), .CK(net7205), .Q(
        \REGISTERS[20][23] ) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n2678), .CK(net7185), .Q(
        \REGISTERS[16][23] ) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n2677), .CK(net7175), .Q(
        \REGISTERS[14][23] ) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n2676), .CK(net7170), .Q(
        \REGISTERS[13][23] ) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n2675), .CK(net7165), .Q(
        \REGISTERS[12][23] ) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n2674), .CK(net7160), .Q(
        \REGISTERS[11][23] ) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n2673), .CK(net7155), .Q(
        \REGISTERS[10][23] ) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n2672), .CK(net7150), .Q(
        \REGISTERS[9][23] ) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n2671), .CK(net7145), .Q(
        \REGISTERS[8][23] ) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n2670), .CK(net7205), .Q(
        \REGISTERS[20][29] ) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n2669), .CK(net7185), .Q(
        \REGISTERS[16][29] ) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n2668), .CK(net7175), .Q(
        \REGISTERS[14][29] ) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n2667), .CK(net7170), .Q(
        \REGISTERS[13][29] ) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n2666), .CK(net7165), .Q(
        \REGISTERS[12][29] ) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n2665), .CK(net7160), .Q(
        \REGISTERS[11][29] ) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n2664), .CK(net7155), .Q(
        \REGISTERS[10][29] ) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n2663), .CK(net7150), .Q(
        \REGISTERS[9][29] ) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n2662), .CK(net7145), .Q(
        \REGISTERS[8][29] ) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n2661), .CK(net7205), .Q(
        \REGISTERS[20][27] ) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n2660), .CK(net7185), .Q(
        \REGISTERS[16][27] ) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n2659), .CK(net7175), .Q(
        \REGISTERS[14][27] ) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n2658), .CK(net7170), .Q(
        \REGISTERS[13][27] ) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n2657), .CK(net7165), .Q(
        \REGISTERS[12][27] ) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n2656), .CK(net7160), .Q(
        \REGISTERS[11][27] ) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n2655), .CK(net7155), .Q(
        \REGISTERS[10][27] ) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n2654), .CK(net7150), .Q(
        \REGISTERS[9][27] ) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n2653), .CK(net7145), .Q(
        \REGISTERS[8][27] ) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n2652), .CK(net7230), .Q(
        \REGISTERS[25][5] ) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n2651), .CK(net7205), .Q(
        \REGISTERS[20][5] ) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n2650), .CK(net7185), .Q(
        \REGISTERS[16][5] ) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n2649), .CK(net7175), .Q(
        \REGISTERS[14][5] ) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n2648), .CK(net7170), .Q(
        \REGISTERS[13][5] ) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n2647), .CK(net7165), .Q(
        \REGISTERS[12][5] ) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n2646), .CK(net7160), .Q(
        \REGISTERS[11][5] ) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n2645), .CK(net7155), .Q(
        \REGISTERS[10][5] ) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n2644), .CK(net7150), .Q(\REGISTERS[9][5] ) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n2643), .CK(net7145), .Q(\REGISTERS[8][5] ) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n2642), .CK(net7205), .Q(
        \REGISTERS[20][21] ) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n2641), .CK(net7185), .Q(
        \REGISTERS[16][21] ) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n2640), .CK(net7175), .Q(
        \REGISTERS[14][21] ) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n2639), .CK(net7170), .Q(
        \REGISTERS[13][21] ) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n2638), .CK(net7165), .Q(
        \REGISTERS[12][21] ) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n2637), .CK(net7160), .Q(
        \REGISTERS[11][21] ) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n2636), .CK(net7155), .Q(
        \REGISTERS[10][21] ) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n2635), .CK(net7150), .Q(
        \REGISTERS[9][21] ) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n2634), .CK(net7145), .Q(
        \REGISTERS[8][21] ) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n2633), .CK(net7205), .Q(
        \REGISTERS[20][24] ) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n2632), .CK(net7185), .Q(
        \REGISTERS[16][24] ) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n2631), .CK(net7175), .Q(
        \REGISTERS[14][24] ) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n2630), .CK(net7170), .Q(
        \REGISTERS[13][24] ) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n2629), .CK(net7165), .Q(
        \REGISTERS[12][24] ) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n2628), .CK(net7160), .Q(
        \REGISTERS[11][24] ) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n2627), .CK(net7155), .Q(
        \REGISTERS[10][24] ) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n2626), .CK(net7150), .Q(
        \REGISTERS[9][24] ) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n2625), .CK(net7145), .Q(
        \REGISTERS[8][24] ) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n2624), .CK(net7205), .Q(
        \REGISTERS[20][17] ) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n2623), .CK(net7195), .Q(
        \REGISTERS[18][17] ) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n2622), .CK(net7185), .Q(
        \REGISTERS[16][17] ) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n2621), .CK(net7175), .Q(
        \REGISTERS[14][17] ) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n2620), .CK(net7170), .Q(
        \REGISTERS[13][17] ) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n2619), .CK(net7165), .Q(
        \REGISTERS[12][17] ) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n2618), .CK(net7160), .Q(
        \REGISTERS[11][17] ) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n2617), .CK(net7155), .Q(
        \REGISTERS[10][17] ) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n2616), .CK(net7150), .Q(
        \REGISTERS[9][17] ) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n2615), .CK(net7145), .Q(
        \REGISTERS[8][17] ) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n2614), .CK(net7205), .Q(
        \REGISTERS[20][8] ) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n2613), .CK(net7195), .Q(
        \REGISTERS[18][8] ) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n2612), .CK(net7185), .Q(
        \REGISTERS[16][8] ) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n2611), .CK(net7175), .Q(
        \REGISTERS[14][8] ) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n2610), .CK(net7170), .Q(
        \REGISTERS[13][8] ) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n2609), .CK(net7165), .Q(
        \REGISTERS[12][8] ) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n2608), .CK(net7160), .Q(
        \REGISTERS[11][8] ) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n2607), .CK(net7155), .Q(
        \REGISTERS[10][8] ) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n2606), .CK(net7150), .Q(\REGISTERS[9][8] ) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n2605), .CK(net7145), .Q(\REGISTERS[8][8] ) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n2604), .CK(net7205), .Q(
        \REGISTERS[20][22] ) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n2603), .CK(net7195), .Q(
        \REGISTERS[18][22] ) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n2602), .CK(net7185), .Q(
        \REGISTERS[16][22] ) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n2601), .CK(net7175), .Q(
        \REGISTERS[14][22] ) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n2600), .CK(net7170), .Q(
        \REGISTERS[13][22] ) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n2599), .CK(net7165), .Q(
        \REGISTERS[12][22] ) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n2598), .CK(net7160), .Q(
        \REGISTERS[11][22] ) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n2597), .CK(net7155), .Q(
        \REGISTERS[10][22] ) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n2596), .CK(net7150), .Q(
        \REGISTERS[9][22] ) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n2595), .CK(net7145), .Q(
        \REGISTERS[8][22] ) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n2594), .CK(net7205), .Q(
        \REGISTERS[20][18] ) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n2593), .CK(net7195), .Q(
        \REGISTERS[18][18] ) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n2592), .CK(net7185), .Q(
        \REGISTERS[16][18] ) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n2591), .CK(net7175), .Q(
        \REGISTERS[14][18] ) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n2590), .CK(net7170), .Q(
        \REGISTERS[13][18] ) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n2589), .CK(net7165), .Q(
        \REGISTERS[12][18] ) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n2588), .CK(net7160), .Q(
        \REGISTERS[11][18] ) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n2587), .CK(net7155), .Q(
        \REGISTERS[10][18] ) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n2586), .CK(net7150), .Q(
        \REGISTERS[9][18] ) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n2585), .CK(net7145), .Q(
        \REGISTERS[8][18] ) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n2584), .CK(net7205), .Q(
        \REGISTERS[20][14] ) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n2583), .CK(net7195), .Q(
        \REGISTERS[18][14] ) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n2582), .CK(net7185), .Q(
        \REGISTERS[16][14] ) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n2581), .CK(net7175), .Q(
        \REGISTERS[14][14] ) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n2580), .CK(net7170), .Q(
        \REGISTERS[13][14] ) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n2579), .CK(net7165), .Q(
        \REGISTERS[12][14] ) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n2578), .CK(net7160), .Q(
        \REGISTERS[11][14] ) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n2577), .CK(net7155), .Q(
        \REGISTERS[10][14] ) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n2576), .CK(net7150), .Q(
        \REGISTERS[9][14] ) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n2575), .CK(net7145), .Q(
        \REGISTERS[8][14] ) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n2574), .CK(net7205), .Q(
        \REGISTERS[20][10] ) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n2573), .CK(net7195), .Q(
        \REGISTERS[18][10] ) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n2572), .CK(net7185), .Q(
        \REGISTERS[16][10] ) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n2571), .CK(net7175), .Q(
        \REGISTERS[14][10] ) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n2570), .CK(net7170), .Q(
        \REGISTERS[13][10] ) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n2569), .CK(net7165), .Q(
        \REGISTERS[12][10] ) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n2568), .CK(net7160), .Q(
        \REGISTERS[11][10] ) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n2567), .CK(net7155), .Q(
        \REGISTERS[10][10] ) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n2566), .CK(net7150), .Q(
        \REGISTERS[9][10] ) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n2565), .CK(net7145), .Q(
        \REGISTERS[8][10] ) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n2564), .CK(net7205), .Q(
        \REGISTERS[20][9] ) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n2563), .CK(net7195), .Q(
        \REGISTERS[18][9] ) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n2562), .CK(net7185), .Q(
        \REGISTERS[16][9] ) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n2561), .CK(net7175), .Q(
        \REGISTERS[14][9] ) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n2560), .CK(net7170), .Q(
        \REGISTERS[13][9] ) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n2559), .CK(net7165), .Q(
        \REGISTERS[12][9] ) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n2558), .CK(net7160), .Q(
        \REGISTERS[11][9] ) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n2557), .CK(net7155), .Q(
        \REGISTERS[10][9] ) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n2556), .CK(net7150), .Q(\REGISTERS[9][9] ) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n2555), .CK(net7145), .Q(\REGISTERS[8][9] ) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n2554), .CK(net7205), .Q(
        \REGISTERS[20][3] ) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n2553), .CK(net7195), .Q(
        \REGISTERS[18][3] ) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n2552), .CK(net7185), .Q(
        \REGISTERS[16][3] ) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n2551), .CK(net7175), .Q(
        \REGISTERS[14][3] ) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n2550), .CK(net7170), .Q(
        \REGISTERS[13][3] ) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n2549), .CK(net7165), .Q(
        \REGISTERS[12][3] ) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n2548), .CK(net7160), .Q(
        \REGISTERS[11][3] ) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n2547), .CK(net7155), .Q(
        \REGISTERS[10][3] ) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n2546), .CK(net7150), .Q(\REGISTERS[9][3] ) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n2545), .CK(net7145), .Q(\REGISTERS[8][3] ) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n2544), .CK(net7205), .Q(
        \REGISTERS[20][12] ) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n2543), .CK(net7195), .Q(
        \REGISTERS[18][12] ) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n2542), .CK(net7185), .Q(
        \REGISTERS[16][12] ) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n2541), .CK(net7175), .Q(
        \REGISTERS[14][12] ) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n2540), .CK(net7170), .Q(
        \REGISTERS[13][12] ) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n2539), .CK(net7165), .Q(
        \REGISTERS[12][12] ) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n2538), .CK(net7160), .Q(
        \REGISTERS[11][12] ) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n2537), .CK(net7155), .Q(
        \REGISTERS[10][12] ) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n2536), .CK(net7150), .Q(
        \REGISTERS[9][12] ) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n2535), .CK(net7145), .Q(
        \REGISTERS[8][12] ) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n2534), .CK(net7205), .Q(
        \REGISTERS[20][26] ) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n2533), .CK(net7195), .Q(
        \REGISTERS[18][26] ) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n2532), .CK(net7185), .Q(
        \REGISTERS[16][26] ) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n2531), .CK(net7175), .Q(
        \REGISTERS[14][26] ) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n2530), .CK(net7170), .Q(
        \REGISTERS[13][26] ) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n2529), .CK(net7165), .Q(
        \REGISTERS[12][26] ) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n2528), .CK(net7160), .Q(
        \REGISTERS[11][26] ) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n2527), .CK(net7155), .Q(
        \REGISTERS[10][26] ) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n2526), .CK(net7150), .Q(
        \REGISTERS[9][26] ) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n2525), .CK(net7145), .Q(
        \REGISTERS[8][26] ) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n2524), .CK(net7205), .Q(
        \REGISTERS[20][19] ) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n2523), .CK(net7195), .Q(
        \REGISTERS[18][19] ) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n2522), .CK(net7185), .Q(
        \REGISTERS[16][19] ) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n2521), .CK(net7175), .Q(
        \REGISTERS[14][19] ) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n2520), .CK(net7170), .Q(
        \REGISTERS[13][19] ) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n2519), .CK(net7165), .Q(
        \REGISTERS[12][19] ) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n2518), .CK(net7160), .Q(
        \REGISTERS[11][19] ) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n2517), .CK(net7155), .Q(
        \REGISTERS[10][19] ) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n2516), .CK(net7150), .Q(
        \REGISTERS[9][19] ) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n2515), .CK(net7145), .Q(
        \REGISTERS[8][19] ) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n2514), .CK(net7160), .Q(
        \REGISTERS[11][16] ) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n2513), .CK(net7155), .Q(
        \REGISTERS[10][16] ) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n2512), .CK(net7150), .Q(
        \REGISTERS[9][16] ) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n2511), .CK(net7145), .Q(
        \REGISTERS[8][16] ) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n2510), .CK(net7165), .Q(
        \REGISTERS[12][13] ) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n2509), .CK(net7160), .Q(
        \REGISTERS[11][13] ) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n2508), .CK(net7155), .Q(
        \REGISTERS[10][13] ) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n2507), .CK(net7150), .Q(
        \REGISTERS[9][13] ) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n2506), .CK(net7145), .Q(
        \REGISTERS[8][13] ) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n2505), .CK(net7165), .Q(
        \REGISTERS[12][11] ) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n2504), .CK(net7160), .Q(
        \REGISTERS[11][11] ) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n2503), .CK(net7155), .Q(
        \REGISTERS[10][11] ) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n2502), .CK(net7150), .Q(
        \REGISTERS[9][11] ) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n2501), .CK(net7145), .Q(
        \REGISTERS[8][11] ) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n2500), .CK(net7205), .Q(
        \REGISTERS[20][1] ) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n2499), .CK(net7185), .Q(
        \REGISTERS[16][1] ) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n2498), .CK(net7175), .Q(
        \REGISTERS[14][1] ) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n2497), .CK(net7170), .Q(
        \REGISTERS[13][1] ) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n2496), .CK(net7165), .Q(
        \REGISTERS[12][1] ) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n2495), .CK(net7160), .Q(
        \REGISTERS[11][1] ) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n2494), .CK(net7155), .Q(
        \REGISTERS[10][1] ) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n2493), .CK(net7150), .Q(\REGISTERS[9][1] ) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n2492), .CK(net7145), .Q(\REGISTERS[8][1] ) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n2491), .CK(net7104), .Q(
        \REGISTERS[0][18] ) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n2490), .CK(net7260), .Q(
        \REGISTERS[31][11] ) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n2489), .CK(net7255), .Q(
        \REGISTERS[30][11] ) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n2488), .CK(net7250), .Q(
        \REGISTERS[29][11] ) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n2487), .CK(net7245), .Q(
        \REGISTERS[28][11] ) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n2486), .CK(net7240), .Q(
        \REGISTERS[27][11] ) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n2485), .CK(net7235), .Q(
        \REGISTERS[26][11] ) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n2484), .CK(net7230), .Q(
        \REGISTERS[25][11] ) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n2483), .CK(net7225), .Q(
        \REGISTERS[24][11] ) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n2482), .CK(net7220), .Q(
        \REGISTERS[23][11] ) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n2481), .CK(net7215), .Q(
        \REGISTERS[22][11] ) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n2480), .CK(net7210), .Q(
        \REGISTERS[21][11] ) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n2479), .CK(net7200), .Q(
        \REGISTERS[19][11] ) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n2478), .CK(net7190), .Q(
        \REGISTERS[17][11] ) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n2477), .CK(net7180), .Q(
        \REGISTERS[15][11] ) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n2476), .CK(net7140), .Q(
        \REGISTERS[7][11] ) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n2475), .CK(net7135), .Q(
        \REGISTERS[6][11] ) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n2474), .CK(net7130), .Q(
        \REGISTERS[5][11] ) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n2473), .CK(net7125), .Q(
        \REGISTERS[4][11] ) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n2472), .CK(net7120), .Q(
        \REGISTERS[3][11] ) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n2471), .CK(net7115), .Q(
        \REGISTERS[2][11] ) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n2470), .CK(net7110), .Q(
        \REGISTERS[1][11] ) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n2469), .CK(net7104), .Q(
        \REGISTERS[0][11] ) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n2468), .CK(net7260), .Q(
        \REGISTERS[31][16] ) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n2467), .CK(net7255), .Q(
        \REGISTERS[30][16] ) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n2466), .CK(net7250), .Q(
        \REGISTERS[29][16] ) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n2465), .CK(net7245), .Q(
        \REGISTERS[28][16] ) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n2464), .CK(net7240), .Q(
        \REGISTERS[27][16] ) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n2463), .CK(net7235), .Q(
        \REGISTERS[26][16] ) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n2462), .CK(net7230), .Q(
        \REGISTERS[25][16] ) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n2461), .CK(net7225), .Q(
        \REGISTERS[24][16] ) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n2460), .CK(net7220), .Q(
        \REGISTERS[23][16] ) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n2459), .CK(net7215), .Q(
        \REGISTERS[22][16] ) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n2458), .CK(net7210), .Q(
        \REGISTERS[21][16] ) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n2457), .CK(net7200), .Q(
        \REGISTERS[19][16] ) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n2456), .CK(net7190), .Q(
        \REGISTERS[17][16] ) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n2455), .CK(net7180), .Q(
        \REGISTERS[15][16] ) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n2454), .CK(net7140), .Q(
        \REGISTERS[7][16] ) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n2453), .CK(net7135), .Q(
        \REGISTERS[6][16] ) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n2452), .CK(net7130), .Q(
        \REGISTERS[5][16] ) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n2451), .CK(net7125), .Q(
        \REGISTERS[4][16] ) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n2450), .CK(net7120), .Q(
        \REGISTERS[3][16] ) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n2449), .CK(net7115), .Q(
        \REGISTERS[2][16] ) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n2448), .CK(net7110), .Q(
        \REGISTERS[1][16] ) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n2447), .CK(net7104), .Q(
        \REGISTERS[0][16] ) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n2446), .CK(net7260), .Q(
        \REGISTERS[31][27] ) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n2445), .CK(net7255), .Q(
        \REGISTERS[30][27] ) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n2444), .CK(net7250), .Q(
        \REGISTERS[29][27] ) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n2443), .CK(net7245), .Q(
        \REGISTERS[28][27] ) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n2442), .CK(net7240), .Q(
        \REGISTERS[27][27] ) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n2441), .CK(net7235), .Q(
        \REGISTERS[26][27] ) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n2440), .CK(net7230), .Q(
        \REGISTERS[25][27] ) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n2439), .CK(net7225), .Q(
        \REGISTERS[24][27] ) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n2438), .CK(net7220), .Q(
        \REGISTERS[23][27] ) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n2437), .CK(net7215), .Q(
        \REGISTERS[22][27] ) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n2436), .CK(net7210), .Q(
        \REGISTERS[21][27] ) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n2435), .CK(net7200), .Q(
        \REGISTERS[19][27] ) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n2434), .CK(net7190), .Q(
        \REGISTERS[17][27] ) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n2433), .CK(net7180), .Q(
        \REGISTERS[15][27] ) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n2432), .CK(net7140), .Q(
        \REGISTERS[7][27] ) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n2431), .CK(net7135), .Q(
        \REGISTERS[6][27] ) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n2430), .CK(net7130), .Q(
        \REGISTERS[5][27] ) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n2429), .CK(net7125), .Q(
        \REGISTERS[4][27] ) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n2428), .CK(net7120), .Q(
        \REGISTERS[3][27] ) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n2427), .CK(net7115), .Q(
        \REGISTERS[2][27] ) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n2426), .CK(net7110), .Q(
        \REGISTERS[1][27] ) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n2425), .CK(net7104), .Q(
        \REGISTERS[0][27] ) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n2424), .CK(net7260), .Q(
        \REGISTERS[31][21] ) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n2423), .CK(net7255), .Q(
        \REGISTERS[30][21] ) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n2422), .CK(net7250), .Q(
        \REGISTERS[29][21] ) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n2421), .CK(net7245), .Q(
        \REGISTERS[28][21] ) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n2420), .CK(net7240), .Q(
        \REGISTERS[27][21] ) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n2419), .CK(net7235), .Q(
        \REGISTERS[26][21] ) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n2418), .CK(net7230), .Q(
        \REGISTERS[25][21] ) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n2417), .CK(net7225), .Q(
        \REGISTERS[24][21] ) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n2416), .CK(net7220), .Q(
        \REGISTERS[23][21] ) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n2415), .CK(net7215), .Q(
        \REGISTERS[22][21] ) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n2414), .CK(net7210), .Q(
        \REGISTERS[21][21] ) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n2413), .CK(net7200), .Q(
        \REGISTERS[19][21] ) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n2412), .CK(net7190), .Q(
        \REGISTERS[17][21] ) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n2411), .CK(net7180), .Q(
        \REGISTERS[15][21] ) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n2410), .CK(net7140), .Q(
        \REGISTERS[7][21] ) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n2409), .CK(net7135), .Q(
        \REGISTERS[6][21] ) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n2408), .CK(net7130), .Q(
        \REGISTERS[5][21] ) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n2407), .CK(net7125), .Q(
        \REGISTERS[4][21] ) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n2406), .CK(net7120), .Q(
        \REGISTERS[3][21] ) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n2405), .CK(net7115), .Q(
        \REGISTERS[2][21] ) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n2404), .CK(net7110), .Q(
        \REGISTERS[1][21] ) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n2403), .CK(net7104), .Q(
        \REGISTERS[0][21] ) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n2402), .CK(net7260), .Q(
        \REGISTERS[31][24] ) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n2401), .CK(net7255), .Q(
        \REGISTERS[30][24] ) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n2400), .CK(net7250), .Q(
        \REGISTERS[29][24] ) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n2399), .CK(net7245), .Q(
        \REGISTERS[28][24] ) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n2398), .CK(net7240), .Q(
        \REGISTERS[27][24] ) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n2397), .CK(net7235), .Q(
        \REGISTERS[26][24] ) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n2396), .CK(net7230), .Q(
        \REGISTERS[25][24] ) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n2395), .CK(net7225), .Q(
        \REGISTERS[24][24] ) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n2394), .CK(net7220), .Q(
        \REGISTERS[23][24] ) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n2393), .CK(net7215), .Q(
        \REGISTERS[22][24] ) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n2392), .CK(net7210), .Q(
        \REGISTERS[21][24] ) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n2391), .CK(net7200), .Q(
        \REGISTERS[19][24] ) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n2390), .CK(net7190), .Q(
        \REGISTERS[17][24] ) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n2389), .CK(net7180), .Q(
        \REGISTERS[15][24] ) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n2388), .CK(net7140), .Q(
        \REGISTERS[7][24] ) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n2387), .CK(net7135), .Q(
        \REGISTERS[6][24] ) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n2386), .CK(net7130), .Q(
        \REGISTERS[5][24] ) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n2385), .CK(net7125), .Q(
        \REGISTERS[4][24] ) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n2384), .CK(net7120), .Q(
        \REGISTERS[3][24] ) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n2383), .CK(net7115), .Q(
        \REGISTERS[2][24] ) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n2382), .CK(net7110), .Q(
        \REGISTERS[1][24] ) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n2381), .CK(net7104), .Q(
        \REGISTERS[0][24] ) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n2380), .CK(net7260), .Q(
        \REGISTERS[31][13] ) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n2379), .CK(net7255), .Q(
        \REGISTERS[30][13] ) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n2378), .CK(net7250), .Q(
        \REGISTERS[29][13] ) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n2377), .CK(net7245), .Q(
        \REGISTERS[28][13] ) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n2376), .CK(net7240), .Q(
        \REGISTERS[27][13] ) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n2375), .CK(net7235), .Q(
        \REGISTERS[26][13] ) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n2374), .CK(net7230), .Q(
        \REGISTERS[25][13] ) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n2373), .CK(net7225), .Q(
        \REGISTERS[24][13] ) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n2372), .CK(net7220), .Q(
        \REGISTERS[23][13] ) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n2371), .CK(net7215), .Q(
        \REGISTERS[22][13] ) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n2370), .CK(net7210), .Q(
        \REGISTERS[21][13] ) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n2369), .CK(net7200), .Q(
        \REGISTERS[19][13] ) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n2368), .CK(net7190), .Q(
        \REGISTERS[17][13] ) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n2367), .CK(net7180), .Q(
        \REGISTERS[15][13] ) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n2366), .CK(net7140), .Q(
        \REGISTERS[7][13] ) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n2365), .CK(net7135), .Q(
        \REGISTERS[6][13] ) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n2364), .CK(net7130), .Q(
        \REGISTERS[5][13] ) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n2363), .CK(net7125), .Q(
        \REGISTERS[4][13] ) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n2362), .CK(net7120), .Q(
        \REGISTERS[3][13] ) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n2361), .CK(net7115), .Q(
        \REGISTERS[2][13] ) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n2360), .CK(net7110), .Q(
        \REGISTERS[1][13] ) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n2359), .CK(net7104), .Q(
        \REGISTERS[0][13] ) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n2358), .CK(net7260), .Q(
        \REGISTERS[31][5] ) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n2357), .CK(net7255), .Q(
        \REGISTERS[30][5] ) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n2356), .CK(net7250), .Q(
        \REGISTERS[29][5] ) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n2355), .CK(net7245), .Q(
        \REGISTERS[28][5] ) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n2354), .CK(net7240), .Q(
        \REGISTERS[27][5] ) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n2353), .CK(net7235), .Q(
        \REGISTERS[26][5] ) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n2352), .CK(net7225), .Q(
        \REGISTERS[24][5] ) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n2351), .CK(net7220), .Q(
        \REGISTERS[23][5] ) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n2350), .CK(net7215), .Q(
        \REGISTERS[22][5] ) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n2349), .CK(net7210), .Q(
        \REGISTERS[21][5] ) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n2348), .CK(net7200), .Q(
        \REGISTERS[19][5] ) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n2347), .CK(net7195), .Q(
        \REGISTERS[18][5] ) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n2346), .CK(net7190), .Q(
        \REGISTERS[17][5] ) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n2345), .CK(net7180), .Q(
        \REGISTERS[15][5] ) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n2344), .CK(net7140), .Q(\REGISTERS[7][5] ) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n2343), .CK(net7135), .Q(\REGISTERS[6][5] ) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n2342), .CK(net7130), .Q(\REGISTERS[5][5] ) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n2341), .CK(net7125), .Q(\REGISTERS[4][5] ) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n2340), .CK(net7120), .Q(\REGISTERS[3][5] ) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n2339), .CK(net7115), .Q(\REGISTERS[2][5] ) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n2338), .CK(net7110), .Q(\REGISTERS[1][5] ) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n2337), .CK(net7104), .Q(\REGISTERS[0][5] ) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n2336), .CK(net7260), .Q(
        \REGISTERS[31][29] ) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n2335), .CK(net7255), .Q(
        \REGISTERS[30][29] ) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n2334), .CK(net7250), .Q(
        \REGISTERS[29][29] ) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n2333), .CK(net7245), .Q(
        \REGISTERS[28][29] ) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n2332), .CK(net7240), .Q(
        \REGISTERS[27][29] ) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n2331), .CK(net7235), .Q(
        \REGISTERS[26][29] ) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n2330), .CK(net7230), .Q(
        \REGISTERS[25][29] ) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n2329), .CK(net7225), .Q(
        \REGISTERS[24][29] ) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n2328), .CK(net7220), .Q(
        \REGISTERS[23][29] ) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n2327), .CK(net7215), .Q(
        \REGISTERS[22][29] ) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n2326), .CK(net7210), .Q(
        \REGISTERS[21][29] ) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n2325), .CK(net7200), .Q(
        \REGISTERS[19][29] ) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n2324), .CK(net7190), .Q(
        \REGISTERS[17][29] ) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n2323), .CK(net7180), .Q(
        \REGISTERS[15][29] ) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n2322), .CK(net7140), .Q(
        \REGISTERS[7][29] ) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n2321), .CK(net7135), .Q(
        \REGISTERS[6][29] ) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n2320), .CK(net7130), .Q(
        \REGISTERS[5][29] ) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n2319), .CK(net7125), .Q(
        \REGISTERS[4][29] ) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n2318), .CK(net7120), .Q(
        \REGISTERS[3][29] ) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n2317), .CK(net7115), .Q(
        \REGISTERS[2][29] ) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n2316), .CK(net7110), .Q(
        \REGISTERS[1][29] ) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n2315), .CK(net7104), .Q(
        \REGISTERS[0][29] ) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n2314), .CK(net7255), .Q(
        \REGISTERS[30][14] ) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n2313), .CK(net7250), .Q(
        \REGISTERS[29][14] ) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n2312), .CK(net7245), .Q(
        \REGISTERS[28][14] ) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n2311), .CK(net7240), .Q(
        \REGISTERS[27][14] ) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n2310), .CK(net7235), .Q(
        \REGISTERS[26][14] ) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n2309), .CK(net7230), .Q(
        \REGISTERS[25][14] ) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n2308), .CK(net7225), .Q(
        \REGISTERS[24][14] ) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n2307), .CK(net7220), .Q(
        \REGISTERS[23][14] ) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n2306), .CK(net7215), .Q(
        \REGISTERS[22][14] ) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n2305), .CK(net7210), .Q(
        \REGISTERS[21][14] ) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n2304), .CK(net7260), .Q(
        \REGISTERS[31][17] ) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n2303), .CK(net7255), .Q(
        \REGISTERS[30][17] ) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n2302), .CK(net7250), .Q(
        \REGISTERS[29][17] ) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n2301), .CK(net7245), .Q(
        \REGISTERS[28][17] ) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n2300), .CK(net7240), .Q(
        \REGISTERS[27][17] ) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n2299), .CK(net7235), .Q(
        \REGISTERS[26][17] ) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n2298), .CK(net7230), .Q(
        \REGISTERS[25][17] ) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n2297), .CK(net7225), .Q(
        \REGISTERS[24][17] ) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n2296), .CK(net7220), .Q(
        \REGISTERS[23][17] ) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n2295), .CK(net7215), .Q(
        \REGISTERS[22][17] ) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n2294), .CK(net7210), .Q(
        \REGISTERS[21][17] ) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n2293), .CK(net7200), .Q(
        \REGISTERS[19][17] ) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n2292), .CK(net7190), .Q(
        \REGISTERS[17][17] ) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n2291), .CK(net7180), .Q(
        \REGISTERS[15][17] ) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n2290), .CK(net7140), .Q(
        \REGISTERS[7][17] ) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n2289), .CK(net7135), .Q(
        \REGISTERS[6][17] ) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n2288), .CK(net7130), .Q(
        \REGISTERS[5][17] ) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n2287), .CK(net7125), .Q(
        \REGISTERS[4][17] ) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n2286), .CK(net7120), .Q(
        \REGISTERS[3][17] ) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n2285), .CK(net7115), .Q(
        \REGISTERS[2][17] ) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n2284), .CK(net7110), .Q(
        \REGISTERS[1][17] ) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n2283), .CK(net7104), .Q(
        \REGISTERS[0][17] ) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n2282), .CK(net7260), .Q(
        \REGISTERS[31][14] ) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n2281), .CK(net7200), .Q(
        \REGISTERS[19][14] ) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n2280), .CK(net7190), .Q(
        \REGISTERS[17][14] ) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n2279), .CK(net7180), .Q(
        \REGISTERS[15][14] ) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n2278), .CK(net7140), .Q(
        \REGISTERS[7][14] ) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n2277), .CK(net7135), .Q(
        \REGISTERS[6][14] ) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n2276), .CK(net7130), .Q(
        \REGISTERS[5][14] ) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n2275), .CK(net7125), .Q(
        \REGISTERS[4][14] ) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n2274), .CK(net7120), .Q(
        \REGISTERS[3][14] ) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n2273), .CK(net7115), .Q(
        \REGISTERS[2][14] ) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n2272), .CK(net7110), .Q(
        \REGISTERS[1][14] ) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n2271), .CK(net7104), .Q(
        \REGISTERS[0][14] ) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n2270), .CK(net7260), .Q(
        \REGISTERS[31][22] ) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n2269), .CK(net7255), .Q(
        \REGISTERS[30][22] ) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n2268), .CK(net7250), .Q(
        \REGISTERS[29][22] ) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n2267), .CK(net7245), .Q(
        \REGISTERS[28][22] ) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n2266), .CK(net7240), .Q(
        \REGISTERS[27][22] ) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n2265), .CK(net7235), .Q(
        \REGISTERS[26][22] ) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n2264), .CK(net7230), .Q(
        \REGISTERS[25][22] ) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n2263), .CK(net7225), .Q(
        \REGISTERS[24][22] ) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n2262), .CK(net7220), .Q(
        \REGISTERS[23][22] ) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n2261), .CK(net7215), .Q(
        \REGISTERS[22][22] ) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n2260), .CK(net7210), .Q(
        \REGISTERS[21][22] ) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n2259), .CK(net7200), .Q(
        \REGISTERS[19][22] ) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n2258), .CK(net7190), .Q(
        \REGISTERS[17][22] ) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n2257), .CK(net7180), .Q(
        \REGISTERS[15][22] ) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n2256), .CK(net7140), .Q(
        \REGISTERS[7][22] ) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n2255), .CK(net7135), .Q(
        \REGISTERS[6][22] ) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n2254), .CK(net7130), .Q(
        \REGISTERS[5][22] ) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n2253), .CK(net7125), .Q(
        \REGISTERS[4][22] ) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n2252), .CK(net7120), .Q(
        \REGISTERS[3][22] ) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n2251), .CK(net7115), .Q(
        \REGISTERS[2][22] ) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n2250), .CK(net7110), .Q(
        \REGISTERS[1][22] ) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n2249), .CK(net7104), .Q(
        \REGISTERS[0][22] ) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n2248), .CK(net7260), .Q(
        \REGISTERS[31][25] ) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n2247), .CK(net7255), .Q(
        \REGISTERS[30][25] ) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n2246), .CK(net7250), .Q(
        \REGISTERS[29][25] ) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n2245), .CK(net7245), .Q(
        \REGISTERS[28][25] ) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n2244), .CK(net7240), .Q(
        \REGISTERS[27][25] ) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n2243), .CK(net7235), .Q(
        \REGISTERS[26][25] ) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n2242), .CK(net7230), .Q(
        \REGISTERS[25][25] ) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n2241), .CK(net7225), .Q(
        \REGISTERS[24][25] ) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n2240), .CK(net7220), .Q(
        \REGISTERS[23][25] ) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n2239), .CK(net7215), .Q(
        \REGISTERS[22][25] ) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n2238), .CK(net7210), .Q(
        \REGISTERS[21][25] ) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n2237), .CK(net7205), .Q(
        \REGISTERS[20][25] ) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n2236), .CK(net7200), .Q(
        \REGISTERS[19][25] ) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n2235), .CK(net7195), .Q(
        \REGISTERS[18][25] ) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n2234), .CK(net7190), .Q(
        \REGISTERS[17][25] ) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n2233), .CK(net7185), .Q(
        \REGISTERS[16][25] ) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n2232), .CK(net7180), .Q(
        \REGISTERS[15][25] ) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n2231), .CK(net7175), .Q(
        \REGISTERS[14][25] ) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n2230), .CK(net7170), .Q(
        \REGISTERS[13][25] ) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n2229), .CK(net7165), .Q(
        \REGISTERS[12][25] ) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n2228), .CK(net7160), .Q(
        \REGISTERS[11][25] ) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n2227), .CK(net7155), .Q(
        \REGISTERS[10][25] ) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n2226), .CK(net7150), .Q(
        \REGISTERS[9][25] ) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n2225), .CK(net7145), .Q(
        \REGISTERS[8][25] ) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n2224), .CK(net7140), .Q(
        \REGISTERS[7][25] ) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n2223), .CK(net7135), .Q(
        \REGISTERS[6][25] ) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n2222), .CK(net7130), .Q(
        \REGISTERS[5][25] ) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n2221), .CK(net7125), .Q(
        \REGISTERS[4][25] ) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n2220), .CK(net7120), .Q(
        \REGISTERS[3][25] ) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n2219), .CK(net7115), .Q(
        \REGISTERS[2][25] ) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n2218), .CK(net7110), .Q(
        \REGISTERS[1][25] ) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n2217), .CK(net7104), .Q(
        \REGISTERS[0][25] ) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n2216), .CK(net7260), .Q(
        \REGISTERS[31][20] ) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n2215), .CK(net7255), .Q(
        \REGISTERS[30][20] ) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n2214), .CK(net7250), .Q(
        \REGISTERS[29][20] ) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n2213), .CK(net7245), .Q(
        \REGISTERS[28][20] ) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n2212), .CK(net7240), .Q(
        \REGISTERS[27][20] ) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n2211), .CK(net7235), .Q(
        \REGISTERS[26][20] ) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n2210), .CK(net7230), .Q(
        \REGISTERS[25][20] ) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n2209), .CK(net7225), .Q(
        \REGISTERS[24][20] ) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n2208), .CK(net7220), .Q(
        \REGISTERS[23][20] ) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n2207), .CK(net7215), .Q(
        \REGISTERS[22][20] ) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n2206), .CK(net7210), .Q(
        \REGISTERS[21][20] ) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n2205), .CK(net7205), .Q(
        \REGISTERS[20][20] ) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n2204), .CK(net7200), .Q(
        \REGISTERS[19][20] ) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n2203), .CK(net7195), .Q(
        \REGISTERS[18][20] ) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n2202), .CK(net7190), .Q(
        \REGISTERS[17][20] ) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n2201), .CK(net7185), .Q(
        \REGISTERS[16][20] ) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n2200), .CK(net7180), .Q(
        \REGISTERS[15][20] ) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n2199), .CK(net7175), .Q(
        \REGISTERS[14][20] ) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n2198), .CK(net7170), .Q(
        \REGISTERS[13][20] ) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n2197), .CK(net7165), .Q(
        \REGISTERS[12][20] ) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n2196), .CK(net7160), .Q(
        \REGISTERS[11][20] ) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n2195), .CK(net7155), .Q(
        \REGISTERS[10][20] ) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n2194), .CK(net7150), .Q(
        \REGISTERS[9][20] ) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n2193), .CK(net7145), .Q(
        \REGISTERS[8][20] ) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n2192), .CK(net7140), .Q(
        \REGISTERS[7][20] ) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n2191), .CK(net7135), .Q(
        \REGISTERS[6][20] ) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n2190), .CK(net7130), .Q(
        \REGISTERS[5][20] ) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n2189), .CK(net7125), .Q(
        \REGISTERS[4][20] ) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n2188), .CK(net7120), .Q(
        \REGISTERS[3][20] ) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n2187), .CK(net7115), .Q(
        \REGISTERS[2][20] ) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n2186), .CK(net7110), .Q(
        \REGISTERS[1][20] ) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n2185), .CK(net7104), .Q(
        \REGISTERS[0][20] ) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n2184), .CK(net7255), .Q(
        \REGISTERS[30][3] ) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n2183), .CK(net7250), .Q(
        \REGISTERS[29][3] ) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n2182), .CK(net7245), .Q(
        \REGISTERS[28][3] ) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n2181), .CK(net7240), .Q(
        \REGISTERS[27][3] ) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n2180), .CK(net7235), .Q(
        \REGISTERS[26][3] ) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n2179), .CK(net7230), .Q(
        \REGISTERS[25][3] ) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n2178), .CK(net7225), .Q(
        \REGISTERS[24][3] ) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n2177), .CK(net7220), .Q(
        \REGISTERS[23][3] ) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n2176), .CK(net7215), .Q(
        \REGISTERS[22][3] ) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n2175), .CK(net7210), .Q(
        \REGISTERS[21][3] ) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n2174), .CK(net7260), .Q(
        \REGISTERS[31][3] ) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n2173), .CK(net7200), .Q(
        \REGISTERS[19][3] ) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n2172), .CK(net7190), .Q(
        \REGISTERS[17][3] ) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n2171), .CK(net7180), .Q(
        \REGISTERS[15][3] ) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n2170), .CK(net7140), .Q(\REGISTERS[7][3] ) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n2169), .CK(net7135), .Q(\REGISTERS[6][3] ) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n2168), .CK(net7130), .Q(\REGISTERS[5][3] ) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n2167), .CK(net7125), .Q(\REGISTERS[4][3] ) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n2166), .CK(net7120), .Q(\REGISTERS[3][3] ) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n2165), .CK(net7115), .Q(\REGISTERS[2][3] ) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n2164), .CK(net7110), .Q(\REGISTERS[1][3] ) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n2163), .CK(net7104), .Q(\REGISTERS[0][3] ) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n2162), .CK(net7260), .Q(
        \REGISTERS[31][2] ) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n2161), .CK(net7255), .Q(
        \REGISTERS[30][2] ) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n2160), .CK(net7250), .Q(
        \REGISTERS[29][2] ) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n2159), .CK(net7245), .Q(
        \REGISTERS[28][2] ) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n2158), .CK(net7240), .Q(
        \REGISTERS[27][2] ) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n2157), .CK(net7235), .Q(
        \REGISTERS[26][2] ) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n2156), .CK(net7230), .Q(
        \REGISTERS[25][2] ) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n2155), .CK(net7225), .Q(
        \REGISTERS[24][2] ) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n2154), .CK(net7220), .Q(
        \REGISTERS[23][2] ) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n2153), .CK(net7215), .Q(
        \REGISTERS[22][2] ) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n2152), .CK(net7210), .Q(
        \REGISTERS[21][2] ) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n2151), .CK(net7200), .Q(
        \REGISTERS[19][2] ) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n2150), .CK(net7190), .Q(
        \REGISTERS[17][2] ) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n2149), .CK(net7180), .Q(
        \REGISTERS[15][2] ) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n2148), .CK(net7140), .Q(\REGISTERS[7][2] ) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n2147), .CK(net7135), .Q(\REGISTERS[6][2] ) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n2146), .CK(net7130), .Q(\REGISTERS[5][2] ) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n2145), .CK(net7125), .Q(\REGISTERS[4][2] ) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n2144), .CK(net7120), .Q(\REGISTERS[3][2] ) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n2143), .CK(net7115), .Q(\REGISTERS[2][2] ) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n2142), .CK(net7110), .Q(\REGISTERS[1][2] ) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n2141), .CK(net7104), .Q(\REGISTERS[0][2] ) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n2140), .CK(net7205), .Q(
        \REGISTERS[20][2] ) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n2139), .CK(net7195), .Q(
        \REGISTERS[18][2] ) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n2138), .CK(net7185), .Q(
        \REGISTERS[16][2] ) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n2137), .CK(net7175), .Q(
        \REGISTERS[14][2] ) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n2136), .CK(net7170), .Q(
        \REGISTERS[13][2] ) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n2135), .CK(net7165), .Q(
        \REGISTERS[12][2] ) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n2134), .CK(net7160), .Q(
        \REGISTERS[11][2] ) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n2133), .CK(net7155), .Q(
        \REGISTERS[10][2] ) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n2132), .CK(net7150), .Q(\REGISTERS[9][2] ) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n2131), .CK(net7145), .Q(\REGISTERS[8][2] ) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n2130), .CK(net7260), .Q(
        \REGISTERS[31][19] ) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n2129), .CK(net7255), .Q(
        \REGISTERS[30][19] ) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n2128), .CK(net7250), .Q(
        \REGISTERS[29][19] ) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n2127), .CK(net7245), .Q(
        \REGISTERS[28][19] ) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n2126), .CK(net7240), .Q(
        \REGISTERS[27][19] ) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n2125), .CK(net7235), .Q(
        \REGISTERS[26][19] ) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n2124), .CK(net7230), .Q(
        \REGISTERS[25][19] ) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n2123), .CK(net7225), .Q(
        \REGISTERS[24][19] ) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n2122), .CK(net7220), .Q(
        \REGISTERS[23][19] ) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n2121), .CK(net7215), .Q(
        \REGISTERS[22][19] ) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n2120), .CK(net7210), .Q(
        \REGISTERS[21][19] ) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n2119), .CK(net7200), .Q(
        \REGISTERS[19][19] ) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n2118), .CK(net7190), .Q(
        \REGISTERS[17][19] ) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n2117), .CK(net7180), .Q(
        \REGISTERS[15][19] ) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n2116), .CK(net7140), .Q(
        \REGISTERS[7][19] ) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n2115), .CK(net7135), .Q(
        \REGISTERS[6][19] ) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n2114), .CK(net7130), .Q(
        \REGISTERS[5][19] ) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n2113), .CK(net7125), .Q(
        \REGISTERS[4][19] ) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n2112), .CK(net7120), .Q(
        \REGISTERS[3][19] ) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n2111), .CK(net7115), .Q(
        \REGISTERS[2][19] ) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n2110), .CK(net7110), .Q(
        \REGISTERS[1][19] ) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n2109), .CK(net7104), .Q(
        \REGISTERS[0][19] ) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n2108), .CK(net7260), .Q(
        \REGISTERS[31][10] ) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n2107), .CK(net7255), .Q(
        \REGISTERS[30][10] ) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n2106), .CK(net7250), .Q(
        \REGISTERS[29][10] ) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n2105), .CK(net7245), .Q(
        \REGISTERS[28][10] ) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n2104), .CK(net7240), .Q(
        \REGISTERS[27][10] ) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n2103), .CK(net7235), .Q(
        \REGISTERS[26][10] ) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n2102), .CK(net7230), .Q(
        \REGISTERS[25][10] ) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n2101), .CK(net7225), .Q(
        \REGISTERS[24][10] ) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n2100), .CK(net7220), .Q(
        \REGISTERS[23][10] ) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n2099), .CK(net7215), .Q(
        \REGISTERS[22][10] ) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n2098), .CK(net7210), .Q(
        \REGISTERS[21][10] ) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n2097), .CK(net7200), .Q(
        \REGISTERS[19][10] ) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n2096), .CK(net7190), .Q(
        \REGISTERS[17][10] ) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n2095), .CK(net7180), .Q(
        \REGISTERS[15][10] ) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n2094), .CK(net7140), .Q(
        \REGISTERS[7][10] ) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n2093), .CK(net7135), .Q(
        \REGISTERS[6][10] ) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n2092), .CK(net7130), .Q(
        \REGISTERS[5][10] ) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n2091), .CK(net7125), .Q(
        \REGISTERS[4][10] ) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n2090), .CK(net7120), .Q(
        \REGISTERS[3][10] ) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n2089), .CK(net7115), .Q(
        \REGISTERS[2][10] ) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n2088), .CK(net7110), .Q(
        \REGISTERS[1][10] ) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n2087), .CK(net7104), .Q(
        \REGISTERS[0][10] ) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n2086), .CK(net7255), .Q(
        \REGISTERS[30][28] ) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n2085), .CK(net7250), .Q(
        \REGISTERS[29][28] ) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n2084), .CK(net7245), .Q(
        \REGISTERS[28][28] ) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n2083), .CK(net7240), .Q(
        \REGISTERS[27][28] ) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n2082), .CK(net7235), .Q(
        \REGISTERS[26][28] ) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n2081), .CK(net7230), .Q(
        \REGISTERS[25][28] ) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n2080), .CK(net7225), .Q(
        \REGISTERS[24][28] ) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n2079), .CK(net7220), .Q(
        \REGISTERS[23][28] ) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n2078), .CK(net7215), .Q(
        \REGISTERS[22][28] ) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n2077), .CK(net7210), .Q(
        \REGISTERS[21][28] ) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n2076), .CK(net7205), .Q(
        \REGISTERS[20][28] ) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n2075), .CK(net7200), .Q(
        \REGISTERS[19][28] ) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n2074), .CK(net7195), .Q(
        \REGISTERS[18][28] ) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n2073), .CK(net7190), .Q(
        \REGISTERS[17][28] ) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n2072), .CK(net7185), .Q(
        \REGISTERS[16][28] ) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n2071), .CK(net7180), .Q(
        \REGISTERS[15][28] ) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n2070), .CK(net7175), .Q(
        \REGISTERS[14][28] ) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n2069), .CK(net7170), .Q(
        \REGISTERS[13][28] ) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n2068), .CK(net7165), .Q(
        \REGISTERS[12][28] ) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n2067), .CK(net7160), .Q(
        \REGISTERS[11][28] ) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n2066), .CK(net7155), .Q(
        \REGISTERS[10][28] ) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n2065), .CK(net7150), .Q(
        \REGISTERS[9][28] ) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n2064), .CK(net7145), .Q(
        \REGISTERS[8][28] ) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n2063), .CK(net7140), .Q(
        \REGISTERS[7][28] ) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n2062), .CK(net7135), .Q(
        \REGISTERS[6][28] ) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n2061), .CK(net7130), .Q(
        \REGISTERS[5][28] ) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n2060), .CK(net7125), .Q(
        \REGISTERS[4][28] ) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n2059), .CK(net7120), .Q(
        \REGISTERS[3][28] ) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n2058), .CK(net7115), .Q(
        \REGISTERS[2][28] ) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n2057), .CK(net7110), .Q(
        \REGISTERS[1][28] ) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n2056), .CK(net7104), .Q(
        \REGISTERS[0][28] ) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n2055), .CK(net7260), .Q(
        \REGISTERS[31][26] ) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n2054), .CK(net7255), .Q(
        \REGISTERS[30][26] ) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n2053), .CK(net7250), .Q(
        \REGISTERS[29][26] ) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n2052), .CK(net7245), .Q(
        \REGISTERS[28][26] ) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n2051), .CK(net7240), .Q(
        \REGISTERS[27][26] ) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n2050), .CK(net7235), .Q(
        \REGISTERS[26][26] ) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n2049), .CK(net7230), .Q(
        \REGISTERS[25][26] ) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n2048), .CK(net7225), .Q(
        \REGISTERS[24][26] ) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n2047), .CK(net7220), .Q(
        \REGISTERS[23][26] ) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n2046), .CK(net7215), .Q(
        \REGISTERS[22][26] ) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n2045), .CK(net7210), .Q(
        \REGISTERS[21][26] ) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n2044), .CK(net7200), .Q(
        \REGISTERS[19][26] ) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n2043), .CK(net7190), .Q(
        \REGISTERS[17][26] ) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n2042), .CK(net7180), .Q(
        \REGISTERS[15][26] ) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n2041), .CK(net7140), .Q(
        \REGISTERS[7][26] ) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n2040), .CK(net7135), .Q(
        \REGISTERS[6][26] ) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n2039), .CK(net7130), .Q(
        \REGISTERS[5][26] ) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n2038), .CK(net7125), .Q(
        \REGISTERS[4][26] ) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n2037), .CK(net7120), .Q(
        \REGISTERS[3][26] ) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n2036), .CK(net7115), .Q(
        \REGISTERS[2][26] ) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n2035), .CK(net7110), .Q(
        \REGISTERS[1][26] ) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n2034), .CK(net7104), .Q(
        \REGISTERS[0][26] ) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n2033), .CK(net7260), .Q(
        \REGISTERS[31][6] ) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n2032), .CK(net7255), .Q(
        \REGISTERS[30][6] ) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n2031), .CK(net7250), .Q(
        \REGISTERS[29][6] ) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n2030), .CK(net7245), .Q(
        \REGISTERS[28][6] ) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n2029), .CK(net7240), .Q(
        \REGISTERS[27][6] ) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n2028), .CK(net7235), .Q(
        \REGISTERS[26][6] ) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n2027), .CK(net7230), .Q(
        \REGISTERS[25][6] ) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n2026), .CK(net7225), .Q(
        \REGISTERS[24][6] ) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n2025), .CK(net7220), .Q(
        \REGISTERS[23][6] ) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n2024), .CK(net7215), .Q(
        \REGISTERS[22][6] ) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n2023), .CK(net7210), .Q(
        \REGISTERS[21][6] ) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n2022), .CK(net7200), .Q(
        \REGISTERS[19][6] ) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n2021), .CK(net7195), .Q(
        \REGISTERS[18][6] ) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n2020), .CK(net7190), .Q(
        \REGISTERS[17][6] ) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n2019), .CK(net7185), .Q(
        \REGISTERS[16][6] ) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n2018), .CK(net7180), .Q(
        \REGISTERS[15][6] ) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n2017), .CK(net7175), .Q(
        \REGISTERS[14][6] ) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n2016), .CK(net7170), .Q(
        \REGISTERS[13][6] ) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n2015), .CK(net7165), .Q(
        \REGISTERS[12][6] ) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n2014), .CK(net7160), .Q(
        \REGISTERS[11][6] ) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n2013), .CK(net7155), .Q(
        \REGISTERS[10][6] ) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n2012), .CK(net7150), .Q(\REGISTERS[9][6] ) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n2011), .CK(net7145), .Q(\REGISTERS[8][6] ) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n2010), .CK(net7140), .Q(\REGISTERS[7][6] ) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n2009), .CK(net7135), .Q(\REGISTERS[6][6] ) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n2008), .CK(net7130), .Q(\REGISTERS[5][6] ) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n2007), .CK(net7125), .Q(\REGISTERS[4][6] ) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n2006), .CK(net7120), .Q(\REGISTERS[3][6] ) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n2005), .CK(net7115), .Q(\REGISTERS[2][6] ) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n2004), .CK(net7110), .Q(\REGISTERS[1][6] ) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n2003), .CK(net7104), .Q(\REGISTERS[0][6] ) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n2002), .CK(net7255), .Q(
        \REGISTERS[30][0] ) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n2001), .CK(net7245), .Q(
        \REGISTERS[28][0] ) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n2000), .CK(net7235), .Q(
        \REGISTERS[26][0] ) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n1999), .CK(net7225), .Q(
        \REGISTERS[24][0] ) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n1998), .CK(net7215), .Q(
        \REGISTERS[22][0] ) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n1997), .CK(net7200), .Q(
        \REGISTERS[19][0] ) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n1996), .CK(net7190), .Q(
        \REGISTERS[17][0] ) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n1995), .CK(net7180), .Q(
        \REGISTERS[15][0] ) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n1994), .CK(net7140), .Q(\REGISTERS[7][0] ) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n1993), .CK(net7135), .Q(\REGISTERS[6][0] ) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n1992), .CK(net7255), .Q(
        \REGISTERS[30][31] ) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n1991), .CK(net7250), .Q(
        \REGISTERS[29][31] ) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n1990), .CK(net7245), .Q(
        \REGISTERS[28][31] ) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n1989), .CK(net7240), .Q(
        \REGISTERS[27][31] ) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n1988), .CK(net7235), .Q(
        \REGISTERS[26][31] ) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n1987), .CK(net7230), .Q(
        \REGISTERS[25][31] ) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n1986), .CK(net7225), .Q(
        \REGISTERS[24][31] ) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n1985), .CK(net7220), .Q(
        \REGISTERS[23][31] ) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n1984), .CK(net7215), .Q(
        \REGISTERS[22][31] ) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n1983), .CK(net7210), .Q(
        \REGISTERS[21][31] ) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n1982), .CK(net7205), .Q(
        \REGISTERS[20][31] ) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n1981), .CK(net7200), .Q(
        \REGISTERS[19][31] ) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n1980), .CK(net7195), .Q(
        \REGISTERS[18][31] ) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n1979), .CK(net7190), .Q(
        \REGISTERS[17][31] ) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n1978), .CK(net7185), .Q(
        \REGISTERS[16][31] ) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n1977), .CK(net7180), .Q(
        \REGISTERS[15][31] ) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n1976), .CK(net7175), .Q(
        \REGISTERS[14][31] ) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n1975), .CK(net7170), .Q(
        \REGISTERS[13][31] ) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n1974), .CK(net7165), .Q(
        \REGISTERS[12][31] ) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n1973), .CK(net7160), .Q(
        \REGISTERS[11][31] ) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n1972), .CK(net7155), .Q(
        \REGISTERS[10][31] ) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n1971), .CK(net7150), .Q(
        \REGISTERS[9][31] ) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n1970), .CK(net7145), .Q(
        \REGISTERS[8][31] ) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n1969), .CK(net7140), .Q(
        \REGISTERS[7][31] ) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n1968), .CK(net7135), .Q(
        \REGISTERS[6][31] ) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n1967), .CK(net7130), .Q(
        \REGISTERS[5][31] ) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n1966), .CK(net7125), .Q(
        \REGISTERS[4][31] ) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n1965), .CK(net7120), .Q(
        \REGISTERS[3][31] ) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n1964), .CK(net7115), .Q(
        \REGISTERS[2][31] ) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n1963), .CK(net7110), .Q(
        \REGISTERS[1][31] ) );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n1962), .CK(net7104), .Q(
        \REGISTERS[0][31] ) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n1961), .CK(net7130), .Q(\REGISTERS[5][0] ) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n1960), .CK(net7125), .Q(\REGISTERS[4][0] ) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n1959), .CK(net7120), .Q(\REGISTERS[3][0] ) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n1958), .CK(net7115), .Q(\REGISTERS[2][0] ) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n1957), .CK(net7110), .Q(\REGISTERS[1][0] ) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n1956), .CK(net7104), .Q(\REGISTERS[0][0] ) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n1955), .CK(net7260), .Q(
        \REGISTERS[31][1] ) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n1954), .CK(net7255), .Q(
        \REGISTERS[30][1] ) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n1953), .CK(net7250), .Q(
        \REGISTERS[29][1] ) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n1952), .CK(net7245), .Q(
        \REGISTERS[28][1] ) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n1951), .CK(net7240), .Q(
        \REGISTERS[27][1] ) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n1950), .CK(net7235), .Q(
        \REGISTERS[26][1] ) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n1949), .CK(net7230), .Q(
        \REGISTERS[25][1] ) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n1948), .CK(net7225), .Q(
        \REGISTERS[24][1] ) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n1947), .CK(net7220), .Q(
        \REGISTERS[23][1] ) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n1946), .CK(net7215), .Q(
        \REGISTERS[22][1] ) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n1945), .CK(net7210), .Q(
        \REGISTERS[21][1] ) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n1944), .CK(net7200), .Q(
        \REGISTERS[19][1] ) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n1943), .CK(net7190), .Q(
        \REGISTERS[17][1] ) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n1942), .CK(net7180), .Q(
        \REGISTERS[15][1] ) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n1941), .CK(net7140), .Q(\REGISTERS[7][1] ) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n1940), .CK(net7135), .Q(\REGISTERS[6][1] ) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n1939), .CK(net7130), .Q(\REGISTERS[5][1] ) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n1938), .CK(net7125), .Q(\REGISTERS[4][1] ) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n1937), .CK(net7120), .Q(\REGISTERS[3][1] ) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n1936), .CK(net7115), .Q(\REGISTERS[2][1] ) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n1935), .CK(net7110), .Q(\REGISTERS[1][1] ) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n1934), .CK(net7104), .Q(\REGISTERS[0][1] ) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n1933), .CK(net7260), .Q(
        \REGISTERS[31][30] ) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n1932), .CK(net7255), .Q(
        \REGISTERS[30][30] ) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n1931), .CK(net7250), .Q(
        \REGISTERS[29][30] ) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n1930), .CK(net7245), .Q(
        \REGISTERS[28][30] ) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n1929), .CK(net7240), .Q(
        \REGISTERS[27][30] ) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n1928), .CK(net7235), .Q(
        \REGISTERS[26][30] ) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n1927), .CK(net7230), .Q(
        \REGISTERS[25][30] ) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n1926), .CK(net7225), .Q(
        \REGISTERS[24][30] ) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n1925), .CK(net7220), .Q(
        \REGISTERS[23][30] ) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n1924), .CK(net7215), .Q(
        \REGISTERS[22][30] ) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n1923), .CK(net7210), .Q(
        \REGISTERS[21][30] ) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n1922), .CK(net7200), .Q(
        \REGISTERS[19][30] ) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n1921), .CK(net7190), .Q(
        \REGISTERS[17][30] ) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n1920), .CK(net7180), .Q(
        \REGISTERS[15][30] ) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n1919), .CK(net7140), .Q(
        \REGISTERS[7][30] ) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n1918), .CK(net7135), .Q(
        \REGISTERS[6][30] ) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n1917), .CK(net7130), .Q(
        \REGISTERS[5][30] ) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n1916), .CK(net7125), .Q(
        \REGISTERS[4][30] ) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n1915), .CK(net7120), .Q(
        \REGISTERS[3][30] ) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n1914), .CK(net7115), .Q(
        \REGISTERS[2][30] ) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n1913), .CK(net7110), .Q(
        \REGISTERS[1][30] ) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n1912), .CK(net7104), .Q(
        \REGISTERS[0][30] ) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n1911), .CK(net7255), .Q(
        \REGISTERS[30][7] ) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n1910), .CK(net7245), .Q(
        \REGISTERS[28][7] ) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n1909), .CK(net7235), .Q(
        \REGISTERS[26][7] ) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n1908), .CK(net7225), .Q(
        \REGISTERS[24][7] ) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n1907), .CK(net7215), .Q(
        \REGISTERS[22][7] ) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n1906), .CK(net7200), .Q(
        \REGISTERS[19][7] ) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n1905), .CK(net7190), .Q(
        \REGISTERS[17][7] ) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n1904), .CK(net7180), .Q(
        \REGISTERS[15][7] ) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n1903), .CK(net7140), .Q(\REGISTERS[7][7] ) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n1902), .CK(net7135), .Q(\REGISTERS[6][7] ) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n1901), .CK(net7130), .Q(\REGISTERS[5][7] ) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n1900), .CK(net7125), .Q(\REGISTERS[4][7] ) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n1899), .CK(net7120), .Q(\REGISTERS[3][7] ) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n1898), .CK(net7115), .Q(\REGISTERS[2][7] ) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n1897), .CK(net7110), .Q(\REGISTERS[1][7] ) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n1896), .CK(net7104), .Q(\REGISTERS[0][7] ) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n1895), .CK(net7140), .Q(
        \REGISTERS[7][15] ) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n1894), .CK(net7135), .Q(
        \REGISTERS[6][15] ) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n1893), .CK(net7130), .Q(
        \REGISTERS[5][15] ) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n1892), .CK(net7125), .Q(
        \REGISTERS[4][15] ) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n1891), .CK(net7120), .Q(
        \REGISTERS[3][15] ) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n1890), .CK(net7115), .Q(
        \REGISTERS[2][15] ) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n1889), .CK(net7255), .Q(
        \REGISTERS[30][15] ) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n1888), .CK(net7245), .Q(
        \REGISTERS[28][15] ) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n1887), .CK(net7235), .Q(
        \REGISTERS[26][15] ) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n1886), .CK(net7225), .Q(
        \REGISTERS[24][15] ) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n1885), .CK(net7215), .Q(
        \REGISTERS[22][15] ) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n1884), .CK(net7200), .Q(
        \REGISTERS[19][15] ) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n1883), .CK(net7190), .Q(
        \REGISTERS[17][15] ) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n1882), .CK(net7180), .Q(
        \REGISTERS[15][15] ) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n1881), .CK(net7110), .Q(
        \REGISTERS[1][15] ) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n1880), .CK(net7104), .Q(
        \REGISTERS[0][15] ) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n1879), .CK(net7255), .Q(
        \REGISTERS[30][23] ) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n1878), .CK(net7250), .Q(
        \REGISTERS[29][23] ) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n1877), .CK(net7245), .Q(
        \REGISTERS[28][23] ) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n1876), .CK(net7240), .Q(
        \REGISTERS[27][23] ) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n1875), .CK(net7235), .Q(
        \REGISTERS[26][23] ) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n1874), .CK(net7230), .Q(
        \REGISTERS[25][23] ) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n1873), .CK(net7225), .Q(
        \REGISTERS[24][23] ) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n1872), .CK(net7220), .Q(
        \REGISTERS[23][23] ) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n1871), .CK(net7215), .Q(
        \REGISTERS[22][23] ) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n1870), .CK(net7210), .Q(
        \REGISTERS[21][23] ) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n1869), .CK(net7260), .Q(
        \REGISTERS[31][8] ) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n1868), .CK(net7255), .Q(
        \REGISTERS[30][8] ) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n1867), .CK(net7250), .Q(
        \REGISTERS[29][8] ) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n1866), .CK(net7245), .Q(
        \REGISTERS[28][8] ) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n1865), .CK(net7240), .Q(
        \REGISTERS[27][8] ) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n1864), .CK(net7235), .Q(
        \REGISTERS[26][8] ) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n1863), .CK(net7230), .Q(
        \REGISTERS[25][8] ) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n1862), .CK(net7225), .Q(
        \REGISTERS[24][8] ) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n1861), .CK(net7220), .Q(
        \REGISTERS[23][8] ) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n1860), .CK(net7215), .Q(
        \REGISTERS[22][8] ) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n1859), .CK(net7210), .Q(
        \REGISTERS[21][8] ) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n1858), .CK(net7200), .Q(
        \REGISTERS[19][8] ) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n1857), .CK(net7190), .Q(
        \REGISTERS[17][8] ) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n1856), .CK(net7180), .Q(
        \REGISTERS[15][8] ) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n1855), .CK(net7140), .Q(\REGISTERS[7][8] ) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n1854), .CK(net7135), .Q(\REGISTERS[6][8] ) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n1853), .CK(net7130), .Q(\REGISTERS[5][8] ) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n1852), .CK(net7125), .Q(\REGISTERS[4][8] ) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n1851), .CK(net7120), .Q(\REGISTERS[3][8] ) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n1850), .CK(net7115), .Q(\REGISTERS[2][8] ) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n1849), .CK(net7110), .Q(\REGISTERS[1][8] ) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n1848), .CK(net7104), .Q(\REGISTERS[0][8] ) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n1847), .CK(net7260), .Q(
        \REGISTERS[31][23] ) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n1846), .CK(net7200), .Q(
        \REGISTERS[19][23] ) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n1845), .CK(net7190), .Q(
        \REGISTERS[17][23] ) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n1844), .CK(net7180), .Q(
        \REGISTERS[15][23] ) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n1843), .CK(net7140), .Q(
        \REGISTERS[7][23] ) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n1842), .CK(net7135), .Q(
        \REGISTERS[6][23] ) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n1841), .CK(net7130), .Q(
        \REGISTERS[5][23] ) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n1840), .CK(net7125), .Q(
        \REGISTERS[4][23] ) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n1839), .CK(net7120), .Q(
        \REGISTERS[3][23] ) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n1838), .CK(net7115), .Q(
        \REGISTERS[2][23] ) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n1837), .CK(net7110), .Q(
        \REGISTERS[1][23] ) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n1836), .CK(net7104), .Q(
        \REGISTERS[0][23] ) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n1835), .CK(net7260), .Q(
        \REGISTERS[31][4] ) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n1834), .CK(net7255), .Q(
        \REGISTERS[30][4] ) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n1833), .CK(net7250), .Q(
        \REGISTERS[29][4] ) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n1832), .CK(net7245), .Q(
        \REGISTERS[28][4] ) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n1831), .CK(net7240), .Q(
        \REGISTERS[27][4] ) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n1830), .CK(net7235), .Q(
        \REGISTERS[26][4] ) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n1829), .CK(net7230), .Q(
        \REGISTERS[25][4] ) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n1828), .CK(net7225), .Q(
        \REGISTERS[24][4] ) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n1827), .CK(net7220), .Q(
        \REGISTERS[23][4] ) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n1826), .CK(net7215), .Q(
        \REGISTERS[22][4] ) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n1825), .CK(net7210), .Q(
        \REGISTERS[21][4] ) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n1824), .CK(net7200), .Q(
        \REGISTERS[19][4] ) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n1823), .CK(net7190), .Q(
        \REGISTERS[17][4] ) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n1822), .CK(net7180), .Q(
        \REGISTERS[15][4] ) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n1821), .CK(net7140), .Q(\REGISTERS[7][4] ) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n1820), .CK(net7135), .Q(\REGISTERS[6][4] ) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n1819), .CK(net7130), .Q(\REGISTERS[5][4] ) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n1818), .CK(net7125), .Q(\REGISTERS[4][4] ) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n1817), .CK(net7120), .Q(\REGISTERS[3][4] ) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n1816), .CK(net7115), .Q(\REGISTERS[2][4] ) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n1815), .CK(net7110), .Q(\REGISTERS[1][4] ) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n1814), .CK(net7104), .Q(\REGISTERS[0][4] ) );
  CLKBUF_X2 U13 ( .A(n144), .Z(n146) );
  CLKBUF_X2 U18 ( .A(n149), .Z(n144) );
  CLKBUF_X2 U19 ( .A(RST), .Z(n139) );
  CLKBUF_X2 U21 ( .A(RST), .Z(n149) );
  AND2_X1 U1906 ( .A1(n127), .A2(RST), .ZN(n1814) );
  AND2_X1 U1907 ( .A1(n127), .A2(RST), .ZN(n1815) );
  AND2_X1 U1908 ( .A1(n127), .A2(n153), .ZN(n1816) );
  AND2_X1 U1909 ( .A1(n127), .A2(n151), .ZN(n1817) );
  AND2_X1 U1910 ( .A1(n127), .A2(n152), .ZN(n1818) );
  AND2_X1 U1911 ( .A1(n127), .A2(RST), .ZN(n1819) );
  AND2_X1 U1912 ( .A1(n127), .A2(n150), .ZN(n1820) );
  AND2_X1 U1913 ( .A1(n127), .A2(n152), .ZN(n1821) );
  AND2_X1 U1914 ( .A1(n127), .A2(RST), .ZN(n1822) );
  AND2_X1 U1915 ( .A1(n127), .A2(n138), .ZN(n1823) );
  AND2_X1 U1916 ( .A1(n127), .A2(RST), .ZN(n1824) );
  AND2_X1 U1917 ( .A1(n127), .A2(RST), .ZN(n1825) );
  AND2_X1 U1918 ( .A1(n127), .A2(RST), .ZN(n1826) );
  AND2_X1 U1919 ( .A1(n127), .A2(n144), .ZN(n1827) );
  AND2_X1 U1920 ( .A1(n127), .A2(n137), .ZN(n1828) );
  AND2_X1 U1921 ( .A1(n127), .A2(RST), .ZN(n1829) );
  AND2_X1 U1922 ( .A1(n127), .A2(n142), .ZN(n1830) );
  AND2_X1 U1923 ( .A1(n127), .A2(n140), .ZN(n1831) );
  AND2_X1 U1924 ( .A1(n127), .A2(n138), .ZN(n1832) );
  AND2_X1 U1925 ( .A1(n127), .A2(n152), .ZN(n1833) );
  AND2_X1 U1926 ( .A1(n127), .A2(RST), .ZN(n1834) );
  AND2_X1 U1927 ( .A1(n127), .A2(n153), .ZN(n1835) );
  AND2_X1 U1928 ( .A1(n89), .A2(n154), .ZN(n1836) );
  AND2_X1 U1929 ( .A1(n89), .A2(n152), .ZN(n1837) );
  AND2_X1 U1930 ( .A1(n89), .A2(n145), .ZN(n1838) );
  AND2_X1 U1931 ( .A1(n89), .A2(n153), .ZN(n1839) );
  AND2_X1 U1932 ( .A1(n89), .A2(n153), .ZN(n1840) );
  AND2_X1 U1933 ( .A1(n89), .A2(n152), .ZN(n1841) );
  AND2_X1 U1934 ( .A1(n89), .A2(n148), .ZN(n1842) );
  AND2_X1 U1935 ( .A1(n89), .A2(n150), .ZN(n1843) );
  AND2_X1 U1936 ( .A1(n89), .A2(n144), .ZN(n1844) );
  AND2_X1 U1937 ( .A1(n89), .A2(n143), .ZN(n1845) );
  AND2_X1 U1938 ( .A1(n89), .A2(RST), .ZN(n1846) );
  AND2_X1 U1939 ( .A1(n89), .A2(n151), .ZN(n1847) );
  AND2_X1 U1940 ( .A1(n119), .A2(n155), .ZN(n1848) );
  AND2_X1 U1941 ( .A1(n119), .A2(RST), .ZN(n1849) );
  AND2_X1 U1942 ( .A1(n119), .A2(n154), .ZN(n1850) );
  AND2_X1 U1943 ( .A1(n119), .A2(n149), .ZN(n1851) );
  AND2_X1 U1944 ( .A1(n119), .A2(RST), .ZN(n1852) );
  AND2_X1 U1945 ( .A1(n119), .A2(n154), .ZN(n1853) );
  AND2_X1 U1946 ( .A1(n119), .A2(n151), .ZN(n1854) );
  AND2_X1 U1947 ( .A1(n119), .A2(n153), .ZN(n1855) );
  AND2_X1 U1948 ( .A1(n119), .A2(n143), .ZN(n1856) );
  AND2_X1 U1949 ( .A1(n119), .A2(n147), .ZN(n1857) );
  AND2_X1 U1950 ( .A1(n119), .A2(n138), .ZN(n1858) );
  AND2_X1 U1951 ( .A1(n119), .A2(RST), .ZN(n1859) );
  AND2_X1 U1952 ( .A1(n119), .A2(n138), .ZN(n1860) );
  AND2_X1 U1953 ( .A1(n119), .A2(n139), .ZN(n1861) );
  AND2_X1 U1954 ( .A1(n119), .A2(RST), .ZN(n1862) );
  AND2_X1 U1955 ( .A1(n119), .A2(n138), .ZN(n1863) );
  AND2_X1 U1956 ( .A1(n119), .A2(n145), .ZN(n1864) );
  AND2_X1 U1957 ( .A1(n119), .A2(n141), .ZN(n1865) );
  AND2_X1 U1958 ( .A1(n119), .A2(n139), .ZN(n1866) );
  AND2_X1 U1959 ( .A1(n119), .A2(n137), .ZN(n1867) );
  AND2_X1 U1960 ( .A1(n119), .A2(RST), .ZN(n1868) );
  AND2_X1 U1961 ( .A1(n119), .A2(n154), .ZN(n1869) );
  AND2_X1 U1962 ( .A1(n89), .A2(RST), .ZN(n1870) );
  AND2_X1 U1963 ( .A1(n89), .A2(RST), .ZN(n1871) );
  AND2_X1 U1964 ( .A1(n89), .A2(RST), .ZN(n1872) );
  AND2_X1 U1965 ( .A1(n89), .A2(n150), .ZN(n1873) );
  AND2_X1 U1966 ( .A1(n89), .A2(n154), .ZN(n1874) );
  AND2_X1 U1967 ( .A1(n89), .A2(n138), .ZN(n1875) );
  AND2_X1 U1968 ( .A1(n89), .A2(n142), .ZN(n1876) );
  AND2_X1 U1969 ( .A1(n89), .A2(n140), .ZN(n1877) );
  AND2_X1 U1970 ( .A1(n89), .A2(n138), .ZN(n1878) );
  AND2_X1 U1971 ( .A1(n89), .A2(n148), .ZN(n1879) );
  AND2_X1 U1972 ( .A1(n105), .A2(n155), .ZN(n1880) );
  AND2_X1 U1973 ( .A1(n105), .A2(RST), .ZN(n1881) );
  AND2_X1 U1974 ( .A1(n105), .A2(n153), .ZN(n1882) );
  AND2_X1 U1975 ( .A1(n105), .A2(RST), .ZN(n1883) );
  AND2_X1 U1976 ( .A1(n105), .A2(n140), .ZN(n1884) );
  AND2_X1 U1977 ( .A1(n105), .A2(n142), .ZN(n1885) );
  AND2_X1 U1978 ( .A1(n105), .A2(n149), .ZN(n1886) );
  AND2_X1 U1979 ( .A1(n105), .A2(n145), .ZN(n1887) );
  AND2_X1 U1980 ( .A1(n105), .A2(n139), .ZN(n1888) );
  AND2_X1 U1981 ( .A1(n105), .A2(RST), .ZN(n1889) );
  AND2_X1 U1982 ( .A1(n105), .A2(n154), .ZN(n1890) );
  AND2_X1 U1983 ( .A1(n105), .A2(n152), .ZN(n1891) );
  AND2_X1 U1984 ( .A1(n105), .A2(RST), .ZN(n1892) );
  AND2_X1 U1985 ( .A1(n105), .A2(RST), .ZN(n1893) );
  AND2_X1 U1986 ( .A1(n105), .A2(n151), .ZN(n1894) );
  AND2_X1 U1987 ( .A1(n105), .A2(n155), .ZN(n1895) );
  AND2_X1 U1988 ( .A1(n121), .A2(n155), .ZN(n1896) );
  AND2_X1 U1989 ( .A1(n121), .A2(RST), .ZN(n1897) );
  AND2_X1 U1990 ( .A1(n121), .A2(n154), .ZN(n1898) );
  AND2_X1 U1991 ( .A1(n121), .A2(RST), .ZN(n1899) );
  AND2_X1 U1992 ( .A1(n121), .A2(RST), .ZN(n1900) );
  AND2_X1 U1993 ( .A1(n121), .A2(RST), .ZN(n1901) );
  AND2_X1 U1994 ( .A1(n121), .A2(n151), .ZN(n1902) );
  AND2_X1 U1995 ( .A1(n121), .A2(RST), .ZN(n1903) );
  AND2_X1 U1996 ( .A1(n121), .A2(n152), .ZN(n1904) );
  AND2_X1 U1997 ( .A1(n121), .A2(n148), .ZN(n1905) );
  AND2_X1 U1998 ( .A1(n121), .A2(n139), .ZN(n1906) );
  AND2_X1 U1999 ( .A1(n121), .A2(n139), .ZN(n1907) );
  AND2_X1 U2000 ( .A1(n121), .A2(n148), .ZN(n1908) );
  AND2_X1 U2001 ( .A1(n121), .A2(RST), .ZN(n1909) );
  AND2_X1 U2002 ( .A1(n121), .A2(n139), .ZN(n1910) );
  AND2_X1 U2003 ( .A1(n121), .A2(RST), .ZN(n1911) );
  AND2_X1 U2004 ( .A1(n75), .A2(RST), .ZN(n1912) );
  AND2_X1 U2005 ( .A1(n75), .A2(n153), .ZN(n1913) );
  AND2_X1 U2006 ( .A1(n75), .A2(RST), .ZN(n1914) );
  AND2_X1 U2007 ( .A1(n75), .A2(n153), .ZN(n1915) );
  AND2_X1 U2008 ( .A1(n75), .A2(n149), .ZN(n1916) );
  AND2_X1 U2009 ( .A1(n75), .A2(n152), .ZN(n1917) );
  AND2_X1 U2010 ( .A1(n75), .A2(n152), .ZN(n1918) );
  AND2_X1 U2011 ( .A1(n75), .A2(n150), .ZN(n1919) );
  AND2_X1 U2012 ( .A1(n75), .A2(n144), .ZN(n1920) );
  AND2_X1 U2013 ( .A1(n75), .A2(n143), .ZN(n1921) );
  AND2_X1 U2014 ( .A1(n75), .A2(n150), .ZN(n1922) );
  AND2_X1 U2015 ( .A1(n75), .A2(RST), .ZN(n1923) );
  AND2_X1 U2016 ( .A1(n75), .A2(RST), .ZN(n1924) );
  AND2_X1 U2017 ( .A1(n75), .A2(n137), .ZN(n1925) );
  AND2_X1 U2018 ( .A1(n75), .A2(RST), .ZN(n1926) );
  AND2_X1 U2019 ( .A1(n75), .A2(RST), .ZN(n1927) );
  AND2_X1 U2020 ( .A1(n75), .A2(n140), .ZN(n1928) );
  AND2_X1 U2021 ( .A1(n75), .A2(n142), .ZN(n1929) );
  AND2_X1 U2022 ( .A1(n75), .A2(n140), .ZN(n1930) );
  AND2_X1 U2023 ( .A1(n75), .A2(n138), .ZN(n1931) );
  AND2_X1 U2024 ( .A1(n75), .A2(RST), .ZN(n1932) );
  AND2_X1 U2025 ( .A1(n75), .A2(n146), .ZN(n1933) );
  AND2_X1 U2026 ( .A1(n133), .A2(n152), .ZN(n1934) );
  AND2_X1 U2027 ( .A1(n133), .A2(n146), .ZN(n1935) );
  AND2_X1 U2028 ( .A1(n133), .A2(n153), .ZN(n1936) );
  AND2_X1 U2029 ( .A1(n133), .A2(n147), .ZN(n1937) );
  AND2_X1 U2030 ( .A1(n133), .A2(n152), .ZN(n1938) );
  AND2_X1 U2031 ( .A1(n133), .A2(n143), .ZN(n1939) );
  AND2_X1 U2032 ( .A1(n133), .A2(n150), .ZN(n1940) );
  AND2_X1 U2033 ( .A1(n133), .A2(n147), .ZN(n1941) );
  AND2_X1 U2034 ( .A1(n133), .A2(RST), .ZN(n1942) );
  AND2_X1 U2035 ( .A1(n133), .A2(n141), .ZN(n1943) );
  AND2_X1 U2036 ( .A1(n133), .A2(n146), .ZN(n1944) );
  AND2_X1 U2037 ( .A1(n133), .A2(n140), .ZN(n1945) );
  AND2_X1 U2038 ( .A1(n133), .A2(RST), .ZN(n1946) );
  AND2_X1 U2039 ( .A1(n133), .A2(n137), .ZN(n1947) );
  AND2_X1 U2040 ( .A1(n133), .A2(n153), .ZN(n1948) );
  AND2_X1 U2041 ( .A1(n133), .A2(n155), .ZN(n1949) );
  AND2_X1 U2042 ( .A1(n133), .A2(n142), .ZN(n1950) );
  AND2_X1 U2043 ( .A1(n133), .A2(n140), .ZN(n1951) );
  AND2_X1 U2044 ( .A1(n133), .A2(n138), .ZN(n1952) );
  AND2_X1 U2045 ( .A1(n133), .A2(n151), .ZN(n1953) );
  AND2_X1 U2046 ( .A1(n133), .A2(RST), .ZN(n1954) );
  AND2_X1 U2047 ( .A1(n133), .A2(RST), .ZN(n1955) );
  AND2_X1 U2048 ( .A1(n135), .A2(n146), .ZN(n1956) );
  AND2_X1 U2049 ( .A1(n135), .A2(n144), .ZN(n1957) );
  AND2_X1 U2050 ( .A1(n135), .A2(n153), .ZN(n1958) );
  AND2_X1 U2051 ( .A1(n135), .A2(n148), .ZN(n1959) );
  AND2_X1 U2052 ( .A1(n135), .A2(n152), .ZN(n1960) );
  AND2_X1 U2053 ( .A1(n135), .A2(n153), .ZN(n1961) );
  AND2_X1 U2054 ( .A1(DATAIN[31]), .A2(n149), .ZN(n1962) );
  AND2_X1 U2055 ( .A1(DATAIN[31]), .A2(n144), .ZN(n1963) );
  AND2_X1 U2056 ( .A1(DATAIN[31]), .A2(n153), .ZN(n1964) );
  AND2_X1 U2057 ( .A1(DATAIN[31]), .A2(n153), .ZN(n1965) );
  AND2_X1 U2058 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1966) );
  AND2_X1 U2059 ( .A1(DATAIN[31]), .A2(n152), .ZN(n1967) );
  AND2_X1 U2060 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1968) );
  AND2_X1 U2061 ( .A1(DATAIN[31]), .A2(n150), .ZN(n1969) );
  AND2_X1 U2062 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1970) );
  AND2_X1 U2063 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1971) );
  AND2_X1 U2064 ( .A1(DATAIN[31]), .A2(n148), .ZN(n1972) );
  AND2_X1 U2065 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1973) );
  AND2_X1 U2066 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1974) );
  AND2_X1 U2067 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1975) );
  AND2_X1 U2068 ( .A1(DATAIN[31]), .A2(n145), .ZN(n1976) );
  AND2_X1 U2069 ( .A1(DATAIN[31]), .A2(n144), .ZN(n1977) );
  AND2_X1 U2070 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1978) );
  AND2_X1 U2071 ( .A1(DATAIN[31]), .A2(n143), .ZN(n1979) );
  AND2_X1 U2072 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1980) );
  AND2_X1 U2073 ( .A1(DATAIN[31]), .A2(n137), .ZN(n1981) );
  AND2_X1 U2074 ( .A1(DATAIN[31]), .A2(n139), .ZN(n1982) );
  AND2_X1 U2075 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1983) );
  AND2_X1 U2076 ( .A1(DATAIN[31]), .A2(n142), .ZN(n1984) );
  AND2_X1 U2077 ( .A1(DATAIN[31]), .A2(n138), .ZN(n1985) );
  AND2_X1 U2078 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1986) );
  AND2_X1 U2079 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1987) );
  AND2_X1 U2080 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1988) );
  AND2_X1 U2081 ( .A1(DATAIN[31]), .A2(n142), .ZN(n1989) );
  AND2_X1 U2082 ( .A1(DATAIN[31]), .A2(n140), .ZN(n1990) );
  AND2_X1 U2083 ( .A1(DATAIN[31]), .A2(n138), .ZN(n1991) );
  AND2_X1 U2084 ( .A1(DATAIN[31]), .A2(RST), .ZN(n1992) );
  AND2_X1 U2085 ( .A1(n135), .A2(n150), .ZN(n1993) );
  AND2_X1 U2086 ( .A1(n135), .A2(n148), .ZN(n1994) );
  AND2_X1 U2087 ( .A1(n135), .A2(RST), .ZN(n1995) );
  AND2_X1 U2088 ( .A1(n135), .A2(n142), .ZN(n1996) );
  AND2_X1 U2089 ( .A1(n135), .A2(n138), .ZN(n1997) );
  AND2_X1 U2090 ( .A1(n135), .A2(n137), .ZN(n1998) );
  AND2_X1 U2091 ( .A1(n135), .A2(RST), .ZN(n1999) );
  AND2_X1 U2092 ( .A1(n135), .A2(n142), .ZN(n2000) );
  AND2_X1 U2093 ( .A1(n135), .A2(n138), .ZN(n2001) );
  AND2_X1 U2094 ( .A1(n135), .A2(n144), .ZN(n2002) );
  AND2_X1 U2095 ( .A1(DATAIN[6]), .A2(n155), .ZN(n2003) );
  AND2_X1 U2096 ( .A1(DATAIN[6]), .A2(RST), .ZN(n2004) );
  AND2_X1 U2097 ( .A1(DATAIN[6]), .A2(n154), .ZN(n2005) );
  AND2_X1 U2098 ( .A1(DATAIN[6]), .A2(RST), .ZN(n2006) );
  AND2_X1 U2099 ( .A1(DATAIN[6]), .A2(RST), .ZN(n2007) );
  AND2_X1 U2100 ( .A1(DATAIN[6]), .A2(n155), .ZN(n2008) );
  AND2_X1 U2101 ( .A1(DATAIN[6]), .A2(n151), .ZN(n2009) );
  AND2_X1 U2102 ( .A1(DATAIN[6]), .A2(n151), .ZN(n2010) );
  AND2_X1 U2103 ( .A1(DATAIN[6]), .A2(RST), .ZN(n2011) );
  AND2_X1 U2104 ( .A1(DATAIN[6]), .A2(n149), .ZN(n2012) );
  AND2_X1 U2105 ( .A1(DATAIN[6]), .A2(n147), .ZN(n2013) );
  AND2_X1 U2106 ( .A1(DATAIN[6]), .A2(RST), .ZN(n2014) );
  AND2_X1 U2107 ( .A1(DATAIN[6]), .A2(n151), .ZN(n2015) );
  AND2_X1 U2108 ( .A1(DATAIN[6]), .A2(n146), .ZN(n2016) );
  AND2_X1 U2109 ( .A1(DATAIN[6]), .A2(RST), .ZN(n2017) );
  AND2_X1 U2110 ( .A1(DATAIN[6]), .A2(n151), .ZN(n2018) );
  AND2_X1 U2111 ( .A1(DATAIN[6]), .A2(n147), .ZN(n2019) );
  AND2_X1 U2112 ( .A1(DATAIN[6]), .A2(n149), .ZN(n2020) );
  AND2_X1 U2113 ( .A1(DATAIN[6]), .A2(n147), .ZN(n2021) );
  AND2_X1 U2114 ( .A1(DATAIN[6]), .A2(n140), .ZN(n2022) );
  AND2_X1 U2115 ( .A1(DATAIN[6]), .A2(RST), .ZN(n2023) );
  AND2_X1 U2116 ( .A1(DATAIN[6]), .A2(n140), .ZN(n2024) );
  AND2_X1 U2117 ( .A1(DATAIN[6]), .A2(n141), .ZN(n2025) );
  AND2_X1 U2118 ( .A1(DATAIN[6]), .A2(n142), .ZN(n2026) );
  AND2_X1 U2119 ( .A1(DATAIN[6]), .A2(n139), .ZN(n2027) );
  AND2_X1 U2120 ( .A1(DATAIN[6]), .A2(n142), .ZN(n2028) );
  AND2_X1 U2121 ( .A1(DATAIN[6]), .A2(n141), .ZN(n2029) );
  AND2_X1 U2122 ( .A1(DATAIN[6]), .A2(n139), .ZN(n2030) );
  AND2_X1 U2123 ( .A1(DATAIN[6]), .A2(n137), .ZN(n2031) );
  AND2_X1 U2124 ( .A1(DATAIN[6]), .A2(n147), .ZN(n2032) );
  AND2_X1 U2125 ( .A1(DATAIN[6]), .A2(n139), .ZN(n2033) );
  AND2_X1 U2126 ( .A1(n83), .A2(RST), .ZN(n2034) );
  AND2_X1 U2127 ( .A1(n83), .A2(RST), .ZN(n2035) );
  AND2_X1 U2128 ( .A1(n83), .A2(n143), .ZN(n2036) );
  AND2_X1 U2129 ( .A1(n83), .A2(n153), .ZN(n2037) );
  AND2_X1 U2130 ( .A1(n83), .A2(RST), .ZN(n2038) );
  AND2_X1 U2131 ( .A1(n83), .A2(n152), .ZN(n2039) );
  AND2_X1 U2132 ( .A1(n83), .A2(RST), .ZN(n2040) );
  AND2_X1 U2133 ( .A1(n83), .A2(n150), .ZN(n2041) );
  AND2_X1 U2134 ( .A1(n83), .A2(n144), .ZN(n2042) );
  AND2_X1 U2135 ( .A1(n83), .A2(n143), .ZN(n2043) );
  AND2_X1 U2136 ( .A1(n83), .A2(RST), .ZN(n2044) );
  AND2_X1 U2137 ( .A1(n83), .A2(RST), .ZN(n2045) );
  AND2_X1 U2138 ( .A1(n83), .A2(RST), .ZN(n2046) );
  AND2_X1 U2139 ( .A1(n83), .A2(n141), .ZN(n2047) );
  AND2_X1 U2140 ( .A1(n83), .A2(n137), .ZN(n2048) );
  AND2_X1 U2141 ( .A1(n83), .A2(n144), .ZN(n2049) );
  AND2_X1 U2142 ( .A1(n83), .A2(n142), .ZN(n2050) );
  AND2_X1 U2143 ( .A1(n83), .A2(n142), .ZN(n2051) );
  AND2_X1 U2144 ( .A1(n83), .A2(n140), .ZN(n2052) );
  AND2_X1 U2145 ( .A1(n83), .A2(n138), .ZN(n2053) );
  AND2_X1 U2146 ( .A1(n83), .A2(n145), .ZN(n2054) );
  AND2_X1 U2147 ( .A1(n83), .A2(n143), .ZN(n2055) );
  AND2_X1 U2148 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2056) );
  AND2_X1 U2149 ( .A1(DATAIN[28]), .A2(n150), .ZN(n2057) );
  AND2_X1 U2150 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2058) );
  AND2_X1 U2151 ( .A1(DATAIN[28]), .A2(n153), .ZN(n2059) );
  AND2_X1 U2152 ( .A1(DATAIN[28]), .A2(n150), .ZN(n2060) );
  AND2_X1 U2153 ( .A1(DATAIN[28]), .A2(n152), .ZN(n2061) );
  AND2_X1 U2154 ( .A1(DATAIN[28]), .A2(n145), .ZN(n2062) );
  AND2_X1 U2155 ( .A1(DATAIN[28]), .A2(n150), .ZN(n2063) );
  AND2_X1 U2156 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2064) );
  AND2_X1 U2157 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2065) );
  AND2_X1 U2158 ( .A1(DATAIN[28]), .A2(n148), .ZN(n2066) );
  AND2_X1 U2159 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2067) );
  AND2_X1 U2160 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2068) );
  AND2_X1 U2161 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2069) );
  AND2_X1 U2162 ( .A1(DATAIN[28]), .A2(n145), .ZN(n2070) );
  AND2_X1 U2163 ( .A1(DATAIN[28]), .A2(n144), .ZN(n2071) );
  AND2_X1 U2164 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2072) );
  AND2_X1 U2165 ( .A1(DATAIN[28]), .A2(n143), .ZN(n2073) );
  AND2_X1 U2166 ( .A1(DATAIN[28]), .A2(n140), .ZN(n2074) );
  AND2_X1 U2167 ( .A1(DATAIN[28]), .A2(n141), .ZN(n2075) );
  AND2_X1 U2168 ( .A1(DATAIN[28]), .A2(n146), .ZN(n2076) );
  AND2_X1 U2169 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2077) );
  AND2_X1 U2170 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2078) );
  AND2_X1 U2171 ( .A1(DATAIN[28]), .A2(n139), .ZN(n2079) );
  AND2_X1 U2172 ( .A1(DATAIN[28]), .A2(n139), .ZN(n2080) );
  AND2_X1 U2173 ( .A1(DATAIN[28]), .A2(n155), .ZN(n2081) );
  AND2_X1 U2174 ( .A1(DATAIN[28]), .A2(n154), .ZN(n2082) );
  AND2_X1 U2175 ( .A1(DATAIN[28]), .A2(n142), .ZN(n2083) );
  AND2_X1 U2176 ( .A1(DATAIN[28]), .A2(n140), .ZN(n2084) );
  AND2_X1 U2177 ( .A1(DATAIN[28]), .A2(n138), .ZN(n2085) );
  AND2_X1 U2178 ( .A1(DATAIN[28]), .A2(n147), .ZN(n2086) );
  AND2_X1 U2179 ( .A1(n1636), .A2(n155), .ZN(n2087) );
  AND2_X1 U2180 ( .A1(n1636), .A2(RST), .ZN(n2088) );
  AND2_X1 U2181 ( .A1(n1636), .A2(n154), .ZN(n2089) );
  AND2_X1 U2182 ( .A1(n1636), .A2(n148), .ZN(n2090) );
  AND2_X1 U2183 ( .A1(n1636), .A2(RST), .ZN(n2091) );
  AND2_X1 U2184 ( .A1(n1636), .A2(RST), .ZN(n2092) );
  AND2_X1 U2185 ( .A1(n1636), .A2(n151), .ZN(n2093) );
  AND2_X1 U2186 ( .A1(n1636), .A2(RST), .ZN(n2094) );
  AND2_X1 U2187 ( .A1(n1636), .A2(n149), .ZN(n2095) );
  AND2_X1 U2188 ( .A1(n1636), .A2(n145), .ZN(n2096) );
  AND2_X1 U2189 ( .A1(n1636), .A2(RST), .ZN(n2097) );
  AND2_X1 U2190 ( .A1(n1636), .A2(RST), .ZN(n2098) );
  AND2_X1 U2191 ( .A1(n1636), .A2(RST), .ZN(n2099) );
  AND2_X1 U2192 ( .A1(n1636), .A2(n137), .ZN(n2100) );
  AND2_X1 U2193 ( .A1(n1636), .A2(n140), .ZN(n2101) );
  AND2_X1 U2194 ( .A1(n1636), .A2(n137), .ZN(n2102) );
  AND2_X1 U2195 ( .A1(n1636), .A2(RST), .ZN(n2103) );
  AND2_X1 U2196 ( .A1(n1636), .A2(n141), .ZN(n2104) );
  AND2_X1 U2197 ( .A1(n1636), .A2(n139), .ZN(n2105) );
  AND2_X1 U2198 ( .A1(n1636), .A2(n137), .ZN(n2106) );
  AND2_X1 U2199 ( .A1(n1636), .A2(RST), .ZN(n2107) );
  AND2_X1 U2200 ( .A1(n1636), .A2(RST), .ZN(n2108) );
  AND2_X1 U2201 ( .A1(n97), .A2(n155), .ZN(n2109) );
  AND2_X1 U2202 ( .A1(n97), .A2(RST), .ZN(n2110) );
  AND2_X1 U2203 ( .A1(n97), .A2(n154), .ZN(n2111) );
  AND2_X1 U2204 ( .A1(n97), .A2(n154), .ZN(n2112) );
  AND2_X1 U2205 ( .A1(n97), .A2(RST), .ZN(n2113) );
  AND2_X1 U2206 ( .A1(n97), .A2(RST), .ZN(n2114) );
  AND2_X1 U2207 ( .A1(n97), .A2(n151), .ZN(n2115) );
  AND2_X1 U2208 ( .A1(n97), .A2(n144), .ZN(n2116) );
  AND2_X1 U2209 ( .A1(n97), .A2(RST), .ZN(n2117) );
  AND2_X1 U2210 ( .A1(n97), .A2(RST), .ZN(n2118) );
  AND2_X1 U2211 ( .A1(n97), .A2(RST), .ZN(n2119) );
  AND2_X1 U2212 ( .A1(n97), .A2(RST), .ZN(n2120) );
  AND2_X1 U2213 ( .A1(n97), .A2(n140), .ZN(n2121) );
  AND2_X1 U2214 ( .A1(n97), .A2(n139), .ZN(n2122) );
  AND2_X1 U2215 ( .A1(n97), .A2(n149), .ZN(n2123) );
  AND2_X1 U2216 ( .A1(n97), .A2(n155), .ZN(n2124) );
  AND2_X1 U2217 ( .A1(n97), .A2(RST), .ZN(n2125) );
  AND2_X1 U2218 ( .A1(n97), .A2(n141), .ZN(n2126) );
  AND2_X1 U2219 ( .A1(n97), .A2(n139), .ZN(n2127) );
  AND2_X1 U2220 ( .A1(n97), .A2(n137), .ZN(n2128) );
  AND2_X1 U2221 ( .A1(n97), .A2(n153), .ZN(n2129) );
  AND2_X1 U2222 ( .A1(n97), .A2(RST), .ZN(n2130) );
  AND2_X1 U2223 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2131) );
  AND2_X1 U2224 ( .A1(DATAIN[2]), .A2(n148), .ZN(n2132) );
  AND2_X1 U2225 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2133) );
  AND2_X1 U2226 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2134) );
  AND2_X1 U2227 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2135) );
  AND2_X1 U2228 ( .A1(DATAIN[2]), .A2(n145), .ZN(n2136) );
  AND2_X1 U2229 ( .A1(DATAIN[2]), .A2(n144), .ZN(n2137) );
  AND2_X1 U2230 ( .A1(DATAIN[2]), .A2(n143), .ZN(n2138) );
  AND2_X1 U2231 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2139) );
  AND2_X1 U2232 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2140) );
  AND2_X1 U2233 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2141) );
  AND2_X1 U2234 ( .A1(DATAIN[2]), .A2(n145), .ZN(n2142) );
  AND2_X1 U2235 ( .A1(DATAIN[2]), .A2(n153), .ZN(n2143) );
  AND2_X1 U2236 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2144) );
  AND2_X1 U2237 ( .A1(DATAIN[2]), .A2(n152), .ZN(n2145) );
  AND2_X1 U2238 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2146) );
  AND2_X1 U2239 ( .A1(DATAIN[2]), .A2(n150), .ZN(n2147) );
  AND2_X1 U2240 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2148) );
  AND2_X1 U2241 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2149) );
  AND2_X1 U2242 ( .A1(DATAIN[2]), .A2(n140), .ZN(n2150) );
  AND2_X1 U2243 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2151) );
  AND2_X1 U2244 ( .A1(DATAIN[2]), .A2(n139), .ZN(n2152) );
  AND2_X1 U2245 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2153) );
  AND2_X1 U2246 ( .A1(DATAIN[2]), .A2(n152), .ZN(n2154) );
  AND2_X1 U2247 ( .A1(DATAIN[2]), .A2(n153), .ZN(n2155) );
  AND2_X1 U2248 ( .A1(DATAIN[2]), .A2(n147), .ZN(n2156) );
  AND2_X1 U2249 ( .A1(DATAIN[2]), .A2(n142), .ZN(n2157) );
  AND2_X1 U2250 ( .A1(DATAIN[2]), .A2(n140), .ZN(n2158) );
  AND2_X1 U2251 ( .A1(DATAIN[2]), .A2(n138), .ZN(n2159) );
  AND2_X1 U2252 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2160) );
  AND2_X1 U2253 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2161) );
  AND2_X1 U2254 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2162) );
  AND2_X1 U2255 ( .A1(n129), .A2(RST), .ZN(n2163) );
  AND2_X1 U2256 ( .A1(n129), .A2(RST), .ZN(n2164) );
  AND2_X1 U2257 ( .A1(n129), .A2(n153), .ZN(n2165) );
  AND2_X1 U2258 ( .A1(n129), .A2(n145), .ZN(n2166) );
  AND2_X1 U2259 ( .A1(n129), .A2(n152), .ZN(n2167) );
  AND2_X1 U2260 ( .A1(n129), .A2(n155), .ZN(n2168) );
  AND2_X1 U2261 ( .A1(n129), .A2(n150), .ZN(n2169) );
  AND2_X1 U2262 ( .A1(n129), .A2(RST), .ZN(n2170) );
  AND2_X1 U2263 ( .A1(n129), .A2(RST), .ZN(n2171) );
  AND2_X1 U2264 ( .A1(n129), .A2(n139), .ZN(n2172) );
  AND2_X1 U2265 ( .A1(n129), .A2(n142), .ZN(n2173) );
  AND2_X1 U2266 ( .A1(n129), .A2(n146), .ZN(n2174) );
  AND2_X1 U2267 ( .A1(n129), .A2(n138), .ZN(n2175) );
  AND2_X1 U2268 ( .A1(n129), .A2(RST), .ZN(n2176) );
  AND2_X1 U2269 ( .A1(n129), .A2(RST), .ZN(n2177) );
  AND2_X1 U2270 ( .A1(n129), .A2(n141), .ZN(n2178) );
  AND2_X1 U2271 ( .A1(n129), .A2(RST), .ZN(n2179) );
  AND2_X1 U2272 ( .A1(n129), .A2(n142), .ZN(n2180) );
  AND2_X1 U2273 ( .A1(n129), .A2(n140), .ZN(n2181) );
  AND2_X1 U2274 ( .A1(n129), .A2(n138), .ZN(n2182) );
  AND2_X1 U2275 ( .A1(n129), .A2(RST), .ZN(n2183) );
  AND2_X1 U2276 ( .A1(n129), .A2(n150), .ZN(n2184) );
  AND2_X1 U2277 ( .A1(DATAIN[20]), .A2(n155), .ZN(n2185) );
  AND2_X1 U2278 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2186) );
  AND2_X1 U2279 ( .A1(DATAIN[20]), .A2(n154), .ZN(n2187) );
  AND2_X1 U2280 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2188) );
  AND2_X1 U2281 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2189) );
  AND2_X1 U2282 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2190) );
  AND2_X1 U2283 ( .A1(DATAIN[20]), .A2(n151), .ZN(n2191) );
  AND2_X1 U2284 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2192) );
  AND2_X1 U2285 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2193) );
  AND2_X1 U2286 ( .A1(DATAIN[20]), .A2(n149), .ZN(n2194) );
  AND2_X1 U2287 ( .A1(DATAIN[20]), .A2(n147), .ZN(n2195) );
  AND2_X1 U2288 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2196) );
  AND2_X1 U2289 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2197) );
  AND2_X1 U2290 ( .A1(DATAIN[20]), .A2(n146), .ZN(n2198) );
  AND2_X1 U2291 ( .A1(DATAIN[20]), .A2(n146), .ZN(n2199) );
  AND2_X1 U2292 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2200) );
  AND2_X1 U2293 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2201) );
  AND2_X1 U2294 ( .A1(DATAIN[20]), .A2(n153), .ZN(n2202) );
  AND2_X1 U2295 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2203) );
  AND2_X1 U2296 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2204) );
  AND2_X1 U2297 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2205) );
  AND2_X1 U2298 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2206) );
  AND2_X1 U2299 ( .A1(DATAIN[20]), .A2(n139), .ZN(n2207) );
  AND2_X1 U2300 ( .A1(DATAIN[20]), .A2(n138), .ZN(n2208) );
  AND2_X1 U2301 ( .A1(DATAIN[20]), .A2(n138), .ZN(n2209) );
  AND2_X1 U2302 ( .A1(DATAIN[20]), .A2(n147), .ZN(n2210) );
  AND2_X1 U2303 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2211) );
  AND2_X1 U2304 ( .A1(DATAIN[20]), .A2(n141), .ZN(n2212) );
  AND2_X1 U2305 ( .A1(DATAIN[20]), .A2(n139), .ZN(n2213) );
  AND2_X1 U2306 ( .A1(DATAIN[20]), .A2(n137), .ZN(n2214) );
  AND2_X1 U2307 ( .A1(DATAIN[20]), .A2(n144), .ZN(n2215) );
  AND2_X1 U2308 ( .A1(DATAIN[20]), .A2(n149), .ZN(n2216) );
  AND2_X1 U2309 ( .A1(DATAIN[25]), .A2(n153), .ZN(n2217) );
  AND2_X1 U2310 ( .A1(DATAIN[25]), .A2(n154), .ZN(n2218) );
  AND2_X1 U2311 ( .A1(DATAIN[25]), .A2(n152), .ZN(n2219) );
  AND2_X1 U2312 ( .A1(DATAIN[25]), .A2(n153), .ZN(n2220) );
  AND2_X1 U2313 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2221) );
  AND2_X1 U2314 ( .A1(DATAIN[25]), .A2(n152), .ZN(n2222) );
  AND2_X1 U2315 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2223) );
  AND2_X1 U2316 ( .A1(DATAIN[25]), .A2(n150), .ZN(n2224) );
  AND2_X1 U2317 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2225) );
  AND2_X1 U2318 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2226) );
  AND2_X1 U2319 ( .A1(DATAIN[25]), .A2(n148), .ZN(n2227) );
  AND2_X1 U2320 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2228) );
  AND2_X1 U2321 ( .A1(DATAIN[25]), .A2(n155), .ZN(n2229) );
  AND2_X1 U2322 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2230) );
  AND2_X1 U2323 ( .A1(DATAIN[25]), .A2(n145), .ZN(n2231) );
  AND2_X1 U2324 ( .A1(DATAIN[25]), .A2(n144), .ZN(n2232) );
  AND2_X1 U2325 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2233) );
  AND2_X1 U2326 ( .A1(DATAIN[25]), .A2(n143), .ZN(n2234) );
  AND2_X1 U2327 ( .A1(DATAIN[25]), .A2(n139), .ZN(n2235) );
  AND2_X1 U2328 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2236) );
  AND2_X1 U2329 ( .A1(DATAIN[25]), .A2(n138), .ZN(n2237) );
  AND2_X1 U2330 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2238) );
  AND2_X1 U2331 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2239) );
  AND2_X1 U2332 ( .A1(DATAIN[25]), .A2(n142), .ZN(n2240) );
  AND2_X1 U2333 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2241) );
  AND2_X1 U2334 ( .A1(DATAIN[25]), .A2(n141), .ZN(n2242) );
  AND2_X1 U2335 ( .A1(DATAIN[25]), .A2(n137), .ZN(n2243) );
  AND2_X1 U2336 ( .A1(DATAIN[25]), .A2(n142), .ZN(n2244) );
  AND2_X1 U2337 ( .A1(DATAIN[25]), .A2(n140), .ZN(n2245) );
  AND2_X1 U2338 ( .A1(DATAIN[25]), .A2(n138), .ZN(n2246) );
  AND2_X1 U2339 ( .A1(DATAIN[25]), .A2(n154), .ZN(n2247) );
  AND2_X1 U2340 ( .A1(DATAIN[25]), .A2(n149), .ZN(n2248) );
  AND2_X1 U2341 ( .A1(n91), .A2(n143), .ZN(n2249) );
  AND2_X1 U2342 ( .A1(n91), .A2(n151), .ZN(n2250) );
  AND2_X1 U2343 ( .A1(n91), .A2(n147), .ZN(n2251) );
  AND2_X1 U2344 ( .A1(n91), .A2(n153), .ZN(n2252) );
  AND2_X1 U2345 ( .A1(n91), .A2(RST), .ZN(n2253) );
  AND2_X1 U2346 ( .A1(n91), .A2(n152), .ZN(n2254) );
  AND2_X1 U2347 ( .A1(n91), .A2(n149), .ZN(n2255) );
  AND2_X1 U2348 ( .A1(n91), .A2(n150), .ZN(n2256) );
  AND2_X1 U2349 ( .A1(n91), .A2(n144), .ZN(n2257) );
  AND2_X1 U2350 ( .A1(n91), .A2(n143), .ZN(n2258) );
  AND2_X1 U2351 ( .A1(n91), .A2(n146), .ZN(n2259) );
  AND2_X1 U2352 ( .A1(n91), .A2(RST), .ZN(n2260) );
  AND2_X1 U2353 ( .A1(n91), .A2(n137), .ZN(n2261) );
  AND2_X1 U2354 ( .A1(n91), .A2(RST), .ZN(n2262) );
  AND2_X1 U2355 ( .A1(n91), .A2(n142), .ZN(n2263) );
  AND2_X1 U2356 ( .A1(n91), .A2(n152), .ZN(n2264) );
  AND2_X1 U2357 ( .A1(n91), .A2(n141), .ZN(n2265) );
  AND2_X1 U2358 ( .A1(n91), .A2(n142), .ZN(n2266) );
  AND2_X1 U2359 ( .A1(n91), .A2(n140), .ZN(n2267) );
  AND2_X1 U2360 ( .A1(n91), .A2(n138), .ZN(n2268) );
  AND2_X1 U2361 ( .A1(n91), .A2(n152), .ZN(n2269) );
  AND2_X1 U2362 ( .A1(n91), .A2(RST), .ZN(n2270) );
  AND2_X1 U2363 ( .A1(n107), .A2(n155), .ZN(n2271) );
  AND2_X1 U2364 ( .A1(n107), .A2(RST), .ZN(n2272) );
  AND2_X1 U2365 ( .A1(n107), .A2(n154), .ZN(n2273) );
  AND2_X1 U2366 ( .A1(n107), .A2(n151), .ZN(n2274) );
  AND2_X1 U2367 ( .A1(n107), .A2(RST), .ZN(n2275) );
  AND2_X1 U2368 ( .A1(n107), .A2(n150), .ZN(n2276) );
  AND2_X1 U2369 ( .A1(n107), .A2(n151), .ZN(n2277) );
  AND2_X1 U2370 ( .A1(n107), .A2(RST), .ZN(n2278) );
  AND2_X1 U2371 ( .A1(n107), .A2(RST), .ZN(n2279) );
  AND2_X1 U2372 ( .A1(n107), .A2(n154), .ZN(n2280) );
  AND2_X1 U2373 ( .A1(n107), .A2(n141), .ZN(n2281) );
  AND2_X1 U2374 ( .A1(n107), .A2(n144), .ZN(n2282) );
  AND2_X1 U2375 ( .A1(n101), .A2(n155), .ZN(n2283) );
  AND2_X1 U2376 ( .A1(n101), .A2(RST), .ZN(n2284) );
  AND2_X1 U2377 ( .A1(n101), .A2(n154), .ZN(n2285) );
  AND2_X1 U2378 ( .A1(n101), .A2(RST), .ZN(n2286) );
  AND2_X1 U2379 ( .A1(n101), .A2(RST), .ZN(n2287) );
  AND2_X1 U2380 ( .A1(n101), .A2(n152), .ZN(n2288) );
  AND2_X1 U2381 ( .A1(n101), .A2(n151), .ZN(n2289) );
  AND2_X1 U2382 ( .A1(n101), .A2(n148), .ZN(n2290) );
  AND2_X1 U2383 ( .A1(n101), .A2(n146), .ZN(n2291) );
  AND2_X1 U2384 ( .A1(n101), .A2(RST), .ZN(n2292) );
  AND2_X1 U2385 ( .A1(n101), .A2(n138), .ZN(n2293) );
  AND2_X1 U2386 ( .A1(n101), .A2(RST), .ZN(n2294) );
  AND2_X1 U2387 ( .A1(n101), .A2(n142), .ZN(n2295) );
  AND2_X1 U2388 ( .A1(n101), .A2(n141), .ZN(n2296) );
  AND2_X1 U2389 ( .A1(n101), .A2(RST), .ZN(n2297) );
  AND2_X1 U2390 ( .A1(n101), .A2(RST), .ZN(n2298) );
  AND2_X1 U2391 ( .A1(n101), .A2(n147), .ZN(n2299) );
  AND2_X1 U2392 ( .A1(n101), .A2(n141), .ZN(n2300) );
  AND2_X1 U2393 ( .A1(n101), .A2(n139), .ZN(n2301) );
  AND2_X1 U2394 ( .A1(n101), .A2(n137), .ZN(n2302) );
  AND2_X1 U2395 ( .A1(n101), .A2(RST), .ZN(n2303) );
  AND2_X1 U2396 ( .A1(n101), .A2(n150), .ZN(n2304) );
  AND2_X1 U2397 ( .A1(n107), .A2(RST), .ZN(n2305) );
  AND2_X1 U2398 ( .A1(n107), .A2(RST), .ZN(n2306) );
  AND2_X1 U2399 ( .A1(n107), .A2(RST), .ZN(n2307) );
  AND2_X1 U2400 ( .A1(n107), .A2(RST), .ZN(n2308) );
  AND2_X1 U2401 ( .A1(n107), .A2(n155), .ZN(n2309) );
  AND2_X1 U2402 ( .A1(n107), .A2(n154), .ZN(n2310) );
  AND2_X1 U2403 ( .A1(n107), .A2(n141), .ZN(n2311) );
  AND2_X1 U2404 ( .A1(n107), .A2(n139), .ZN(n2312) );
  AND2_X1 U2405 ( .A1(n107), .A2(n137), .ZN(n2313) );
  AND2_X1 U2406 ( .A1(n107), .A2(n148), .ZN(n2314) );
  AND2_X1 U2407 ( .A1(n77), .A2(n149), .ZN(n2315) );
  AND2_X1 U2408 ( .A1(n77), .A2(RST), .ZN(n2316) );
  AND2_X1 U2409 ( .A1(n77), .A2(n150), .ZN(n2317) );
  AND2_X1 U2410 ( .A1(n77), .A2(n153), .ZN(n2318) );
  AND2_X1 U2411 ( .A1(n77), .A2(RST), .ZN(n2319) );
  AND2_X1 U2412 ( .A1(n77), .A2(n152), .ZN(n2320) );
  AND2_X1 U2413 ( .A1(n77), .A2(n151), .ZN(n2321) );
  AND2_X1 U2414 ( .A1(n77), .A2(n150), .ZN(n2322) );
  AND2_X1 U2415 ( .A1(n77), .A2(n144), .ZN(n2323) );
  AND2_X1 U2416 ( .A1(n77), .A2(n143), .ZN(n2324) );
  AND2_X1 U2417 ( .A1(n77), .A2(RST), .ZN(n2325) );
  AND2_X1 U2418 ( .A1(n77), .A2(RST), .ZN(n2326) );
  AND2_X1 U2419 ( .A1(n77), .A2(RST), .ZN(n2327) );
  AND2_X1 U2420 ( .A1(n77), .A2(n138), .ZN(n2328) );
  AND2_X1 U2421 ( .A1(n77), .A2(RST), .ZN(n2329) );
  AND2_X1 U2422 ( .A1(n77), .A2(RST), .ZN(n2330) );
  AND2_X1 U2423 ( .A1(n77), .A2(n147), .ZN(n2331) );
  AND2_X1 U2424 ( .A1(n77), .A2(n142), .ZN(n2332) );
  AND2_X1 U2425 ( .A1(n77), .A2(n140), .ZN(n2333) );
  AND2_X1 U2426 ( .A1(n77), .A2(n138), .ZN(n2334) );
  AND2_X1 U2427 ( .A1(n77), .A2(RST), .ZN(n2335) );
  AND2_X1 U2428 ( .A1(n77), .A2(RST), .ZN(n2336) );
  AND2_X1 U2429 ( .A1(n125), .A2(n155), .ZN(n2337) );
  AND2_X1 U2430 ( .A1(n125), .A2(RST), .ZN(n2338) );
  AND2_X1 U2431 ( .A1(n125), .A2(n154), .ZN(n2339) );
  AND2_X1 U2432 ( .A1(n125), .A2(n154), .ZN(n2340) );
  AND2_X1 U2433 ( .A1(n125), .A2(RST), .ZN(n2341) );
  AND2_X1 U2434 ( .A1(n125), .A2(RST), .ZN(n2342) );
  AND2_X1 U2435 ( .A1(n125), .A2(n151), .ZN(n2343) );
  AND2_X1 U2436 ( .A1(n125), .A2(n145), .ZN(n2344) );
  AND2_X1 U2437 ( .A1(n125), .A2(n145), .ZN(n2345) );
  AND2_X1 U2438 ( .A1(n125), .A2(RST), .ZN(n2346) );
  AND2_X1 U2439 ( .A1(n125), .A2(RST), .ZN(n2347) );
  AND2_X1 U2440 ( .A1(n125), .A2(n141), .ZN(n2348) );
  AND2_X1 U2441 ( .A1(n125), .A2(n137), .ZN(n2349) );
  AND2_X1 U2442 ( .A1(n125), .A2(n141), .ZN(n2350) );
  AND2_X1 U2443 ( .A1(n125), .A2(n142), .ZN(n2351) );
  AND2_X1 U2444 ( .A1(n125), .A2(n139), .ZN(n2352) );
  AND2_X1 U2445 ( .A1(n125), .A2(n137), .ZN(n2353) );
  AND2_X1 U2446 ( .A1(n125), .A2(n141), .ZN(n2354) );
  AND2_X1 U2447 ( .A1(n125), .A2(n139), .ZN(n2355) );
  AND2_X1 U2448 ( .A1(n125), .A2(n137), .ZN(n2356) );
  AND2_X1 U2449 ( .A1(n125), .A2(n155), .ZN(n2357) );
  AND2_X1 U2450 ( .A1(n125), .A2(n151), .ZN(n2358) );
  AND2_X1 U2451 ( .A1(n109), .A2(n155), .ZN(n2359) );
  AND2_X1 U2452 ( .A1(n109), .A2(RST), .ZN(n2360) );
  AND2_X1 U2453 ( .A1(n109), .A2(n154), .ZN(n2361) );
  AND2_X1 U2454 ( .A1(n109), .A2(n145), .ZN(n2362) );
  AND2_X1 U2455 ( .A1(n109), .A2(RST), .ZN(n2363) );
  AND2_X1 U2456 ( .A1(n109), .A2(n146), .ZN(n2364) );
  AND2_X1 U2457 ( .A1(n109), .A2(n151), .ZN(n2365) );
  AND2_X1 U2458 ( .A1(n109), .A2(n154), .ZN(n2366) );
  AND2_X1 U2459 ( .A1(n109), .A2(n150), .ZN(n2367) );
  AND2_X1 U2460 ( .A1(n109), .A2(n143), .ZN(n2368) );
  AND2_X1 U2461 ( .A1(n109), .A2(n142), .ZN(n2369) );
  AND2_X1 U2462 ( .A1(n109), .A2(RST), .ZN(n2370) );
  AND2_X1 U2463 ( .A1(n109), .A2(RST), .ZN(n2371) );
  AND2_X1 U2464 ( .A1(n109), .A2(RST), .ZN(n2372) );
  AND2_X1 U2465 ( .A1(n109), .A2(RST), .ZN(n2373) );
  AND2_X1 U2466 ( .A1(n109), .A2(n143), .ZN(n2374) );
  AND2_X1 U2467 ( .A1(n109), .A2(n143), .ZN(n2375) );
  AND2_X1 U2468 ( .A1(n109), .A2(n141), .ZN(n2376) );
  AND2_X1 U2469 ( .A1(n109), .A2(n139), .ZN(n2377) );
  AND2_X1 U2470 ( .A1(n109), .A2(n137), .ZN(n2378) );
  AND2_X1 U2471 ( .A1(n109), .A2(RST), .ZN(n2379) );
  AND2_X1 U2472 ( .A1(n109), .A2(n153), .ZN(n2380) );
  AND2_X1 U2473 ( .A1(n87), .A2(n150), .ZN(n2381) );
  AND2_X1 U2474 ( .A1(n87), .A2(n143), .ZN(n2382) );
  AND2_X1 U2475 ( .A1(n87), .A2(n151), .ZN(n2383) );
  AND2_X1 U2476 ( .A1(n87), .A2(n153), .ZN(n2384) );
  AND2_X1 U2477 ( .A1(n87), .A2(RST), .ZN(n2385) );
  AND2_X1 U2478 ( .A1(n87), .A2(n152), .ZN(n2386) );
  AND2_X1 U2479 ( .A1(n87), .A2(n147), .ZN(n2387) );
  AND2_X1 U2480 ( .A1(n87), .A2(n150), .ZN(n2388) );
  AND2_X1 U2481 ( .A1(n87), .A2(n144), .ZN(n2389) );
  AND2_X1 U2482 ( .A1(n87), .A2(n143), .ZN(n2390) );
  AND2_X1 U2483 ( .A1(n87), .A2(n146), .ZN(n2391) );
  AND2_X1 U2484 ( .A1(n87), .A2(RST), .ZN(n2392) );
  AND2_X1 U2485 ( .A1(n87), .A2(RST), .ZN(n2393) );
  AND2_X1 U2486 ( .A1(n87), .A2(n137), .ZN(n2394) );
  AND2_X1 U2487 ( .A1(n87), .A2(RST), .ZN(n2395) );
  AND2_X1 U2488 ( .A1(n87), .A2(n139), .ZN(n2396) );
  AND2_X1 U2489 ( .A1(n87), .A2(n140), .ZN(n2397) );
  AND2_X1 U2490 ( .A1(n87), .A2(n142), .ZN(n2398) );
  AND2_X1 U2491 ( .A1(n87), .A2(n140), .ZN(n2399) );
  AND2_X1 U2492 ( .A1(n87), .A2(n138), .ZN(n2400) );
  AND2_X1 U2493 ( .A1(n87), .A2(n143), .ZN(n2401) );
  AND2_X1 U2494 ( .A1(n87), .A2(n149), .ZN(n2402) );
  AND2_X1 U2495 ( .A1(n93), .A2(n152), .ZN(n2403) );
  AND2_X1 U2496 ( .A1(n93), .A2(n145), .ZN(n2404) );
  AND2_X1 U2497 ( .A1(n93), .A2(n148), .ZN(n2405) );
  AND2_X1 U2498 ( .A1(n93), .A2(n153), .ZN(n2406) );
  AND2_X1 U2499 ( .A1(n93), .A2(n150), .ZN(n2407) );
  AND2_X1 U2500 ( .A1(n93), .A2(n152), .ZN(n2408) );
  AND2_X1 U2501 ( .A1(n93), .A2(RST), .ZN(n2409) );
  AND2_X1 U2502 ( .A1(n93), .A2(n150), .ZN(n2410) );
  AND2_X1 U2503 ( .A1(n93), .A2(n144), .ZN(n2411) );
  AND2_X1 U2504 ( .A1(n93), .A2(n143), .ZN(n2412) );
  AND2_X1 U2505 ( .A1(n93), .A2(RST), .ZN(n2413) );
  AND2_X1 U2506 ( .A1(n93), .A2(RST), .ZN(n2414) );
  AND2_X1 U2507 ( .A1(n93), .A2(n138), .ZN(n2415) );
  AND2_X1 U2508 ( .A1(n93), .A2(RST), .ZN(n2416) );
  AND2_X1 U2509 ( .A1(n93), .A2(n140), .ZN(n2417) );
  AND2_X1 U2510 ( .A1(n93), .A2(n140), .ZN(n2418) );
  AND2_X1 U2511 ( .A1(n93), .A2(n139), .ZN(n2419) );
  AND2_X1 U2512 ( .A1(n93), .A2(n142), .ZN(n2420) );
  AND2_X1 U2513 ( .A1(n93), .A2(n140), .ZN(n2421) );
  AND2_X1 U2514 ( .A1(n93), .A2(n138), .ZN(n2422) );
  AND2_X1 U2515 ( .A1(n93), .A2(RST), .ZN(n2423) );
  AND2_X1 U2516 ( .A1(n93), .A2(RST), .ZN(n2424) );
  AND2_X1 U2517 ( .A1(n81), .A2(RST), .ZN(n2425) );
  AND2_X1 U2518 ( .A1(n81), .A2(RST), .ZN(n2426) );
  AND2_X1 U2519 ( .A1(n81), .A2(n154), .ZN(n2427) );
  AND2_X1 U2520 ( .A1(n81), .A2(n153), .ZN(n2428) );
  AND2_X1 U2521 ( .A1(n81), .A2(n155), .ZN(n2429) );
  AND2_X1 U2522 ( .A1(n81), .A2(n152), .ZN(n2430) );
  AND2_X1 U2523 ( .A1(n81), .A2(n146), .ZN(n2431) );
  AND2_X1 U2524 ( .A1(n81), .A2(n150), .ZN(n2432) );
  AND2_X1 U2525 ( .A1(n81), .A2(n144), .ZN(n2433) );
  AND2_X1 U2526 ( .A1(n81), .A2(n143), .ZN(n2434) );
  AND2_X1 U2527 ( .A1(n81), .A2(n149), .ZN(n2435) );
  AND2_X1 U2528 ( .A1(n81), .A2(RST), .ZN(n2436) );
  AND2_X1 U2529 ( .A1(n81), .A2(RST), .ZN(n2437) );
  AND2_X1 U2530 ( .A1(n81), .A2(n140), .ZN(n2438) );
  AND2_X1 U2531 ( .A1(n81), .A2(RST), .ZN(n2439) );
  AND2_X1 U2532 ( .A1(n81), .A2(RST), .ZN(n2440) );
  AND2_X1 U2533 ( .A1(n81), .A2(RST), .ZN(n2441) );
  AND2_X1 U2534 ( .A1(n81), .A2(n142), .ZN(n2442) );
  AND2_X1 U2535 ( .A1(n81), .A2(n140), .ZN(n2443) );
  AND2_X1 U2536 ( .A1(n81), .A2(n138), .ZN(n2444) );
  AND2_X1 U2537 ( .A1(n81), .A2(n155), .ZN(n2445) );
  AND2_X1 U2538 ( .A1(n81), .A2(RST), .ZN(n2446) );
  AND2_X1 U2539 ( .A1(n103), .A2(n155), .ZN(n2447) );
  AND2_X1 U2540 ( .A1(n103), .A2(RST), .ZN(n2448) );
  AND2_X1 U2541 ( .A1(n103), .A2(n154), .ZN(n2449) );
  AND2_X1 U2542 ( .A1(n103), .A2(n143), .ZN(n2450) );
  AND2_X1 U2543 ( .A1(n103), .A2(RST), .ZN(n2451) );
  AND2_X1 U2544 ( .A1(n103), .A2(RST), .ZN(n2452) );
  AND2_X1 U2545 ( .A1(n103), .A2(n151), .ZN(n2453) );
  AND2_X1 U2546 ( .A1(n103), .A2(n148), .ZN(n2454) );
  AND2_X1 U2547 ( .A1(n103), .A2(n144), .ZN(n2455) );
  AND2_X1 U2548 ( .A1(n103), .A2(n149), .ZN(n2456) );
  AND2_X1 U2549 ( .A1(n103), .A2(n139), .ZN(n2457) );
  AND2_X1 U2550 ( .A1(n103), .A2(RST), .ZN(n2458) );
  AND2_X1 U2551 ( .A1(n103), .A2(RST), .ZN(n2459) );
  AND2_X1 U2552 ( .A1(n103), .A2(n142), .ZN(n2460) );
  AND2_X1 U2553 ( .A1(n103), .A2(n141), .ZN(n2461) );
  AND2_X1 U2554 ( .A1(n103), .A2(RST), .ZN(n2462) );
  AND2_X1 U2555 ( .A1(n103), .A2(n155), .ZN(n2463) );
  AND2_X1 U2556 ( .A1(n103), .A2(n141), .ZN(n2464) );
  AND2_X1 U2557 ( .A1(n103), .A2(n139), .ZN(n2465) );
  AND2_X1 U2558 ( .A1(n103), .A2(n137), .ZN(n2466) );
  AND2_X1 U2559 ( .A1(n103), .A2(RST), .ZN(n2467) );
  AND2_X1 U2560 ( .A1(n103), .A2(RST), .ZN(n2468) );
  AND2_X1 U2561 ( .A1(n113), .A2(n155), .ZN(n2469) );
  AND2_X1 U2562 ( .A1(n113), .A2(RST), .ZN(n2470) );
  AND2_X1 U2563 ( .A1(n113), .A2(n154), .ZN(n2471) );
  AND2_X1 U2564 ( .A1(n113), .A2(n147), .ZN(n2472) );
  AND2_X1 U2565 ( .A1(n113), .A2(RST), .ZN(n2473) );
  AND2_X1 U2566 ( .A1(n113), .A2(RST), .ZN(n2474) );
  AND2_X1 U2567 ( .A1(n113), .A2(n151), .ZN(n2475) );
  AND2_X1 U2568 ( .A1(n113), .A2(n155), .ZN(n2476) );
  AND2_X1 U2569 ( .A1(n113), .A2(RST), .ZN(n2477) );
  AND2_X1 U2570 ( .A1(n113), .A2(n151), .ZN(n2478) );
  AND2_X1 U2571 ( .A1(n113), .A2(RST), .ZN(n2479) );
  AND2_X1 U2572 ( .A1(n113), .A2(RST), .ZN(n2480) );
  AND2_X1 U2573 ( .A1(n113), .A2(RST), .ZN(n2481) );
  AND2_X1 U2574 ( .A1(n113), .A2(n137), .ZN(n2482) );
  AND2_X1 U2575 ( .A1(n113), .A2(RST), .ZN(n2483) );
  AND2_X1 U2576 ( .A1(n113), .A2(n142), .ZN(n2484) );
  AND2_X1 U2577 ( .A1(n113), .A2(n152), .ZN(n2485) );
  AND2_X1 U2578 ( .A1(n113), .A2(n141), .ZN(n2486) );
  AND2_X1 U2579 ( .A1(n113), .A2(n139), .ZN(n2487) );
  AND2_X1 U2580 ( .A1(n113), .A2(n137), .ZN(n2488) );
  AND2_X1 U2581 ( .A1(n113), .A2(n151), .ZN(n2489) );
  AND2_X1 U2582 ( .A1(n113), .A2(RST), .ZN(n2490) );
  AND2_X1 U2583 ( .A1(n99), .A2(n155), .ZN(n2491) );
  AND2_X1 U2584 ( .A1(n1640), .A2(RST), .ZN(n2492) );
  AND2_X1 U2585 ( .A1(n1640), .A2(n148), .ZN(n2493) );
  AND2_X1 U2586 ( .A1(n1640), .A2(RST), .ZN(n2494) );
  AND2_X1 U2587 ( .A1(n1640), .A2(RST), .ZN(n2495) );
  AND2_X1 U2588 ( .A1(n1640), .A2(RST), .ZN(n2496) );
  AND2_X1 U2589 ( .A1(n1640), .A2(n145), .ZN(n2497) );
  AND2_X1 U2590 ( .A1(n1640), .A2(n144), .ZN(n2498) );
  AND2_X1 U2591 ( .A1(n1640), .A2(n143), .ZN(n2499) );
  AND2_X1 U2592 ( .A1(n1640), .A2(RST), .ZN(n2500) );
  AND2_X1 U2593 ( .A1(n1635), .A2(n151), .ZN(n2501) );
  AND2_X1 U2594 ( .A1(n1635), .A2(n149), .ZN(n2502) );
  AND2_X1 U2595 ( .A1(n1635), .A2(n147), .ZN(n2503) );
  AND2_X1 U2596 ( .A1(n1635), .A2(RST), .ZN(n2504) );
  AND2_X1 U2597 ( .A1(n1635), .A2(n143), .ZN(n2505) );
  AND2_X1 U2598 ( .A1(n1634), .A2(RST), .ZN(n2506) );
  AND2_X1 U2599 ( .A1(n1634), .A2(n149), .ZN(n2507) );
  AND2_X1 U2600 ( .A1(n1634), .A2(n147), .ZN(n2508) );
  AND2_X1 U2601 ( .A1(n1634), .A2(RST), .ZN(n2509) );
  AND2_X1 U2602 ( .A1(n1634), .A2(n155), .ZN(n2510) );
  AND2_X1 U2603 ( .A1(n1633), .A2(n155), .ZN(n2511) );
  AND2_X1 U2604 ( .A1(n1633), .A2(n149), .ZN(n2512) );
  AND2_X1 U2605 ( .A1(n1633), .A2(n147), .ZN(n2513) );
  AND2_X1 U2606 ( .A1(n1633), .A2(RST), .ZN(n2514) );
  AND2_X1 U2607 ( .A1(n1645), .A2(n155), .ZN(n2515) );
  AND2_X1 U2608 ( .A1(n1645), .A2(n149), .ZN(n2516) );
  AND2_X1 U2609 ( .A1(n1645), .A2(n147), .ZN(n2517) );
  AND2_X1 U2610 ( .A1(n1645), .A2(RST), .ZN(n2518) );
  AND2_X1 U2611 ( .A1(n1645), .A2(n149), .ZN(n2519) );
  AND2_X1 U2612 ( .A1(n1645), .A2(n146), .ZN(n2520) );
  AND2_X1 U2613 ( .A1(n1645), .A2(RST), .ZN(n2521) );
  AND2_X1 U2614 ( .A1(n1645), .A2(n146), .ZN(n2522) );
  AND2_X1 U2615 ( .A1(n1645), .A2(RST), .ZN(n2523) );
  AND2_X1 U2616 ( .A1(n1645), .A2(RST), .ZN(n2524) );
  AND2_X1 U2617 ( .A1(n1792), .A2(n148), .ZN(n2525) );
  AND2_X1 U2618 ( .A1(n1792), .A2(RST), .ZN(n2526) );
  AND2_X1 U2619 ( .A1(n1792), .A2(n148), .ZN(n2527) );
  AND2_X1 U2620 ( .A1(n1792), .A2(RST), .ZN(n2528) );
  AND2_X1 U2621 ( .A1(n1792), .A2(RST), .ZN(n2529) );
  AND2_X1 U2622 ( .A1(n1792), .A2(RST), .ZN(n2530) );
  AND2_X1 U2623 ( .A1(n1792), .A2(n145), .ZN(n2531) );
  AND2_X1 U2624 ( .A1(n1792), .A2(RST), .ZN(n2532) );
  AND2_X1 U2625 ( .A1(n1792), .A2(n138), .ZN(n2533) );
  AND2_X1 U2626 ( .A1(n1792), .A2(n146), .ZN(n2534) );
  AND2_X1 U2627 ( .A1(n1794), .A2(n152), .ZN(n2535) );
  AND2_X1 U2628 ( .A1(n1794), .A2(n149), .ZN(n2536) );
  AND2_X1 U2629 ( .A1(n1794), .A2(n147), .ZN(n2537) );
  AND2_X1 U2630 ( .A1(n1794), .A2(RST), .ZN(n2538) );
  AND2_X1 U2631 ( .A1(n1794), .A2(RST), .ZN(n2539) );
  AND2_X1 U2632 ( .A1(n1794), .A2(n146), .ZN(n2540) );
  AND2_X1 U2633 ( .A1(n1794), .A2(RST), .ZN(n2541) );
  AND2_X1 U2634 ( .A1(n1794), .A2(RST), .ZN(n2542) );
  AND2_X1 U2635 ( .A1(n1794), .A2(RST), .ZN(n2543) );
  AND2_X1 U2636 ( .A1(n1794), .A2(n151), .ZN(n2544) );
  AND2_X1 U2637 ( .A1(n1631), .A2(RST), .ZN(n2545) );
  AND2_X1 U2638 ( .A1(n1631), .A2(n148), .ZN(n2546) );
  AND2_X1 U2639 ( .A1(n1631), .A2(RST), .ZN(n2547) );
  AND2_X1 U2640 ( .A1(n1631), .A2(n149), .ZN(n2548) );
  AND2_X1 U2641 ( .A1(n1631), .A2(RST), .ZN(n2549) );
  AND2_X1 U2642 ( .A1(n1631), .A2(n145), .ZN(n2550) );
  AND2_X1 U2643 ( .A1(n1631), .A2(n144), .ZN(n2551) );
  AND2_X1 U2644 ( .A1(n1631), .A2(n143), .ZN(n2552) );
  AND2_X1 U2645 ( .A1(n1631), .A2(n151), .ZN(n2553) );
  AND2_X1 U2646 ( .A1(n1631), .A2(RST), .ZN(n2554) );
  AND2_X1 U2647 ( .A1(n1790), .A2(RST), .ZN(n2555) );
  AND2_X1 U2648 ( .A1(n1790), .A2(n149), .ZN(n2556) );
  AND2_X1 U2649 ( .A1(n1790), .A2(n147), .ZN(n2557) );
  AND2_X1 U2650 ( .A1(n1790), .A2(RST), .ZN(n2558) );
  AND2_X1 U2651 ( .A1(n1790), .A2(RST), .ZN(n2559) );
  AND2_X1 U2652 ( .A1(n1790), .A2(n146), .ZN(n2560) );
  AND2_X1 U2653 ( .A1(n1790), .A2(RST), .ZN(n2561) );
  AND2_X1 U2654 ( .A1(n1790), .A2(n152), .ZN(n2562) );
  AND2_X1 U2655 ( .A1(n1790), .A2(RST), .ZN(n2563) );
  AND2_X1 U2656 ( .A1(n1790), .A2(n140), .ZN(n2564) );
  AND2_X1 U2657 ( .A1(DATAIN[10]), .A2(n145), .ZN(n2565) );
  AND2_X1 U2658 ( .A1(DATAIN[10]), .A2(n149), .ZN(n2566) );
  AND2_X1 U2659 ( .A1(DATAIN[10]), .A2(n147), .ZN(n2567) );
  AND2_X1 U2660 ( .A1(DATAIN[10]), .A2(RST), .ZN(n2568) );
  AND2_X1 U2661 ( .A1(DATAIN[10]), .A2(n153), .ZN(n2569) );
  AND2_X1 U2662 ( .A1(DATAIN[10]), .A2(n146), .ZN(n2570) );
  AND2_X1 U2663 ( .A1(DATAIN[10]), .A2(n144), .ZN(n2571) );
  AND2_X1 U2664 ( .A1(DATAIN[10]), .A2(n143), .ZN(n2572) );
  AND2_X1 U2665 ( .A1(DATAIN[10]), .A2(n139), .ZN(n2573) );
  AND2_X1 U2666 ( .A1(DATAIN[10]), .A2(n144), .ZN(n2574) );
  AND2_X1 U2667 ( .A1(n1630), .A2(n143), .ZN(n2575) );
  AND2_X1 U2668 ( .A1(n1630), .A2(n149), .ZN(n2576) );
  AND2_X1 U2669 ( .A1(n1630), .A2(n147), .ZN(n2577) );
  AND2_X1 U2670 ( .A1(n1630), .A2(RST), .ZN(n2578) );
  AND2_X1 U2671 ( .A1(n1630), .A2(RST), .ZN(n2579) );
  AND2_X1 U2672 ( .A1(n1630), .A2(n146), .ZN(n2580) );
  AND2_X1 U2673 ( .A1(n1630), .A2(RST), .ZN(n2581) );
  AND2_X1 U2674 ( .A1(n1630), .A2(RST), .ZN(n2582) );
  AND2_X1 U2675 ( .A1(n1630), .A2(n144), .ZN(n2583) );
  AND2_X1 U2676 ( .A1(n1630), .A2(n142), .ZN(n2584) );
  AND2_X1 U2677 ( .A1(n1791), .A2(n154), .ZN(n2585) );
  AND2_X1 U2678 ( .A1(n1791), .A2(n149), .ZN(n2586) );
  AND2_X1 U2679 ( .A1(n1791), .A2(n147), .ZN(n2587) );
  AND2_X1 U2680 ( .A1(n1791), .A2(RST), .ZN(n2588) );
  AND2_X1 U2681 ( .A1(n1791), .A2(RST), .ZN(n2589) );
  AND2_X1 U2682 ( .A1(n1791), .A2(n146), .ZN(n2590) );
  AND2_X1 U2683 ( .A1(n1791), .A2(RST), .ZN(n2591) );
  AND2_X1 U2684 ( .A1(n1791), .A2(n153), .ZN(n2592) );
  AND2_X1 U2685 ( .A1(n1791), .A2(RST), .ZN(n2593) );
  AND2_X1 U2686 ( .A1(n1791), .A2(n144), .ZN(n2594) );
  AND2_X1 U2687 ( .A1(n1793), .A2(RST), .ZN(n2595) );
  AND2_X1 U2688 ( .A1(n1793), .A2(RST), .ZN(n2596) );
  AND2_X1 U2689 ( .A1(n1793), .A2(n148), .ZN(n2597) );
  AND2_X1 U2690 ( .A1(n1793), .A2(RST), .ZN(n2598) );
  AND2_X1 U2691 ( .A1(n1793), .A2(RST), .ZN(n2599) );
  AND2_X1 U2692 ( .A1(n1793), .A2(RST), .ZN(n2600) );
  AND2_X1 U2693 ( .A1(n1793), .A2(n145), .ZN(n2601) );
  AND2_X1 U2694 ( .A1(n1793), .A2(RST), .ZN(n2602) );
  AND2_X1 U2695 ( .A1(n1793), .A2(n142), .ZN(n2603) );
  AND2_X1 U2696 ( .A1(n1793), .A2(RST), .ZN(n2604) );
  AND2_X1 U2697 ( .A1(n1789), .A2(RST), .ZN(n2605) );
  AND2_X1 U2698 ( .A1(n1789), .A2(n149), .ZN(n2606) );
  AND2_X1 U2699 ( .A1(n1789), .A2(n147), .ZN(n2607) );
  AND2_X1 U2700 ( .A1(n1789), .A2(RST), .ZN(n2608) );
  AND2_X1 U2701 ( .A1(n1789), .A2(n152), .ZN(n2609) );
  AND2_X1 U2702 ( .A1(n1789), .A2(n146), .ZN(n2610) );
  AND2_X1 U2703 ( .A1(n1789), .A2(n147), .ZN(n2611) );
  AND2_X1 U2704 ( .A1(n1789), .A2(n151), .ZN(n2612) );
  AND2_X1 U2705 ( .A1(n1789), .A2(RST), .ZN(n2613) );
  AND2_X1 U2706 ( .A1(n1789), .A2(n141), .ZN(n2614) );
  AND2_X1 U2707 ( .A1(n1644), .A2(RST), .ZN(n2615) );
  AND2_X1 U2708 ( .A1(n1644), .A2(n149), .ZN(n2616) );
  AND2_X1 U2709 ( .A1(n1644), .A2(n147), .ZN(n2617) );
  AND2_X1 U2710 ( .A1(n1644), .A2(RST), .ZN(n2618) );
  AND2_X1 U2711 ( .A1(n1644), .A2(n150), .ZN(n2619) );
  AND2_X1 U2712 ( .A1(n1644), .A2(n146), .ZN(n2620) );
  AND2_X1 U2713 ( .A1(n1644), .A2(n147), .ZN(n2621) );
  AND2_X1 U2714 ( .A1(n1644), .A2(RST), .ZN(n2622) );
  AND2_X1 U2715 ( .A1(n1644), .A2(RST), .ZN(n2623) );
  AND2_X1 U2716 ( .A1(n1644), .A2(RST), .ZN(n2624) );
  AND2_X1 U2717 ( .A1(n1642), .A2(n150), .ZN(n2625) );
  AND2_X1 U2718 ( .A1(n1642), .A2(RST), .ZN(n2626) );
  AND2_X1 U2719 ( .A1(n1642), .A2(n148), .ZN(n2627) );
  AND2_X1 U2720 ( .A1(n1642), .A2(RST), .ZN(n2628) );
  AND2_X1 U2721 ( .A1(n1642), .A2(RST), .ZN(n2629) );
  AND2_X1 U2722 ( .A1(n1642), .A2(RST), .ZN(n2630) );
  AND2_X1 U2723 ( .A1(n1642), .A2(n145), .ZN(n2631) );
  AND2_X1 U2724 ( .A1(n1642), .A2(RST), .ZN(n2632) );
  AND2_X1 U2725 ( .A1(n1642), .A2(n150), .ZN(n2633) );
  AND2_X1 U2726 ( .A1(n1643), .A2(n144), .ZN(n2634) );
  AND2_X1 U2727 ( .A1(n1643), .A2(RST), .ZN(n2635) );
  AND2_X1 U2728 ( .A1(n1643), .A2(n148), .ZN(n2636) );
  AND2_X1 U2729 ( .A1(n1643), .A2(RST), .ZN(n2637) );
  AND2_X1 U2730 ( .A1(n1643), .A2(n153), .ZN(n2638) );
  AND2_X1 U2731 ( .A1(n1643), .A2(RST), .ZN(n2639) );
  AND2_X1 U2732 ( .A1(n1643), .A2(n145), .ZN(n2640) );
  AND2_X1 U2733 ( .A1(n1643), .A2(RST), .ZN(n2641) );
  AND2_X1 U2734 ( .A1(n1643), .A2(n141), .ZN(n2642) );
  AND2_X1 U2735 ( .A1(n1632), .A2(n149), .ZN(n2643) );
  AND2_X1 U2736 ( .A1(n1632), .A2(n149), .ZN(n2644) );
  AND2_X1 U2737 ( .A1(n1632), .A2(n147), .ZN(n2645) );
  AND2_X1 U2738 ( .A1(n1632), .A2(RST), .ZN(n2646) );
  AND2_X1 U2739 ( .A1(n1632), .A2(n145), .ZN(n2647) );
  AND2_X1 U2740 ( .A1(n1632), .A2(n146), .ZN(n2648) );
  AND2_X1 U2741 ( .A1(n1632), .A2(RST), .ZN(n2649) );
  AND2_X1 U2742 ( .A1(n1632), .A2(n148), .ZN(n2650) );
  AND2_X1 U2743 ( .A1(n1632), .A2(n146), .ZN(n2651) );
  AND2_X1 U2744 ( .A1(n1632), .A2(RST), .ZN(n2652) );
  AND2_X1 U2745 ( .A1(n1641), .A2(n143), .ZN(n2653) );
  AND2_X1 U2746 ( .A1(n1641), .A2(RST), .ZN(n2654) );
  AND2_X1 U2747 ( .A1(n1641), .A2(n148), .ZN(n2655) );
  AND2_X1 U2748 ( .A1(n1641), .A2(RST), .ZN(n2656) );
  AND2_X1 U2749 ( .A1(n1641), .A2(RST), .ZN(n2657) );
  AND2_X1 U2750 ( .A1(n1641), .A2(RST), .ZN(n2658) );
  AND2_X1 U2751 ( .A1(n1641), .A2(n145), .ZN(n2659) );
  AND2_X1 U2752 ( .A1(n1641), .A2(RST), .ZN(n2660) );
  AND2_X1 U2753 ( .A1(n1641), .A2(RST), .ZN(n2661) );
  AND2_X1 U2754 ( .A1(n1638), .A2(n144), .ZN(n2662) );
  AND2_X1 U2755 ( .A1(n1638), .A2(RST), .ZN(n2663) );
  AND2_X1 U2756 ( .A1(n1638), .A2(n148), .ZN(n2664) );
  AND2_X1 U2757 ( .A1(n1638), .A2(RST), .ZN(n2665) );
  AND2_X1 U2758 ( .A1(n1638), .A2(RST), .ZN(n2666) );
  AND2_X1 U2759 ( .A1(n1638), .A2(RST), .ZN(n2667) );
  AND2_X1 U2760 ( .A1(n1638), .A2(n145), .ZN(n2668) );
  AND2_X1 U2761 ( .A1(n1638), .A2(RST), .ZN(n2669) );
  AND2_X1 U2762 ( .A1(n1638), .A2(RST), .ZN(n2670) );
  AND2_X1 U2763 ( .A1(DATAIN[23]), .A2(n146), .ZN(n2671) );
  AND2_X1 U2764 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2672) );
  AND2_X1 U2765 ( .A1(DATAIN[23]), .A2(n148), .ZN(n2673) );
  AND2_X1 U2766 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2674) );
  AND2_X1 U2767 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2675) );
  AND2_X1 U2768 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2676) );
  AND2_X1 U2769 ( .A1(DATAIN[23]), .A2(n145), .ZN(n2677) );
  AND2_X1 U2770 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2678) );
  AND2_X1 U2771 ( .A1(DATAIN[23]), .A2(n151), .ZN(n2679) );
  AND2_X1 U2772 ( .A1(DATAIN[30]), .A2(n153), .ZN(n2680) );
  AND2_X1 U2773 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2681) );
  AND2_X1 U2774 ( .A1(DATAIN[30]), .A2(n148), .ZN(n2682) );
  AND2_X1 U2775 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2683) );
  AND2_X1 U2776 ( .A1(DATAIN[30]), .A2(n144), .ZN(n2684) );
  AND2_X1 U2777 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2685) );
  AND2_X1 U2778 ( .A1(DATAIN[30]), .A2(n145), .ZN(n2686) );
  AND2_X1 U2779 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2687) );
  AND2_X1 U2780 ( .A1(DATAIN[30]), .A2(n150), .ZN(n2688) );
  AND2_X1 U2781 ( .A1(DATAIN[4]), .A2(RST), .ZN(n2689) );
  AND2_X1 U2782 ( .A1(DATAIN[4]), .A2(n148), .ZN(n2690) );
  AND2_X1 U2783 ( .A1(DATAIN[4]), .A2(RST), .ZN(n2691) );
  AND2_X1 U2784 ( .A1(DATAIN[4]), .A2(n145), .ZN(n2692) );
  AND2_X1 U2785 ( .A1(DATAIN[4]), .A2(RST), .ZN(n2693) );
  AND2_X1 U2786 ( .A1(DATAIN[4]), .A2(n145), .ZN(n2694) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_0 \clk_gate_REGISTERS_reg[0]  ( 
        .CLK(CLK), .EN(N144), .ENCLK(net7104), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_31 \clk_gate_REGISTERS_reg[1]  ( 
        .CLK(CLK), .EN(N143), .ENCLK(net7110), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_30 \clk_gate_REGISTERS_reg[2]  ( 
        .CLK(CLK), .EN(N142), .ENCLK(net7115), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_29 \clk_gate_REGISTERS_reg[3]  ( 
        .CLK(CLK), .EN(N141), .ENCLK(net7120), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_28 \clk_gate_REGISTERS_reg[4]  ( 
        .CLK(CLK), .EN(N140), .ENCLK(net7125), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_27 \clk_gate_REGISTERS_reg[5]  ( 
        .CLK(CLK), .EN(N139), .ENCLK(net7130), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_26 \clk_gate_REGISTERS_reg[6]  ( 
        .CLK(CLK), .EN(N138), .ENCLK(net7135), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_25 \clk_gate_REGISTERS_reg[7]  ( 
        .CLK(CLK), .EN(N137), .ENCLK(net7140), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_24 \clk_gate_REGISTERS_reg[8]  ( 
        .CLK(CLK), .EN(N136), .ENCLK(net7145), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_23 \clk_gate_REGISTERS_reg[9]  ( 
        .CLK(CLK), .EN(N135), .ENCLK(net7150), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_22 \clk_gate_REGISTERS_reg[10]  ( 
        .CLK(CLK), .EN(N134), .ENCLK(net7155), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_21 \clk_gate_REGISTERS_reg[11]  ( 
        .CLK(CLK), .EN(N133), .ENCLK(net7160), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_20 \clk_gate_REGISTERS_reg[12]  ( 
        .CLK(CLK), .EN(N132), .ENCLK(net7165), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_19 \clk_gate_REGISTERS_reg[13]  ( 
        .CLK(CLK), .EN(N131), .ENCLK(net7170), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_18 \clk_gate_REGISTERS_reg[14]  ( 
        .CLK(CLK), .EN(N130), .ENCLK(net7175), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_17 \clk_gate_REGISTERS_reg[15]  ( 
        .CLK(CLK), .EN(N129), .ENCLK(net7180), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_16 \clk_gate_REGISTERS_reg[16]  ( 
        .CLK(CLK), .EN(N128), .ENCLK(net7185), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_15 \clk_gate_REGISTERS_reg[17]  ( 
        .CLK(CLK), .EN(N127), .ENCLK(net7190), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_14 \clk_gate_REGISTERS_reg[18]  ( 
        .CLK(CLK), .EN(N126), .ENCLK(net7195), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_13 \clk_gate_REGISTERS_reg[19]  ( 
        .CLK(CLK), .EN(N125), .ENCLK(net7200), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_12 \clk_gate_REGISTERS_reg[20]  ( 
        .CLK(CLK), .EN(N124), .ENCLK(net7205), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_11 \clk_gate_REGISTERS_reg[21]  ( 
        .CLK(CLK), .EN(N123), .ENCLK(net7210), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_10 \clk_gate_REGISTERS_reg[22]  ( 
        .CLK(CLK), .EN(N122), .ENCLK(net7215), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_9 \clk_gate_REGISTERS_reg[23]  ( 
        .CLK(CLK), .EN(N121), .ENCLK(net7220), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_8 \clk_gate_REGISTERS_reg[24]  ( 
        .CLK(CLK), .EN(N120), .ENCLK(net7225), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_7 \clk_gate_REGISTERS_reg[25]  ( 
        .CLK(CLK), .EN(N119), .ENCLK(net7230), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_6 \clk_gate_REGISTERS_reg[26]  ( 
        .CLK(CLK), .EN(N118), .ENCLK(net7235), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_5 \clk_gate_REGISTERS_reg[27]  ( 
        .CLK(CLK), .EN(N117), .ENCLK(net7240), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_4 \clk_gate_REGISTERS_reg[28]  ( 
        .CLK(CLK), .EN(N116), .ENCLK(net7245), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_3 \clk_gate_REGISTERS_reg[29]  ( 
        .CLK(CLK), .EN(N115), .ENCLK(net7250), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_2 \clk_gate_REGISTERS_reg[30]  ( 
        .CLK(CLK), .EN(N114), .ENCLK(net7255), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_1 \clk_gate_REGISTERS_reg[31]  ( 
        .CLK(CLK), .EN(N81), .ENCLK(net7260), .TE(1'b0) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n2695), .CK(net7170), .Q(
        \REGISTERS[13][13] ) );
  AND2_X1 U1902 ( .A1(DATAIN[13]), .A2(n146), .ZN(n2695) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH5_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7070, net7072, net7074, net7075, net7078, net7081;
  assign net7070 = EN;
  assign net7072 = CLK;
  assign ENCLK = net7074;
  assign net7081 = TE;

  DLL_X1 latch ( .D(net7075), .GN(net7072), .Q(net7078) );
  OR2_X1 test_or ( .A1(net7070), .A2(net7081), .ZN(net7075) );
  AND2_X1 main_gate ( .A1(net7078), .A2(net7072), .ZN(net7074) );
endmodule


module SNPS_CLOCK_GATE_HIGH_FFD_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7016, net7018, net7020, net7021, net7024, net7027;
  assign net7016 = EN;
  assign net7018 = CLK;
  assign ENCLK = net7020;
  assign net7027 = TE;

  DLL_X1 latch ( .D(net7021), .GN(net7018), .Q(net7024) );
  OR2_X1 test_or ( .A1(net7016), .A2(net7027), .ZN(net7021) );
  AND2_X1 main_gate ( .A1(net7024), .A2(net7018), .ZN(net7020) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_12 ( CLK, EN, ENCLK, TE
 );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  OR2_X1 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
  AND2_X2 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_11 ( CLK, EN, ENCLK, TE
 );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  AND2_X2 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
  OR2_X2 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_10 ( CLK, EN, ENCLK, TE
 );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  OR2_X1 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
  AND2_X1 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  OR2_X1 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
  AND2_X1 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  OR2_X1 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
  AND2_X1 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  OR2_X1 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
  AND2_X1 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  OR2_X1 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
  AND2_X1 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  OR2_X1 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
  AND2_X1 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  OR2_X1 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
  AND2_X1 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH5_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7070, net7072, net7074, net7075, net7078, net7081;
  assign net7070 = EN;
  assign net7072 = CLK;
  assign ENCLK = net7074;
  assign net7081 = TE;

  DLL_X1 latch ( .D(net7075), .GN(net7072), .Q(net7078) );
  OR2_X1 test_or ( .A1(net7070), .A2(net7081), .ZN(net7075) );
  AND2_X1 main_gate ( .A1(net7078), .A2(net7072), .ZN(net7074) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  OR2_X1 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
  AND2_X1 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  OR2_X1 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
  AND2_X1 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH5_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7070, net7072, net7074, net7075, net7078, net7081;
  assign net7070 = EN;
  assign net7072 = CLK;
  assign ENCLK = net7074;
  assign net7081 = TE;

  DLL_X1 latch ( .D(net7075), .GN(net7072), .Q(net7078) );
  OR2_X1 test_or ( .A1(net7070), .A2(net7081), .ZN(net7075) );
  AND2_X1 main_gate ( .A1(net7078), .A2(net7072), .ZN(net7074) );
endmodule


module SNPS_CLOCK_GATE_HIGH_FFD_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7016, net7018, net7020, net7021, net7024, net7027;
  assign net7016 = EN;
  assign net7018 = CLK;
  assign ENCLK = net7020;
  assign net7027 = TE;

  DLL_X1 latch ( .D(net7021), .GN(net7018), .Q(net7024) );
  OR2_X1 test_or ( .A1(net7016), .A2(net7027), .ZN(net7021) );
  AND2_X1 main_gate ( .A1(net7024), .A2(net7018), .ZN(net7020) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net7052, net7054, net7056, net7057, net7060, net7063;
  assign net7052 = EN;
  assign net7054 = CLK;
  assign ENCLK = net7056;
  assign net7063 = TE;

  DLL_X1 latch ( .D(net7057), .GN(net7054), .Q(net7060) );
  OR2_X1 test_or ( .A1(net7052), .A2(net7063), .ZN(net7057) );
  AND2_X1 main_gate ( .A1(net7060), .A2(net7054), .ZN(net7056) );
endmodule


module DLX_WIDTH32 ( CLK, RST, IROM_ADDR, IROM_DATA, DRAM_EN, DRAM_RW, 
        DRAM_ADDR, DRAM_DATA_IN, DRAM_DATA_OUT );
  output [11:0] IROM_ADDR;
  input [31:0] IROM_DATA;
  output [11:0] DRAM_ADDR;
  input [31:0] DRAM_DATA_IN;
  output [31:0] DRAM_DATA_OUT;
  input CLK, RST;
  output DRAM_EN, DRAM_RW;
  wire   w_IF_EN, w_RF_RD1, w_RF_RD2, w_EX_EN, w_MuxA_SEL, w_MuxB_SEL,
         w_JUMP_EQ, w_RegME_LATCH_EN, w_RegRD2_LATCH_EN, w_RF_WE_EX, w_SIGN_LD,
         w_RegALU2_LATCH_EN, w_RegLMD_LATCH_EN, w_RegRD3_LATCH_EN, w_MuxWB_SEL,
         w_RF_WE, \PC/N34 , \PC/N33 , \PC/N32 , \PC/N31 , \PC/N30 , \PC/N29 ,
         \PC/N28 , \PC/N27 , \PC/N26 , \PC/N25 , \PC/N24 , \PC/N23 , \PC/N22 ,
         \PC/N21 , \PC/N20 , \PC/N19 , \PC/N18 , \PC/N17 , \PC/N16 , \PC/N15 ,
         \PC/N14 , \PC/N13 , \PC/N12 , \PC/N11 , \PC/N10 , \PC/N9 , \PC/N8 ,
         \PC/N7 , \PC/N6 , \PC/N5 , \PC/N4 , \PC/N3 , \PC/N2 , \CU/N89 ,
         \CU/N88 , \CU/N87 , \CU/N86 , \CU/N85 , \CU/N82 , \CU/N81 , \CU/N80 ,
         \CU/N79 , \CU/N78 , \CU/N77 , \CU/N76 , \CU/N75 , \CU/N74 , \CU/N73 ,
         \CU/N72 , \CU/N71 , \CU/N70 , \CU/N69 , \CU/N68 , \CU/N67 , \CU/N66 ,
         \CU/N65 , \CU/N64 , \CU/N63 , \CU/N62 , \CU/N61 , \CU/N60 , \CU/N59 ,
         \CU/N58 , \CU/N56 , \CU/N55 , \CU/N54 , \CU/N52 , \CU/N51 , \CU/N50 ,
         \CU/N49 , \CU/N48 , \CU/N47 , \CU/N46 , \CU/N45 , \CU/N42 ,
         \CU/cw2[2] , \CU/cw2[1] , \CU/cw1[14] , \CU/cw1[13] , \CU/cw1[12] ,
         \CU/cw1[11] , \CU/cw1[10] , \CU/cw1[9] , \CU/cw1[8] , \CU/cw1[7] ,
         \CU/cw1[6] , \CU/cw1[5] , \CU/cw1[4] , \CU/cw1[3] , \CU/cw1[2] ,
         \CU/cw1[1] , \CU/JUMP3 , \CU/JUMP2 , \DP/RegLMD_out[31] ,
         \DP/RegLMD_out[30] , \DP/RegLMD_out[29] , \DP/RegLMD_out[28] ,
         \DP/RegLMD_out[27] , \DP/RegLMD_out[26] , \DP/RegLMD_out[25] ,
         \DP/RegLMD_out[24] , \DP/RegLMD_out[23] , \DP/RegLMD_out[22] ,
         \DP/RegLMD_out[21] , \DP/RegLMD_out[20] , \DP/RegLMD_out[19] ,
         \DP/RegLMD_out[18] , \DP/RegLMD_out[17] , \DP/RegLMD_out[16] ,
         \DP/RegLMD_out[15] , \DP/RegLMD_out[14] , \DP/RegLMD_out[13] ,
         \DP/RegLMD_out[12] , \DP/RegLMD_out[11] , \DP/RegLMD_out[10] ,
         \DP/RegLMD_out[9] , \DP/RegLMD_out[8] , \DP/RegLMD_out[7] ,
         \DP/RegLMD_out[6] , \DP/RegLMD_out[5] , \DP/RegLMD_out[4] ,
         \DP/RegLMD_out[3] , \DP/RegLMD_out[2] , \DP/RegLMD_out[1] ,
         \DP/RegLMD_out[0] , \DP/RegALU2_out[31] , \DP/RegALU2_out[30] ,
         \DP/RegALU2_out[29] , \DP/RegALU2_out[28] , \DP/RegALU2_out[27] ,
         \DP/RegALU2_out[26] , \DP/RegALU2_out[25] , \DP/RegALU2_out[24] ,
         \DP/RegALU2_out[23] , \DP/RegALU2_out[22] , \DP/RegALU2_out[21] ,
         \DP/RegALU2_out[20] , \DP/RegALU2_out[19] , \DP/RegALU2_out[18] ,
         \DP/RegALU2_out[17] , \DP/RegALU2_out[16] , \DP/RegALU2_out[15] ,
         \DP/RegALU2_out[14] , \DP/RegALU2_out[13] , \DP/RegALU2_out[12] ,
         \DP/RegALU2_out[11] , \DP/RegALU2_out[10] , \DP/RegALU2_out[9] ,
         \DP/RegALU2_out[8] , \DP/RegALU2_out[7] , \DP/RegALU2_out[6] ,
         \DP/RegALU2_out[5] , \DP/RegALU2_out[4] , \DP/RegALU2_out[3] ,
         \DP/RegALU2_out[2] , \DP/RegALU2_out[1] , \DP/RegALU2_out[0] ,
         \DP/LOAD8[7] , \DP/LOAD8[6] , \DP/LOAD8[5] , \DP/LOAD8[4] ,
         \DP/LOAD8[3] , \DP/LOAD8[2] , \DP/LOAD8[1] , \DP/LOAD8[0] ,
         \DP/LOAD16[15] , \DP/LOAD16[14] , \DP/LOAD16[13] , \DP/LOAD16[12] ,
         \DP/LOAD16[11] , \DP/LOAD16[10] , \DP/LOAD16[9] , \DP/LOAD16[8] ,
         \DP/FwdD , \DP/RD2[0] , \DP/RD2[1] , \DP/RD2[2] , \DP/RegME_out[31] ,
         \DP/RegME_out[30] , \DP/RegME_out[29] , \DP/RegME_out[28] ,
         \DP/RegME_out[27] , \DP/RegME_out[26] , \DP/RegME_out[25] ,
         \DP/RegME_out[24] , \DP/RegME_out[23] , \DP/RegME_out[22] ,
         \DP/RegME_out[21] , \DP/RegME_out[20] , \DP/RegME_out[19] ,
         \DP/RegME_out[18] , \DP/RegME_out[17] , \DP/RegME_out[16] ,
         \DP/RegME_out[15] , \DP/RegME_out[14] , \DP/RegME_out[13] ,
         \DP/RegME_out[12] , \DP/RegME_out[11] , \DP/RegME_out[10] ,
         \DP/RegME_out[9] , \DP/RegME_out[8] , \DP/RegME_out[7] ,
         \DP/NPC3[31] , \DP/NPC3[30] , \DP/NPC3[29] , \DP/NPC3[28] ,
         \DP/NPC3[27] , \DP/NPC3[26] , \DP/NPC3[25] , \DP/NPC3[24] ,
         \DP/NPC3[23] , \DP/NPC3[22] , \DP/NPC3[21] , \DP/NPC3[20] ,
         \DP/NPC3[19] , \DP/NPC3[18] , \DP/NPC3[17] , \DP/NPC3[16] ,
         \DP/NPC3[15] , \DP/NPC3[14] , \DP/NPC3[13] , \DP/NPC3[12] ,
         \DP/NPC3[11] , \DP/NPC3[10] , \DP/NPC3[9] , \DP/NPC3[8] ,
         \DP/NPC3[7] , \DP/NPC3[6] , \DP/NPC3[5] , \DP/NPC3[4] , \DP/NPC3[3] ,
         \DP/NPC3[2] , \DP/NPC3[1] , \DP/NPC3[0] , \DP/JREG , \DP/JL1 ,
         \DP/RegA1_out[31] , \DP/RegA1_out[30] , \DP/RegA1_out[29] ,
         \DP/RegA1_out[28] , \DP/RegA1_out[27] , \DP/RegA1_out[26] ,
         \DP/RegA1_out[25] , \DP/RegA1_out[24] , \DP/RegA1_out[23] ,
         \DP/RegA1_out[22] , \DP/RegA1_out[21] , \DP/RegA1_out[20] ,
         \DP/RegA1_out[19] , \DP/RegA1_out[18] , \DP/RegA1_out[17] ,
         \DP/RegA1_out[16] , \DP/RegA1_out[15] , \DP/RegA1_out[14] ,
         \DP/RegA1_out[13] , \DP/RegA1_out[12] , \DP/RegA1_out[11] ,
         \DP/RegA1_out[10] , \DP/RegA1_out[9] , \DP/RegA1_out[8] ,
         \DP/RegA1_out[7] , \DP/RegA1_out[6] , \DP/RegA1_out[5] ,
         \DP/RegA1_out[4] , \DP/RegA1_out[3] , \DP/RegA1_out[2] ,
         \DP/RegA1_out[1] , \DP/RegA1_out[0] , \DP/RES[31] , \DP/RES[30] ,
         \DP/RES[29] , \DP/RES[28] , \DP/RES[27] , \DP/RES[26] , \DP/RES[25] ,
         \DP/RES[24] , \DP/RES[23] , \DP/RES[22] , \DP/RES[21] , \DP/RES[20] ,
         \DP/RES[19] , \DP/RES[18] , \DP/RES[17] , \DP/RES[16] , \DP/RES[15] ,
         \DP/RES[14] , \DP/RES[13] , \DP/RES[12] , \DP/RES[11] , \DP/RES[10] ,
         \DP/RES[9] , \DP/RES[8] , \DP/RES[7] , \DP/RES[6] , \DP/RES[5] ,
         \DP/RES[4] , \DP/RES[3] , \DP/RES[2] , \DP/RES[1] , \DP/RES[0] ,
         \DP/FwdC[1] , \DP/B[31] , \DP/B[30] , \DP/B[29] , \DP/B[28] ,
         \DP/B[27] , \DP/B[26] , \DP/B[25] , \DP/B[24] , \DP/B[23] ,
         \DP/B[22] , \DP/B[21] , \DP/B[20] , \DP/B[19] , \DP/B[18] ,
         \DP/B[17] , \DP/B[16] , \DP/B[15] , \DP/B[14] , \DP/B[13] ,
         \DP/B[12] , \DP/B[11] , \DP/B[10] , \DP/B[9] , \DP/B[8] , \DP/B[7] ,
         \DP/B[6] , \DP/B[5] , \DP/B[4] , \DP/B[3] , \DP/B[2] , \DP/B[1] ,
         \DP/B[0] , \DP/FwdB[1] , \DP/FwdB[0] , \DP/A[31] , \DP/A[30] ,
         \DP/A[29] , \DP/A[28] , \DP/A[27] , \DP/A[26] , \DP/A[25] ,
         \DP/A[24] , \DP/A[23] , \DP/A[22] , \DP/A[21] , \DP/A[20] ,
         \DP/A[19] , \DP/A[18] , \DP/A[17] , \DP/A[16] , \DP/A[15] ,
         \DP/A[14] , \DP/A[13] , \DP/A[12] , \DP/A[11] , \DP/A[10] , \DP/A[9] ,
         \DP/A[8] , \DP/A[7] , \DP/A[6] , \DP/A[5] , \DP/A[4] , \DP/A[3] ,
         \DP/A[2] , \DP/A[1] , \DP/A[0] , \DP/FwdA[2] , \DP/RegALU1_out[12] ,
         \DP/RegALU1_out[13] , \DP/RegALU1_out[14] , \DP/RegALU1_out[15] ,
         \DP/RegALU1_out[16] , \DP/RegALU1_out[17] , \DP/RegALU1_out[18] ,
         \DP/RegALU1_out[19] , \DP/RegALU1_out[20] , \DP/RegALU1_out[21] ,
         \DP/RegALU1_out[22] , \DP/RegALU1_out[23] , \DP/RegALU1_out[24] ,
         \DP/RegALU1_out[25] , \DP/RegALU1_out[26] , \DP/RegALU1_out[27] ,
         \DP/RegALU1_out[28] , \DP/RegALU1_out[29] , \DP/RegALU1_out[30] ,
         \DP/RegALU1_out[31] , \DP/RD1[0] , \DP/RD1[1] , \DP/RD1[2] ,
         \DP/RD1[3] , \DP/RD1[4] , \DP/RegIMM_out[31] , \DP/RegIMM_out[24] ,
         \DP/RegIMM_out[23] , \DP/RegIMM_out[22] , \DP/RegIMM_out[21] ,
         \DP/RegIMM_out[20] , \DP/RegIMM_out[19] , \DP/RegIMM_out[18] ,
         \DP/RegIMM_out[17] , \DP/RegIMM_out[16] , \DP/RegIMM_out[15] ,
         \DP/RegIMM_out[14] , \DP/RegIMM_out[13] , \DP/RegIMM_out[12] ,
         \DP/RegIMM_out[11] , \DP/RegIMM_out[10] , \DP/RegIMM_out[9] ,
         \DP/RegIMM_out[8] , \DP/RegIMM_out[7] , \DP/RegIMM_out[6] ,
         \DP/RegIMM_out[5] , \DP/RegIMM_out[4] , \DP/RegIMM_out[3] ,
         \DP/RegIMM_out[2] , \DP/RegIMM_out[1] , \DP/RegIMM_out[0] ,
         \DP/RegB_out[0] , \DP/RegB_out[1] , \DP/RegB_out[2] ,
         \DP/RegB_out[3] , \DP/RegB_out[4] , \DP/RegB_out[5] ,
         \DP/RegB_out[6] , \DP/RegB_out[7] , \DP/RegB_out[8] ,
         \DP/RegB_out[9] , \DP/RegB_out[10] , \DP/RegB_out[11] ,
         \DP/RegB_out[12] , \DP/RegB_out[13] , \DP/RegB_out[14] ,
         \DP/RegB_out[15] , \DP/RegB_out[16] , \DP/RegB_out[17] ,
         \DP/RegB_out[18] , \DP/RegB_out[19] , \DP/RegB_out[20] ,
         \DP/RegB_out[21] , \DP/RegB_out[22] , \DP/RegB_out[23] ,
         \DP/RegB_out[24] , \DP/RegB_out[25] , \DP/RegB_out[26] ,
         \DP/RegB_out[27] , \DP/RegB_out[28] , \DP/RegB_out[29] ,
         \DP/RegB_out[30] , \DP/RegB_out[31] , \DP/RegA_out[0] ,
         \DP/RegA_out[1] , \DP/RegA_out[2] , \DP/RegA_out[3] ,
         \DP/RegA_out[4] , \DP/RegA_out[5] , \DP/RegA_out[6] ,
         \DP/RegA_out[7] , \DP/RegA_out[8] , \DP/RegA_out[9] ,
         \DP/RegA_out[10] , \DP/RegA_out[11] , \DP/RegA_out[12] ,
         \DP/RegA_out[13] , \DP/RegA_out[14] , \DP/RegA_out[15] ,
         \DP/RegA_out[16] , \DP/RegA_out[17] , \DP/RegA_out[18] ,
         \DP/RegA_out[19] , \DP/RegA_out[20] , \DP/RegA_out[21] ,
         \DP/RegA_out[22] , \DP/RegA_out[23] , \DP/RegA_out[24] ,
         \DP/RegA_out[25] , \DP/RegA_out[26] , \DP/RegA_out[27] ,
         \DP/RegA_out[28] , \DP/RegA_out[29] , \DP/RegA_out[30] ,
         \DP/RegA_out[31] , \DP/NPC2[0] , \DP/NPC2[1] , \DP/NPC2[2] ,
         \DP/NPC2[3] , \DP/NPC2[4] , \DP/NPC2[5] , \DP/NPC2[6] , \DP/NPC2[7] ,
         \DP/NPC2[8] , \DP/NPC2[9] , \DP/NPC2[10] , \DP/NPC2[11] ,
         \DP/NPC2[12] , \DP/NPC2[13] , \DP/NPC2[14] , \DP/NPC2[15] ,
         \DP/NPC2[16] , \DP/NPC2[17] , \DP/NPC2[18] , \DP/NPC2[19] ,
         \DP/NPC2[20] , \DP/NPC2[21] , \DP/NPC2[22] , \DP/NPC2[23] ,
         \DP/NPC2[24] , \DP/NPC2[25] , \DP/NPC2[26] , \DP/NPC2[27] ,
         \DP/NPC2[28] , \DP/NPC2[29] , \DP/NPC2[30] , \DP/NPC2[31] ,
         \DP/RegB_in[31] , \DP/RegB_in[30] , \DP/RegB_in[29] ,
         \DP/RegB_in[28] , \DP/RegB_in[27] , \DP/RegB_in[26] ,
         \DP/RegB_in[25] , \DP/RegB_in[24] , \DP/RegB_in[23] ,
         \DP/RegB_in[22] , \DP/RegB_in[21] , \DP/RegB_in[20] ,
         \DP/RegB_in[19] , \DP/RegB_in[18] , \DP/RegB_in[17] ,
         \DP/RegB_in[16] , \DP/RegB_in[15] , \DP/RegB_in[14] ,
         \DP/RegB_in[13] , \DP/RegB_in[12] , \DP/RegB_in[11] ,
         \DP/RegB_in[10] , \DP/RegB_in[9] , \DP/RegB_in[8] , \DP/RegB_in[7] ,
         \DP/RegB_in[6] , \DP/RegB_in[5] , \DP/RegB_in[4] , \DP/RegB_in[3] ,
         \DP/RegB_in[2] , \DP/RegB_in[1] , \DP/RegB_in[0] , \DP/RegA_in[31] ,
         \DP/RegA_in[30] , \DP/RegA_in[29] , \DP/RegA_in[28] ,
         \DP/RegA_in[27] , \DP/RegA_in[26] , \DP/RegA_in[25] ,
         \DP/RegA_in[24] , \DP/RegA_in[23] , \DP/RegA_in[22] ,
         \DP/RegA_in[21] , \DP/RegA_in[20] , \DP/RegA_in[19] ,
         \DP/RegA_in[18] , \DP/RegA_in[17] , \DP/RegA_in[16] ,
         \DP/RegA_in[15] , \DP/RegA_in[14] , \DP/RegA_in[13] ,
         \DP/RegA_in[12] , \DP/RegA_in[11] , \DP/RegA_in[10] , \DP/RegA_in[9] ,
         \DP/RegA_in[8] , \DP/RegA_in[7] , \DP/RegA_in[6] , \DP/RegA_in[5] ,
         \DP/RegA_in[4] , \DP/RegA_in[3] , \DP/RegA_in[2] , \DP/RegA_in[1] ,
         \DP/RegA_in[0] , \DP/RF_ADDR[4] , \DP/RF_ADDR[3] , \DP/RF_ADDR[2] ,
         \DP/RF_ADDR[1] , \DP/RF_ADDR[0] , \DP/RD3[4] , \DP/RD3[3] ,
         \DP/RD3[2] , \DP/RD3[1] , \DP/RD3[0] , \DP/RF_DATA[31] ,
         \DP/RF_DATA[30] , \DP/RF_DATA[29] , \DP/RF_DATA[28] ,
         \DP/RF_DATA[27] , \DP/RF_DATA[26] , \DP/RF_DATA[25] ,
         \DP/RF_DATA[24] , \DP/RF_DATA[23] , \DP/RF_DATA[22] ,
         \DP/RF_DATA[21] , \DP/RF_DATA[20] , \DP/RF_DATA[19] ,
         \DP/RF_DATA[18] , \DP/RF_DATA[17] , \DP/RF_DATA[16] ,
         \DP/RF_DATA[15] , \DP/RF_DATA[14] , \DP/RF_DATA[13] ,
         \DP/RF_DATA[12] , \DP/RF_DATA[11] , \DP/RF_DATA[10] , \DP/RF_DATA[9] ,
         \DP/RF_DATA[8] , \DP/RF_DATA[7] , \DP/RF_DATA[6] , \DP/RF_DATA[5] ,
         \DP/RF_DATA[4] , \DP/RF_DATA[3] , \DP/RF_DATA[2] , \DP/RF_DATA[1] ,
         \DP/RF_DATA[0] , \DP/JL2 , \DP/NPC_out[31] , \DP/NPC_out[30] ,
         \DP/NPC_out[29] , \DP/NPC_out[28] , \DP/NPC_out[27] ,
         \DP/NPC_out[26] , \DP/NPC_out[25] , \DP/NPC_out[24] ,
         \DP/NPC_out[23] , \DP/NPC_out[22] , \DP/NPC_out[21] ,
         \DP/NPC_out[20] , \DP/NPC_out[19] , \DP/NPC_out[18] ,
         \DP/NPC_out[17] , \DP/NPC_out[16] , \DP/NPC_out[15] ,
         \DP/NPC_out[14] , \DP/NPC_out[13] , \DP/NPC_out[12] ,
         \DP/NPC_out[11] , \DP/NPC_out[10] , \DP/NPC_out[9] , \DP/NPC_out[8] ,
         \DP/NPC_out[7] , \DP/NPC_out[6] , \DP/NPC_out[5] , \DP/NPC_out[4] ,
         \DP/NPC_out[3] , \DP/NPC_out[2] , \DP/NPC_out[1] , \DP/NPC_out[0] ,
         \DP/RF_EN , \DP/NPC1[31] , \DP/NPC1[30] , \DP/NPC1[29] ,
         \DP/NPC1[28] , \DP/NPC1[27] , \DP/NPC1[26] , \DP/NPC1[25] ,
         \DP/NPC1[24] , \DP/NPC1[23] , \DP/NPC1[22] , \DP/NPC1[20] ,
         \DP/NPC1[19] , \DP/NPC1[18] , \DP/NPC1[17] , \DP/NPC1[16] ,
         \DP/NPC1[15] , \DP/NPC1[14] , \DP/NPC1[13] , \DP/NPC1[12] ,
         \DP/NPC1[11] , \DP/NPC1[10] , \DP/NPC1[9] , \DP/NPC1[8] ,
         \DP/NPC1[7] , \DP/NPC1[6] , \DP/NPC1[5] , \DP/NPC1[4] , \DP/NPC1[3] ,
         \DP/NPC1[2] , \DP/NPC1[1] , \DP/NPC1[0] , \DP/OUTCOME , \IR/N34 ,
         \IR/N33 , \IR/N32 , \IR/N31 , \IR/N30 , \IR/N29 , \IR/N28 , \IR/N27 ,
         \IR/N26 , \IR/N25 , \IR/N24 , \IR/N23 , \IR/N22 , \IR/N21 , \IR/N20 ,
         \IR/N19 , \IR/N18 , \IR/N17 , \IR/N16 , \IR/N15 , \IR/N14 , \IR/N13 ,
         \IR/N12 , \IR/N11 , \IR/N10 , \IR/N9 , \IR/N8 , \IR/N7 , \IR/N6 ,
         \IR/N5 , \IR/N4 , \IR/N3 , \DP/RegRD1/net7086 , \DP/RegRD1/N7 ,
         \DP/RegRD1/N6 , \DP/RegRD1/N5 , \DP/RegRD1/N4 , \DP/RegRD1/N3 ,
         \DP/RegRD1/N2 , \DP/FFDBRANCH/net7032 , \DP/FFDBRANCH/N3 ,
         \DP/FFDBRANCH/N2 , \DP/RegNPC/net7068 , \DP/RegNPC1/net7068 ,
         \DP/RegNPC1/N34 , \DP/RegNPC1/N33 , \DP/RegNPC1/N32 ,
         \DP/RegNPC1/N31 , \DP/RegNPC1/N30 , \DP/RegNPC1/N29 ,
         \DP/RegNPC1/N28 , \DP/RegNPC1/N27 , \DP/RegNPC1/N26 ,
         \DP/RegNPC1/N25 , \DP/RegNPC1/N24 , \DP/RegNPC1/N23 ,
         \DP/RegNPC1/N22 , \DP/RegNPC1/N21 , \DP/RegNPC1/N20 ,
         \DP/RegNPC1/N19 , \DP/RegNPC1/N18 , \DP/RegNPC1/N17 ,
         \DP/RegNPC1/N16 , \DP/RegNPC1/N15 , \DP/RegNPC1/N14 ,
         \DP/RegNPC1/N13 , \DP/RegNPC1/N12 , \DP/RegNPC1/N11 ,
         \DP/RegNPC1/N10 , \DP/RegNPC1/N9 , \DP/RegNPC1/N8 , \DP/RegNPC1/N7 ,
         \DP/RegNPC1/N6 , \DP/RegNPC1/N5 , \DP/RegNPC1/N4 , \DP/RegNPC1/N3 ,
         \DP/RegNPC1/N2 , \DP/RegA/net7068 , \DP/RegA/N34 , \DP/RegA/N33 ,
         \DP/RegA/N32 , \DP/RegA/N31 , \DP/RegA/N30 , \DP/RegA/N29 ,
         \DP/RegA/N28 , \DP/RegA/N27 , \DP/RegA/N26 , \DP/RegA/N25 ,
         \DP/RegA/N24 , \DP/RegA/N23 , \DP/RegA/N22 , \DP/RegA/N21 ,
         \DP/RegA/N20 , \DP/RegA/N19 , \DP/RegA/N18 , \DP/RegA/N17 ,
         \DP/RegA/N16 , \DP/RegA/N15 , \DP/RegA/N14 , \DP/RegA/N13 ,
         \DP/RegA/N12 , \DP/RegA/N11 , \DP/RegA/N10 , \DP/RegA/N9 ,
         \DP/RegA/N8 , \DP/RegA/N7 , \DP/RegA/N6 , \DP/RegA/N5 , \DP/RegA/N4 ,
         \DP/RegA/N3 , \DP/RegA/N2 , \DP/RegB/net7068 , \DP/RegB/N34 ,
         \DP/RegB/N33 , \DP/RegB/N32 , \DP/RegB/N31 , \DP/RegB/N30 ,
         \DP/RegB/N29 , \DP/RegB/N28 , \DP/RegB/N27 , \DP/RegB/N26 ,
         \DP/RegB/N25 , \DP/RegB/N24 , \DP/RegB/N23 , \DP/RegB/N22 ,
         \DP/RegB/N21 , \DP/RegB/N20 , \DP/RegB/N19 , \DP/RegB/N18 ,
         \DP/RegB/N17 , \DP/RegB/N16 , \DP/RegB/N15 , \DP/RegB/N14 ,
         \DP/RegB/N13 , \DP/RegB/N12 , \DP/RegB/N11 , \DP/RegB/N10 ,
         \DP/RegB/N9 , \DP/RegB/N8 , \DP/RegB/N7 , \DP/RegB/N6 , \DP/RegB/N5 ,
         \DP/RegB/N4 , \DP/RegB/N3 , \DP/RegB/N2 , \DP/RegIMM/net7068 ,
         \DP/RegIMM/N34 , \DP/RegIMM/N27 , \DP/RegIMM/N26 , \DP/RegIMM/N25 ,
         \DP/RegIMM/N24 , \DP/RegIMM/N23 , \DP/RegIMM/N22 , \DP/RegIMM/N21 ,
         \DP/RegIMM/N20 , \DP/RegIMM/N19 , \DP/RegIMM/N13 , \DP/RegIMM/N12 ,
         \DP/RegIMM/N11 , \DP/RegIMM/N10 , \DP/RegIMM/N9 , \DP/RegIMM/N8 ,
         \DP/RegIMM/N7 , \DP/RegIMM/N6 , \DP/RegIMM/N5 , \DP/RegIMM/N4 ,
         \DP/RegIMM/N3 , \DP/RegIMM/N2 , \DP/RegA1/net7068 , \DP/RegA1/N34 ,
         \DP/RegA1/N33 , \DP/RegA1/N32 , \DP/RegA1/N31 , \DP/RegA1/N30 ,
         \DP/RegA1/N29 , \DP/RegA1/N28 , \DP/RegA1/N27 , \DP/RegA1/N26 ,
         \DP/RegA1/N25 , \DP/RegA1/N24 , \DP/RegA1/N23 , \DP/RegA1/N22 ,
         \DP/RegA1/N21 , \DP/RegA1/N20 , \DP/RegA1/N19 , \DP/RegA1/N18 ,
         \DP/RegA1/N17 , \DP/RegA1/N16 , \DP/RegA1/N15 , \DP/RegA1/N14 ,
         \DP/RegA1/N13 , \DP/RegA1/N12 , \DP/RegA1/N11 , \DP/RegA1/N10 ,
         \DP/RegA1/N9 , \DP/RegA1/N8 , \DP/RegA1/N7 , \DP/RegA1/N6 ,
         \DP/RegA1/N5 , \DP/RegA1/N4 , \DP/RegA1/N3 , \DP/RegA1/N2 ,
         \DP/FFDJL1/N3 , \DP/FFDJREG/N3 , \DP/RegNPC2/net7068 ,
         \DP/RegNPC2/N34 , \DP/RegNPC2/N33 , \DP/RegNPC2/N32 ,
         \DP/RegNPC2/N31 , \DP/RegNPC2/N30 , \DP/RegNPC2/N29 ,
         \DP/RegNPC2/N28 , \DP/RegNPC2/N27 , \DP/RegNPC2/N26 ,
         \DP/RegNPC2/N25 , \DP/RegNPC2/N24 , \DP/RegNPC2/N23 ,
         \DP/RegNPC2/N22 , \DP/RegNPC2/N21 , \DP/RegNPC2/N20 ,
         \DP/RegNPC2/N19 , \DP/RegNPC2/N18 , \DP/RegNPC2/N17 ,
         \DP/RegNPC2/N16 , \DP/RegNPC2/N15 , \DP/RegNPC2/N14 ,
         \DP/RegNPC2/N13 , \DP/RegNPC2/N12 , \DP/RegNPC2/N11 ,
         \DP/RegNPC2/N10 , \DP/RegNPC2/N9 , \DP/RegNPC2/N8 , \DP/RegNPC2/N7 ,
         \DP/RegNPC2/N6 , \DP/RegNPC2/N5 , \DP/RegNPC2/N4 , \DP/RegNPC2/N3 ,
         \DP/RegNPC2/N2 , \DP/RegALU1/net7068 , \DP/RegALU1/N34 ,
         \DP/RegALU1/N33 , \DP/RegALU1/N32 , \DP/RegALU1/N31 ,
         \DP/RegALU1/N30 , \DP/RegALU1/N29 , \DP/RegALU1/N28 ,
         \DP/RegALU1/N27 , \DP/RegALU1/N26 , \DP/RegALU1/N25 ,
         \DP/RegALU1/N24 , \DP/RegALU1/N23 , \DP/RegALU1/N22 ,
         \DP/RegALU1/N21 , \DP/RegALU1/N20 , \DP/RegALU1/N19 ,
         \DP/RegALU1/N18 , \DP/RegALU1/N17 , \DP/RegALU1/N16 ,
         \DP/RegALU1/N15 , \DP/RegALU1/N14 , \DP/RegALU1/N13 ,
         \DP/RegALU1/N12 , \DP/RegALU1/N11 , \DP/RegALU1/N10 , \DP/RegALU1/N9 ,
         \DP/RegALU1/N8 , \DP/RegALU1/N7 , \DP/RegALU1/N6 , \DP/RegALU1/N5 ,
         \DP/RegALU1/N4 , \DP/RegALU1/N3 , \DP/RegALU1/N2 , \DP/RegME/net7068 ,
         \DP/RegME/N34 , \DP/RegME/N33 , \DP/RegME/N32 , \DP/RegME/N31 ,
         \DP/RegME/N30 , \DP/RegME/N29 , \DP/RegME/N28 , \DP/RegME/N27 ,
         \DP/RegME/N26 , \DP/RegME/N25 , \DP/RegME/N24 , \DP/RegME/N23 ,
         \DP/RegME/N22 , \DP/RegME/N21 , \DP/RegME/N20 , \DP/RegME/N19 ,
         \DP/RegME/N18 , \DP/RegME/N17 , \DP/RegME/N16 , \DP/RegME/N15 ,
         \DP/RegME/N14 , \DP/RegME/N13 , \DP/RegME/N12 , \DP/RegME/N11 ,
         \DP/RegME/N10 , \DP/RegME/N9 , \DP/RegME/N8 , \DP/RegME/N7 ,
         \DP/RegME/N6 , \DP/RegME/N5 , \DP/RegME/N4 , \DP/RegME/N3 ,
         \DP/RegME/N2 , \DP/RegRD2/net7086 , \DP/RegRD2/N7 , \DP/RegRD2/N6 ,
         \DP/RegRD2/N5 , \DP/RegRD2/N4 , \DP/RegRD2/N2 , \DP/RegALU2/net7068 ,
         \DP/RegALU2/N34 , \DP/RegALU2/N33 , \DP/RegALU2/N32 ,
         \DP/RegALU2/N31 , \DP/RegALU2/N30 , \DP/RegALU2/N29 ,
         \DP/RegALU2/N28 , \DP/RegALU2/N27 , \DP/RegALU2/N26 ,
         \DP/RegALU2/N25 , \DP/RegALU2/N24 , \DP/RegALU2/N23 ,
         \DP/RegALU2/N22 , \DP/RegALU2/N21 , \DP/RegALU2/N20 ,
         \DP/RegALU2/N19 , \DP/RegALU2/N18 , \DP/RegALU2/N17 ,
         \DP/RegALU2/N16 , \DP/RegALU2/N15 , \DP/RegALU2/N14 ,
         \DP/RegALU2/N13 , \DP/RegALU2/N12 , \DP/RegALU2/N11 ,
         \DP/RegALU2/N10 , \DP/RegALU2/N9 , \DP/RegALU2/N8 , \DP/RegALU2/N7 ,
         \DP/RegALU2/N6 , \DP/RegALU2/N5 , \DP/RegALU2/N4 , \DP/RegALU2/N3 ,
         \DP/RegALU2/N2 , \DP/RegLMD/net7068 , \DP/RegLMD/N34 ,
         \DP/RegLMD/N33 , \DP/RegLMD/N32 , \DP/RegLMD/N31 , \DP/RegLMD/N30 ,
         \DP/RegLMD/N29 , \DP/RegLMD/N28 , \DP/RegLMD/N27 , \DP/RegLMD/N26 ,
         \DP/RegLMD/N25 , \DP/RegLMD/N23 , \DP/RegLMD/N22 , \DP/RegLMD/N21 ,
         \DP/RegLMD/N20 , \DP/RegLMD/N19 , \DP/RegLMD/N18 , \DP/RegLMD/N17 ,
         \DP/RegLMD/N16 , \DP/RegLMD/N15 , \DP/RegLMD/N14 , \DP/RegLMD/N13 ,
         \DP/RegLMD/N12 , \DP/RegLMD/N11 , \DP/RegLMD/N10 , \DP/RegLMD/N9 ,
         \DP/RegLMD/N8 , \DP/RegLMD/N7 , \DP/RegLMD/N6 , \DP/RegLMD/N5 ,
         \DP/RegLMD/N4 , \DP/RegLMD/N3 , \DP/RegLMD/N2 , \DP/RegRD3/net7086 ,
         \DP/RegRD3/N7 , \DP/RegRD3/N6 , \DP/RegRD3/N5 , \DP/RegRD3/N4 ,
         \DP/RegRD3/N3 , \DP/RegRD3/N2 , \DP/FFDJL2/net7032 , \DP/FFDJL2/N3 ,
         \DP/FFDJL2/N2 , \DP/RegNPC3/net7068 , \DP/RegNPC3/N34 ,
         \DP/RegNPC3/N33 , \DP/RegNPC3/N32 , \DP/RegNPC3/N31 ,
         \DP/RegNPC3/N30 , \DP/RegNPC3/N29 , \DP/RegNPC3/N28 ,
         \DP/RegNPC3/N27 , \DP/RegNPC3/N26 , \DP/RegNPC3/N25 ,
         \DP/RegNPC3/N24 , \DP/RegNPC3/N23 , \DP/RegNPC3/N22 ,
         \DP/RegNPC3/N21 , \DP/RegNPC3/N20 , \DP/RegNPC3/N19 ,
         \DP/RegNPC3/N18 , \DP/RegNPC3/N17 , \DP/RegNPC3/N16 ,
         \DP/RegNPC3/N15 , \DP/RegNPC3/N14 , \DP/RegNPC3/N13 ,
         \DP/RegNPC3/N12 , \DP/RegNPC3/N11 , \DP/RegNPC3/N10 , \DP/RegNPC3/N9 ,
         \DP/RegNPC3/N8 , \DP/RegNPC3/N7 , \DP/RegNPC3/N6 , \DP/RegNPC3/N5 ,
         \DP/RegNPC3/N4 , \DP/RegNPC3/N3 , \DP/RegNPC3/N2 , \DP/RegFB/N4 ,
         \DP/RegFB/N3 , \DP/RegFC/N5 , \DP/RegFC/N4 , \DP/RegFC/N3 ,
         \DP/FFDFD/N3 , n12, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n53, n57, n58, n59, n62, n69, n72, n73, n75, n76, n77, n181, n184,
         n186, n188, n190, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n628, n629, n630, n631, n632,
         n633, n634, n635, n638, n639, n640, n641, n645, n648, n652, n653,
         n654, n655, n656, n657, n659, n660, n661, n662, n663, n665, n666,
         n668, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n686, n687, n688, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n706, n707, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n721, n722,
         n723, n724, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n929, n933,
         n935, n936, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1015,
         n1016, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1163, n1164, n1165, n1167, n1170, n1171, n1172,
         n1173, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1208, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1274, n1275, n1276, n1277,
         n1278, n1280, n1282, n1284, n1285, n1286, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1400, n1401, n1402, n1403, n1404, n1407, n1408,
         n1409, n1410, n1411, n1412, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1476, n1477, n1478, n1479, n1480, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1492, n1493, n1494, n1495, n1497,
         n1498, n1499, n1500, n1501, n1506, n1507, n1508, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1594, n1595, n1596,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1829, n1830, n1839, n1840,
         n1843, n1844, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862;
  wire   [31:12] w_PC_OUT;
  wire   [31:0] IR_OUT;
  wire   [4:0] w_ALU_OPCODE;
  wire   [2:0] w_STORE_SIZE;
  wire   [2:0] w_LOAD_SIZE;
  assign \DP/LOAD8[7]  = DRAM_DATA_IN[7];
  assign \DP/LOAD8[6]  = DRAM_DATA_IN[6];
  assign \DP/LOAD8[5]  = DRAM_DATA_IN[5];
  assign \DP/LOAD8[4]  = DRAM_DATA_IN[4];
  assign \DP/LOAD8[3]  = DRAM_DATA_IN[3];
  assign \DP/LOAD8[2]  = DRAM_DATA_IN[2];
  assign \DP/LOAD8[1]  = DRAM_DATA_IN[1];
  assign \DP/LOAD8[0]  = DRAM_DATA_IN[0];
  assign \DP/LOAD16[15]  = DRAM_DATA_IN[15];
  assign \DP/LOAD16[14]  = DRAM_DATA_IN[14];
  assign \DP/LOAD16[13]  = DRAM_DATA_IN[13];
  assign \DP/LOAD16[12]  = DRAM_DATA_IN[12];
  assign \DP/LOAD16[11]  = DRAM_DATA_IN[11];
  assign \DP/LOAD16[10]  = DRAM_DATA_IN[10];
  assign \DP/LOAD16[9]  = DRAM_DATA_IN[9];
  assign \DP/LOAD16[8]  = DRAM_DATA_IN[8];
  assign IROM_ADDR[6] = \DP/NPC1[6] ;
  assign IROM_ADDR[4] = \DP/NPC1[4] ;
  assign IROM_ADDR[3] = \DP/NPC1[3] ;
  assign IROM_ADDR[2] = \DP/NPC1[2] ;
  assign IROM_ADDR[1] = \DP/NPC1[1] ;

  DFF_X1 \CU/IF_EN_reg  ( .D(n641), .CK(CLK), .QN(w_IF_EN) );
  DFF_X1 \IR/DOUT_reg[0]  ( .D(\IR/N3 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[0]), .QN(n1447) );
  DFF_X1 \IR/DOUT_reg[1]  ( .D(\IR/N4 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[1]) );
  DFF_X1 \IR/DOUT_reg[2]  ( .D(\IR/N5 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[2]) );
  DFF_X1 \IR/DOUT_reg[3]  ( .D(\IR/N6 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[3]) );
  DFF_X1 \IR/DOUT_reg[4]  ( .D(\IR/N7 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[4]), .QN(n595) );
  DFF_X1 \IR/DOUT_reg[5]  ( .D(\IR/N8 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[5]) );
  DFF_X1 \IR/DOUT_reg[6]  ( .D(\IR/N9 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[6]) );
  DFF_X1 \IR/DOUT_reg[7]  ( .D(\IR/N10 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[7]) );
  DFF_X1 \IR/DOUT_reg[8]  ( .D(\IR/N11 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[8]) );
  DFF_X1 \IR/DOUT_reg[9]  ( .D(\IR/N12 ), .CK(\DP/RegNPC/net7068 ), .Q(n1468), 
        .QN(n600) );
  DFF_X1 \IR/DOUT_reg[10]  ( .D(\IR/N13 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[10]) );
  DFF_X1 \IR/DOUT_reg[11]  ( .D(\IR/N14 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[11]) );
  DFF_X1 \IR/DOUT_reg[12]  ( .D(\IR/N15 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[12]) );
  DFF_X1 \IR/DOUT_reg[13]  ( .D(\IR/N16 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[13]) );
  DFF_X1 \IR/DOUT_reg[14]  ( .D(\IR/N17 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[14]) );
  DFF_X1 \IR/DOUT_reg[15]  ( .D(\IR/N18 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[15]) );
  DFF_X1 \IR/DOUT_reg[16]  ( .D(\IR/N19 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[16]) );
  DFF_X1 \IR/DOUT_reg[17]  ( .D(\IR/N20 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[17]) );
  DFF_X1 \IR/DOUT_reg[18]  ( .D(\IR/N21 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[18]) );
  DFF_X1 \IR/DOUT_reg[19]  ( .D(\IR/N22 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[19]) );
  DFF_X1 \IR/DOUT_reg[20]  ( .D(\IR/N23 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[20]) );
  DFF_X1 \IR/DOUT_reg[21]  ( .D(\IR/N24 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[21]) );
  DFF_X1 \IR/DOUT_reg[22]  ( .D(\IR/N25 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[22]) );
  DFF_X1 \IR/DOUT_reg[23]  ( .D(\IR/N26 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[23]) );
  DFF_X1 \IR/DOUT_reg[24]  ( .D(\IR/N27 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[24]) );
  DFF_X1 \IR/DOUT_reg[25]  ( .D(\IR/N28 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[25]) );
  DFF_X1 \IR/DOUT_reg[26]  ( .D(\IR/N29 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[26]), .QN(n586) );
  DFF_X1 \IR/DOUT_reg[27]  ( .D(\IR/N30 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[27]) );
  DFF_X1 \IR/DOUT_reg[28]  ( .D(\IR/N31 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[28]) );
  DFF_X1 \IR/DOUT_reg[29]  ( .D(\IR/N32 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[29]) );
  DFF_X1 \IR/DOUT_reg[30]  ( .D(\IR/N33 ), .CK(\DP/RegNPC/net7068 ), .Q(n592), 
        .QN(n62) );
  DFF_X1 \IR/DOUT_reg[31]  ( .D(\IR/N34 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IR_OUT[31]) );
  DFF_X1 \CU/cw1_reg[17]  ( .D(n12), .CK(CLK), .Q(n590) );
  DFF_X1 \CU/cw1_reg[19]  ( .D(\CU/N59 ), .CK(CLK), .Q(w_JUMP_EQ) );
  DFF_X1 \CU/cw1_reg[16]  ( .D(\CU/N56 ), .CK(CLK), .Q(w_RegME_LATCH_EN) );
  DFF_X1 \CU/cw1_reg[13]  ( .D(\CU/N56 ), .CK(CLK), .Q(\CU/cw1[13] ) );
  DFF_X1 \CU/cw1_reg[12]  ( .D(\CU/N52 ), .CK(CLK), .Q(\CU/cw1[12] ) );
  DFF_X1 \CU/cw2_reg[12]  ( .D(\CU/N76 ), .CK(CLK), .QN(n57) );
  DFF_X1 \CU/cw1_reg[11]  ( .D(\CU/N51 ), .CK(CLK), .Q(\CU/cw1[11] ) );
  DFF_X1 \CU/cw1_reg[10]  ( .D(\CU/N50 ), .CK(CLK), .Q(\CU/cw1[10] ) );
  DFF_X1 \CU/cw1_reg[20]  ( .D(\CU/N60 ), .CK(CLK), .QN(n59) );
  DFF_X1 \CU/cw1_reg[18]  ( .D(\CU/N58 ), .CK(CLK), .QN(n58) );
  DFF_X1 \CU/cw1_reg[9]  ( .D(\CU/N49 ), .CK(CLK), .Q(\CU/cw1[9] ) );
  DFF_X1 \CU/cw1_reg[8]  ( .D(\CU/N48 ), .CK(CLK), .Q(\CU/cw1[8] ) );
  DFF_X1 \CU/cw1_reg[7]  ( .D(\CU/N47 ), .CK(CLK), .Q(\CU/cw1[7] ) );
  DFF_X1 \CU/cw1_reg[6]  ( .D(\CU/N46 ), .CK(CLK), .Q(\CU/cw1[6] ) );
  DFF_X1 \CU/cw1_reg[14]  ( .D(\CU/N54 ), .CK(CLK), .Q(\CU/cw1[14] ) );
  DFF_X1 \CU/aluOpcode1_reg[3]  ( .D(\CU/N88 ), .CK(CLK), .Q(w_ALU_OPCODE[3])
         );
  DFF_X1 \CU/aluOpcode1_reg[0]  ( .D(\CU/N85 ), .CK(CLK), .Q(w_ALU_OPCODE[0])
         );
  DFF_X1 \CU/aluOpcode1_reg[2]  ( .D(\CU/N87 ), .CK(CLK), .Q(w_ALU_OPCODE[2])
         );
  DFF_X1 \CU/aluOpcode1_reg[1]  ( .D(\CU/N86 ), .CK(CLK), .Q(w_ALU_OPCODE[1])
         );
  DFF_X1 \CU/aluOpcode1_reg[4]  ( .D(\CU/N89 ), .CK(CLK), .Q(w_ALU_OPCODE[4])
         );
  DFF_X1 \CU/cw1_reg[23]  ( .D(\CU/N63 ), .CK(CLK), .Q(w_EX_EN) );
  DFF_X1 \CU/cw1_reg[15]  ( .D(n1486), .CK(CLK), .Q(w_RegRD2_LATCH_EN) );
  DFF_X1 \CU/cw1_reg[3]  ( .D(n1486), .CK(CLK), .Q(\CU/cw1[3] ) );
  DFF_X1 \CU/cw2_reg[0]  ( .D(\CU/N64 ), .CK(CLK), .QN(n601) );
  DFF_X1 \CU/cw1_reg[5]  ( .D(\CU/N45 ), .CK(CLK), .Q(\CU/cw1[5] ) );
  DFF_X1 \DP/RegRD1/DOUT_reg[0]  ( .D(\DP/RegRD1/N3 ), .CK(\DP/RegRD1/net7086 ), .Q(\DP/RD1[0] ) );
  DFF_X1 \DP/RegRD1/DOUT_reg[3]  ( .D(\DP/RegRD1/N6 ), .CK(\DP/RegRD1/net7086 ), .Q(\DP/RD1[3] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[0]  ( .D(\DP/RegIMM/N3 ), .CK(\DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[0] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[1]  ( .D(\DP/RegIMM/N4 ), .CK(\DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[1] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[2]  ( .D(\DP/RegIMM/N5 ), .CK(\DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[2] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[3]  ( .D(\DP/RegIMM/N6 ), .CK(\DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[3] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[4]  ( .D(\DP/RegIMM/N7 ), .CK(\DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[4] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[5]  ( .D(\DP/RegIMM/N8 ), .CK(\DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[5] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[6]  ( .D(\DP/RegIMM/N9 ), .CK(\DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[6] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[7]  ( .D(\DP/RegIMM/N10 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[7] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[8]  ( .D(\DP/RegIMM/N11 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[8] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[9]  ( .D(\DP/RegIMM/N12 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[9] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[10]  ( .D(\DP/RegIMM/N13 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[10] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[11]  ( .D(n190), .CK(\DP/RegIMM/net7068 ), .QN(
        \DP/RegIMM_out[11] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[12]  ( .D(n188), .CK(\DP/RegIMM/net7068 ), .QN(
        \DP/RegIMM_out[12] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[13]  ( .D(n186), .CK(\DP/RegIMM/net7068 ), .QN(
        \DP/RegIMM_out[13] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[14]  ( .D(n184), .CK(\DP/RegIMM/net7068 ), .QN(
        \DP/RegIMM_out[14] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[15]  ( .D(n181), .CK(\DP/RegIMM/net7068 ), .QN(
        \DP/RegIMM_out[15] ) );
  DFF_X1 \DP/FFDJL1/Q_reg  ( .D(\DP/FFDJL1/N3 ), .CK(\DP/FFDJL2/net7032 ), .Q(
        \DP/JL1 ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[0]  ( .D(\DP/RegLMD/N3 ), .CK(\DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[0] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[1]  ( .D(\DP/RegLMD/N4 ), .CK(\DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[1] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[2]  ( .D(\DP/RegLMD/N5 ), .CK(\DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[2] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[3]  ( .D(\DP/RegLMD/N6 ), .CK(\DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[3] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[4]  ( .D(\DP/RegLMD/N7 ), .CK(\DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[4] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[5]  ( .D(\DP/RegLMD/N8 ), .CK(\DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[5] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[6]  ( .D(\DP/RegLMD/N9 ), .CK(\DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[6] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[7]  ( .D(\DP/RegLMD/N10 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[7] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[8]  ( .D(\DP/RegLMD/N11 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[8] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[9]  ( .D(\DP/RegLMD/N12 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[9] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[10]  ( .D(\DP/RegLMD/N13 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[10] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[11]  ( .D(\DP/RegLMD/N14 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[11] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[12]  ( .D(\DP/RegLMD/N15 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[12] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[13]  ( .D(\DP/RegLMD/N16 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[13] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[14]  ( .D(\DP/RegLMD/N17 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[14] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[15]  ( .D(\DP/RegLMD/N18 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[15] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[16]  ( .D(\DP/RegLMD/N19 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[16] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[17]  ( .D(\DP/RegLMD/N20 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[17] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[18]  ( .D(\DP/RegLMD/N21 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[18] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[19]  ( .D(\DP/RegLMD/N22 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[19] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[20]  ( .D(\DP/RegLMD/N23 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[20] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[22]  ( .D(\DP/RegLMD/N25 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[22] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[23]  ( .D(\DP/RegLMD/N26 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[23] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[24]  ( .D(\DP/RegLMD/N27 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[24] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[25]  ( .D(\DP/RegLMD/N28 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[25] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[26]  ( .D(\DP/RegLMD/N29 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[26] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[27]  ( .D(\DP/RegLMD/N30 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[27] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[28]  ( .D(\DP/RegLMD/N31 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[28] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[29]  ( .D(\DP/RegLMD/N32 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[29] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[30]  ( .D(\DP/RegLMD/N33 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[30] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[31]  ( .D(\DP/RegLMD/N34 ), .CK(
        \DP/RegLMD/net7068 ), .Q(\DP/RegLMD_out[31] ) );
  DFF_X1 \DP/RegRD3/DOUT_reg[4]  ( .D(\DP/RegRD3/N7 ), .CK(\DP/RegRD3/net7086 ), .Q(\DP/RD3[4] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[18]  ( .D(\DP/RegA1/N21 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[18] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[6]  ( .D(\PC/N9 ), .CK(n635), .Q(\DP/NPC1[6] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[6]  ( .D(\DP/RegNPC1/N9 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[6] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[6]  ( .D(\DP/RegNPC2/N9 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[6] ) );
  DFF_X1 \DP/RegB/DOUT_reg[0]  ( .D(\DP/RegB/N3 ), .CK(\DP/RegB/net7068 ), .Q(
        \DP/RegB_out[0] ) );
  DFF_X1 \DP/RegME/DOUT_reg[0]  ( .D(\DP/RegME/N3 ), .CK(\DP/RegME/net7068 ), 
        .QN(n611) );
  DFF_X1 \DP/RegB/DOUT_reg[1]  ( .D(\DP/RegB/N4 ), .CK(\DP/RegB/net7068 ), .Q(
        \DP/RegB_out[1] ) );
  DFF_X1 \DP/RegME/DOUT_reg[1]  ( .D(\DP/RegME/N4 ), .CK(\DP/RegME/net7068 ), 
        .QN(n612) );
  DFF_X1 \DP/RegB/DOUT_reg[2]  ( .D(\DP/RegB/N5 ), .CK(\DP/RegB/net7068 ), .Q(
        \DP/RegB_out[2] ) );
  DFF_X1 \DP/RegME/DOUT_reg[2]  ( .D(\DP/RegME/N5 ), .CK(\DP/RegME/net7068 ), 
        .QN(n613) );
  DFF_X1 \DP/RegB/DOUT_reg[3]  ( .D(\DP/RegB/N6 ), .CK(\DP/RegB/net7068 ), .Q(
        \DP/RegB_out[3] ) );
  DFF_X1 \DP/RegME/DOUT_reg[3]  ( .D(\DP/RegME/N6 ), .CK(\DP/RegME/net7068 ), 
        .QN(n614) );
  DFF_X1 \DP/RegB/DOUT_reg[4]  ( .D(\DP/RegB/N7 ), .CK(\DP/RegB/net7068 ), .Q(
        \DP/RegB_out[4] ) );
  DFF_X1 \DP/RegME/DOUT_reg[4]  ( .D(\DP/RegME/N7 ), .CK(\DP/RegME/net7068 ), 
        .QN(n615) );
  DFF_X1 \DP/RegB/DOUT_reg[5]  ( .D(\DP/RegB/N8 ), .CK(\DP/RegB/net7068 ), .Q(
        \DP/RegB_out[5] ) );
  DFF_X1 \DP/RegME/DOUT_reg[5]  ( .D(\DP/RegME/N8 ), .CK(\DP/RegME/net7068 ), 
        .QN(n616) );
  DFF_X1 \DP/RegB/DOUT_reg[6]  ( .D(\DP/RegB/N9 ), .CK(\DP/RegB/net7068 ), .Q(
        \DP/RegB_out[6] ) );
  DFF_X1 \DP/RegME/DOUT_reg[6]  ( .D(\DP/RegME/N9 ), .CK(\DP/RegME/net7068 ), 
        .QN(n617) );
  DFF_X1 \DP/RegB/DOUT_reg[7]  ( .D(\DP/RegB/N10 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[7] ) );
  DFF_X1 \DP/RegB/DOUT_reg[8]  ( .D(\DP/RegB/N11 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[8] ) );
  DFF_X1 \DP/RegME/DOUT_reg[8]  ( .D(\DP/RegME/N11 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[8] ) );
  DFF_X1 \DP/RegB/DOUT_reg[9]  ( .D(\DP/RegB/N12 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[9] ) );
  DFF_X1 \DP/RegME/DOUT_reg[9]  ( .D(\DP/RegME/N12 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[9] ) );
  DFF_X1 \DP/RegB/DOUT_reg[10]  ( .D(\DP/RegB/N13 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[10] ) );
  DFF_X1 \DP/RegME/DOUT_reg[10]  ( .D(\DP/RegME/N13 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[10] ) );
  DFF_X1 \DP/RegB/DOUT_reg[11]  ( .D(\DP/RegB/N14 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[11] ) );
  DFF_X1 \DP/RegME/DOUT_reg[11]  ( .D(\DP/RegME/N14 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[11] ) );
  DFF_X1 \DP/RegB/DOUT_reg[12]  ( .D(\DP/RegB/N15 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[12] ) );
  DFF_X1 \DP/RegME/DOUT_reg[12]  ( .D(\DP/RegME/N15 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[12] ) );
  DFF_X1 \DP/RegB/DOUT_reg[13]  ( .D(\DP/RegB/N16 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[13] ) );
  DFF_X1 \DP/RegME/DOUT_reg[13]  ( .D(\DP/RegME/N16 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[13] ) );
  DFF_X1 \DP/RegB/DOUT_reg[14]  ( .D(\DP/RegB/N17 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[14] ) );
  DFF_X1 \DP/RegME/DOUT_reg[14]  ( .D(\DP/RegME/N17 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[14] ) );
  DFF_X1 \DP/RegB/DOUT_reg[15]  ( .D(\DP/RegB/N18 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[15] ) );
  DFF_X1 \DP/RegME/DOUT_reg[15]  ( .D(\DP/RegME/N18 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[15] ) );
  DFF_X1 \DP/RegB/DOUT_reg[16]  ( .D(\DP/RegB/N19 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[16] ) );
  DFF_X1 \DP/RegME/DOUT_reg[16]  ( .D(\DP/RegME/N19 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[16] ) );
  DFF_X1 \DP/RegB/DOUT_reg[17]  ( .D(\DP/RegB/N20 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[17] ) );
  DFF_X1 \DP/RegME/DOUT_reg[17]  ( .D(\DP/RegME/N20 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[17] ) );
  DFF_X1 \DP/RegB/DOUT_reg[18]  ( .D(\DP/RegB/N21 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[18] ) );
  DFF_X1 \DP/RegME/DOUT_reg[18]  ( .D(\DP/RegME/N21 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[18] ) );
  DFF_X1 \DP/RegB/DOUT_reg[19]  ( .D(\DP/RegB/N22 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[19] ) );
  DFF_X1 \DP/RegME/DOUT_reg[19]  ( .D(\DP/RegME/N22 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[19] ) );
  DFF_X1 \DP/RegB/DOUT_reg[20]  ( .D(\DP/RegB/N23 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[20] ) );
  DFF_X1 \DP/RegME/DOUT_reg[20]  ( .D(\DP/RegME/N23 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[20] ) );
  DFF_X1 \DP/RegB/DOUT_reg[21]  ( .D(\DP/RegB/N24 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[21] ) );
  DFF_X1 \DP/RegME/DOUT_reg[21]  ( .D(\DP/RegME/N24 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[21] ) );
  DFF_X1 \DP/RegB/DOUT_reg[22]  ( .D(\DP/RegB/N25 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[22] ) );
  DFF_X1 \DP/RegME/DOUT_reg[22]  ( .D(\DP/RegME/N25 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[22] ) );
  DFF_X1 \DP/RegB/DOUT_reg[23]  ( .D(\DP/RegB/N26 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[23] ) );
  DFF_X1 \DP/RegME/DOUT_reg[23]  ( .D(\DP/RegME/N26 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[23] ) );
  DFF_X1 \DP/RegB/DOUT_reg[24]  ( .D(\DP/RegB/N27 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[24] ) );
  DFF_X1 \DP/RegME/DOUT_reg[24]  ( .D(\DP/RegME/N27 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[24] ) );
  DFF_X1 \DP/RegB/DOUT_reg[25]  ( .D(\DP/RegB/N28 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[25] ) );
  DFF_X1 \DP/RegME/DOUT_reg[25]  ( .D(\DP/RegME/N28 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[25] ) );
  DFF_X1 \DP/RegB/DOUT_reg[26]  ( .D(\DP/RegB/N29 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[26] ) );
  DFF_X1 \DP/RegME/DOUT_reg[26]  ( .D(\DP/RegME/N29 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[26] ) );
  DFF_X1 \DP/RegB/DOUT_reg[27]  ( .D(\DP/RegB/N30 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[27] ) );
  DFF_X1 \DP/RegME/DOUT_reg[27]  ( .D(\DP/RegME/N30 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[27] ) );
  DFF_X1 \DP/RegB/DOUT_reg[28]  ( .D(\DP/RegB/N31 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[28] ) );
  DFF_X1 \DP/RegME/DOUT_reg[28]  ( .D(\DP/RegME/N31 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[28] ) );
  DFF_X1 \DP/RegB/DOUT_reg[29]  ( .D(\DP/RegB/N32 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[29] ) );
  DFF_X1 \DP/RegME/DOUT_reg[29]  ( .D(\DP/RegME/N32 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[29] ) );
  DFF_X1 \DP/RegB/DOUT_reg[30]  ( .D(\DP/RegB/N33 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[30] ) );
  DFF_X1 \DP/RegME/DOUT_reg[30]  ( .D(\DP/RegME/N33 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[30] ) );
  DFF_X1 \DP/RegB/DOUT_reg[31]  ( .D(\DP/RegB/N34 ), .CK(\DP/RegB/net7068 ), 
        .Q(\DP/RegB_out[31] ) );
  DFF_X1 \DP/RegME/DOUT_reg[31]  ( .D(\DP/RegME/N34 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[31] ) );
  DFF_X1 \DP/RegA/DOUT_reg[0]  ( .D(\DP/RegA/N3 ), .CK(\DP/RegA/net7068 ), .Q(
        \DP/RegA_out[0] ), .QN(n1427) );
  DFF_X1 \DP/RegA/DOUT_reg[1]  ( .D(\DP/RegA/N4 ), .CK(\DP/RegA/net7068 ), .Q(
        \DP/RegA_out[1] ), .QN(n1395) );
  DFF_X1 \DP/RegA/DOUT_reg[2]  ( .D(\DP/RegA/N5 ), .CK(\DP/RegA/net7068 ), .Q(
        \DP/RegA_out[2] ), .QN(n1394) );
  DFF_X1 \DP/RegA/DOUT_reg[3]  ( .D(\DP/RegA/N6 ), .CK(\DP/RegA/net7068 ), .Q(
        \DP/RegA_out[3] ), .QN(n1445) );
  DFF_X1 \DP/RegA/DOUT_reg[4]  ( .D(\DP/RegA/N7 ), .CK(\DP/RegA/net7068 ), .Q(
        \DP/RegA_out[4] ), .QN(n1444) );
  DFF_X1 \DP/RegA/DOUT_reg[5]  ( .D(\DP/RegA/N8 ), .CK(\DP/RegA/net7068 ), .Q(
        \DP/RegA_out[5] ), .QN(n1443) );
  DFF_X1 \DP/RegA/DOUT_reg[6]  ( .D(\DP/RegA/N9 ), .CK(\DP/RegA/net7068 ), .Q(
        \DP/RegA_out[6] ), .QN(n1442) );
  DFF_X1 \DP/RegA/DOUT_reg[7]  ( .D(\DP/RegA/N10 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[7] ), .QN(n1410) );
  DFF_X1 \DP/RegA/DOUT_reg[8]  ( .D(\DP/RegA/N11 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[8] ), .QN(n1409) );
  DFF_X1 \DP/RegA/DOUT_reg[9]  ( .D(\DP/RegA/N12 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[9] ), .QN(n1408) );
  DFF_X1 \DP/RegA/DOUT_reg[10]  ( .D(\DP/RegA/N13 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[10] ), .QN(n1407) );
  DFF_X1 \DP/RegA/DOUT_reg[11]  ( .D(\DP/RegA/N14 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[11] ), .QN(n1385) );
  DFF_X1 \DP/RegA/DOUT_reg[12]  ( .D(\DP/RegA/N15 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[12] ), .QN(n1384) );
  DFF_X1 \DP/RegA/DOUT_reg[13]  ( .D(\DP/RegA/N16 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[13] ), .QN(n1383) );
  DFF_X1 \DP/RegA/DOUT_reg[14]  ( .D(\DP/RegA/N17 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[14] ), .QN(n1382) );
  DFF_X1 \DP/RegA/DOUT_reg[15]  ( .D(\DP/RegA/N18 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[15] ) );
  DFF_X1 \DP/RegA/DOUT_reg[16]  ( .D(\DP/RegA/N19 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[16] ) );
  DFF_X1 \DP/RegA/DOUT_reg[17]  ( .D(\DP/RegA/N20 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[17] ) );
  DFF_X1 \DP/RegA/DOUT_reg[18]  ( .D(\DP/RegA/N21 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[18] ) );
  DFF_X1 \DP/RegA/DOUT_reg[19]  ( .D(\DP/RegA/N22 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[19] ), .QN(n1404) );
  DFF_X1 \DP/RegA/DOUT_reg[20]  ( .D(\DP/RegA/N23 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[20] ), .QN(n1403) );
  DFF_X1 \DP/RegA/DOUT_reg[21]  ( .D(\DP/RegA/N24 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[21] ), .QN(n1402) );
  DFF_X1 \DP/RegA/DOUT_reg[22]  ( .D(\DP/RegA/N25 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[22] ), .QN(n1401) );
  DFF_X1 \DP/RegA/DOUT_reg[23]  ( .D(\DP/RegA/N26 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[23] ), .QN(n1437) );
  DFF_X1 \DP/RegA/DOUT_reg[24]  ( .D(\DP/RegA/N27 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[24] ), .QN(n1436) );
  DFF_X1 \DP/RegA/DOUT_reg[25]  ( .D(\DP/RegA/N28 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[25] ), .QN(n1435) );
  DFF_X1 \DP/RegA/DOUT_reg[26]  ( .D(\DP/RegA/N29 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[26] ), .QN(n1434) );
  DFF_X1 \DP/RegA/DOUT_reg[27]  ( .D(\DP/RegA/N30 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[27] ), .QN(n1426) );
  DFF_X1 \DP/RegA/DOUT_reg[28]  ( .D(\DP/RegA/N31 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[28] ), .QN(n1425) );
  DFF_X1 \DP/RegA/DOUT_reg[29]  ( .D(\DP/RegA/N32 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[29] ), .QN(n1424) );
  DFF_X1 \DP/RegA/DOUT_reg[30]  ( .D(\DP/RegA/N33 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[30] ), .QN(n1397) );
  DFF_X1 \DP/RegA/DOUT_reg[31]  ( .D(\DP/RegA/N34 ), .CK(\DP/RegA/net7068 ), 
        .Q(\DP/RegA_out[31] ), .QN(n1396) );
  DFF_X1 \DP/RegA1/DOUT_reg[31]  ( .D(\DP/RegA1/N34 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[31] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[31]  ( .D(\PC/N34 ), .CK(n635), .Q(\DP/NPC1[31] )
         );
  DFF_X1 \DP/RegNPC1/DOUT_reg[31]  ( .D(\DP/RegNPC1/N34 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[31] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[0]  ( .D(\DP/RegALU2/N3 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[0] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[0]  ( .D(\DP/RegA1/N3 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[0] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[0]  ( .D(\PC/N3 ), .CK(n635), .Q(\DP/NPC1[0] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[1]  ( .D(\DP/RegALU1/N4 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[1]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[1]  ( .D(\DP/RegALU2/N4 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[1] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[1]  ( .D(\DP/RegA1/N4 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[1] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[1]  ( .D(\DP/RegNPC1/N4 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[1] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[1]  ( .D(\DP/RegNPC2/N4 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[1] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[2]  ( .D(\DP/RegALU1/N5 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[2]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[2]  ( .D(\DP/RegALU2/N5 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[2] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[2]  ( .D(\DP/RegA1/N5 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[2] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[2]  ( .D(\PC/N5 ), .CK(n635), .Q(\DP/NPC1[2] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[2]  ( .D(\DP/RegNPC1/N5 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[2] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[2]  ( .D(\DP/RegNPC2/N5 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[2] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[3]  ( .D(\DP/RegALU2/N6 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[3] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[3]  ( .D(\DP/RegA1/N6 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[3] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[3]  ( .D(\PC/N6 ), .CK(n635), .Q(\DP/NPC1[3] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[3]  ( .D(\DP/RegNPC1/N6 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[3] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[3]  ( .D(\DP/RegNPC2/N6 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[3] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[4]  ( .D(\DP/RegALU1/N7 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[4]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[4]  ( .D(\DP/RegALU2/N7 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[4] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[4]  ( .D(\DP/RegA1/N7 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[4] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[4]  ( .D(\PC/N7 ), .CK(n635), .Q(\DP/NPC1[4] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[4]  ( .D(\DP/RegNPC1/N7 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[4] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[4]  ( .D(\DP/RegNPC2/N7 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[4] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[5]  ( .D(\DP/RegALU1/N8 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[5]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[5]  ( .D(\DP/RegALU2/N8 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[5] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[5]  ( .D(\DP/RegA1/N8 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[5] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[5]  ( .D(\PC/N8 ), .CK(n635), .Q(\DP/NPC1[5] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[5]  ( .D(\DP/RegNPC2/N8 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[5] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[6]  ( .D(\DP/RegALU1/N9 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[6]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[6]  ( .D(\DP/RegALU2/N9 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[6] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[6]  ( .D(\DP/RegA1/N9 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[6] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[7]  ( .D(\DP/RegALU2/N10 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[7] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[7]  ( .D(\DP/RegA1/N10 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[7] ) );
  DFF_X1 \PC/DOUT_reg[7]  ( .D(\PC/N10 ), .CK(n635), .Q(IROM_ADDR[7]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[7]  ( .D(\PC/N10 ), .CK(\DP/RegNPC/net7068 ), .Q(
        \DP/NPC1[7] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[7]  ( .D(\DP/RegNPC2/N10 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[7] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[8]  ( .D(\DP/RegALU2/N11 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[8] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[8]  ( .D(\DP/RegA1/N11 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[8] ) );
  DFF_X1 \PC/DOUT_reg[8]  ( .D(\PC/N11 ), .CK(n635), .Q(IROM_ADDR[8]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[8]  ( .D(\PC/N11 ), .CK(\DP/RegNPC/net7068 ), .Q(
        \DP/NPC1[8] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[8]  ( .D(\DP/RegNPC2/N11 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[8] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[9]  ( .D(\DP/RegALU2/N12 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[9] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[9]  ( .D(\DP/RegA1/N12 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[9] ) );
  DFF_X1 \PC/DOUT_reg[9]  ( .D(\PC/N12 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IROM_ADDR[9]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[9]  ( .D(\PC/N12 ), .CK(n635), .Q(\DP/NPC1[9] )
         );
  DFF_X1 \DP/RegNPC2/DOUT_reg[9]  ( .D(\DP/RegNPC2/N12 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[9] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[10]  ( .D(\DP/RegALU2/N13 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[10] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[10]  ( .D(\DP/RegA1/N13 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[10] ) );
  DFF_X1 \PC/DOUT_reg[10]  ( .D(\PC/N13 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IROM_ADDR[10]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[10]  ( .D(\PC/N13 ), .CK(n635), .Q(\DP/NPC1[10] )
         );
  DFF_X1 \DP/RegNPC2/DOUT_reg[10]  ( .D(\DP/RegNPC2/N13 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[10] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[11]  ( .D(\DP/RegALU2/N14 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[11] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[11]  ( .D(\DP/RegA1/N14 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[11] ) );
  DFF_X1 \PC/DOUT_reg[11]  ( .D(\PC/N14 ), .CK(n635), .Q(IROM_ADDR[11]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[11]  ( .D(\PC/N14 ), .CK(\DP/RegNPC/net7068 ), 
        .Q(\DP/NPC1[11] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[11]  ( .D(\DP/RegNPC2/N14 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[11] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[12]  ( .D(\DP/RegALU2/N15 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[12] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[12]  ( .D(\DP/RegA1/N15 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[12] ) );
  DFF_X1 \PC/DOUT_reg[12]  ( .D(\PC/N15 ), .CK(\DP/RegNPC/net7068 ), .Q(
        w_PC_OUT[12]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[12]  ( .D(\PC/N15 ), .CK(n635), .Q(\DP/NPC1[12] )
         );
  DFF_X1 \DP/RegNPC2/DOUT_reg[12]  ( .D(\DP/RegNPC2/N15 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[12] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[13]  ( .D(\DP/RegALU2/N16 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[13] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[13]  ( .D(\DP/RegA1/N16 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[13] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[13]  ( .D(\PC/N16 ), .CK(n635), .Q(\DP/NPC1[13] )
         );
  DFF_X1 \DP/RegNPC1/DOUT_reg[13]  ( .D(\DP/RegNPC1/N16 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[13] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[13]  ( .D(\DP/RegNPC2/N16 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[13] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[14]  ( .D(\DP/RegALU2/N17 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[14] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[14]  ( .D(\DP/RegA1/N17 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[14] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[14]  ( .D(\PC/N17 ), .CK(n635), .Q(\DP/NPC1[14] )
         );
  DFF_X1 \DP/RegNPC1/DOUT_reg[14]  ( .D(\DP/RegNPC1/N17 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[14] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[14]  ( .D(\DP/RegNPC2/N17 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[14] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[15]  ( .D(\DP/RegALU2/N18 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[15] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[15]  ( .D(\DP/RegA1/N18 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[15] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[15]  ( .D(\PC/N18 ), .CK(\DP/RegNPC/net7068 ), 
        .Q(\DP/NPC1[15] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[15]  ( .D(\DP/RegNPC1/N18 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[15] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[15]  ( .D(\DP/RegNPC2/N18 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[15] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[16]  ( .D(\DP/RegALU2/N19 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[16] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[16]  ( .D(\DP/RegA1/N19 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[16] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[16]  ( .D(\PC/N19 ), .CK(n635), .Q(\DP/NPC1[16] )
         );
  DFF_X1 \DP/RegNPC1/DOUT_reg[16]  ( .D(\DP/RegNPC1/N19 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[16] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[16]  ( .D(\DP/RegNPC2/N19 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[16] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[17]  ( .D(\DP/RegALU2/N20 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[17] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[17]  ( .D(\DP/RegA1/N20 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[17] ) );
  DFF_X1 \PC/DOUT_reg[17]  ( .D(n1460), .CK(\DP/RegNPC/net7068 ), .Q(
        w_PC_OUT[17]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[17]  ( .D(\PC/N20 ), .CK(n635), .Q(\DP/NPC1[17] )
         );
  DFF_X1 \DP/RegNPC2/DOUT_reg[17]  ( .D(\DP/RegNPC2/N20 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[17] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[18]  ( .D(\DP/RegALU2/N21 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[18] ) );
  DFF_X1 \PC/DOUT_reg[18]  ( .D(\PC/N21 ), .CK(n635), .Q(w_PC_OUT[18]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[18]  ( .D(\PC/N21 ), .CK(\DP/RegNPC/net7068 ), 
        .Q(\DP/NPC1[18] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[18]  ( .D(\DP/RegNPC2/N21 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[18] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[19]  ( .D(\DP/RegALU2/N22 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[19] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[19]  ( .D(\DP/RegA1/N22 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[19] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[19]  ( .D(\PC/N22 ), .CK(n635), .Q(\DP/NPC1[19] )
         );
  DFF_X1 \DP/RegNPC1/DOUT_reg[19]  ( .D(\DP/RegNPC1/N22 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[19] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[19]  ( .D(\DP/RegNPC2/N22 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[19] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[20]  ( .D(\DP/RegALU2/N23 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[20] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[20]  ( .D(\DP/RegA1/N23 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[20] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[20]  ( .D(\DP/RegNPC1/N23 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[20] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[20]  ( .D(\DP/RegNPC2/N23 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[20] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[21]  ( .D(\DP/RegALU2/N24 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[21] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[21]  ( .D(\DP/RegA1/N24 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[21] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[21]  ( .D(\DP/RegNPC2/N24 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[21] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[22]  ( .D(\DP/RegALU2/N25 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[22] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[22]  ( .D(\DP/RegA1/N25 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[22] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[22]  ( .D(\PC/N25 ), .CK(n635), .Q(\DP/NPC1[22] )
         );
  DFF_X1 \DP/RegNPC1/DOUT_reg[22]  ( .D(\DP/RegNPC1/N25 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[22] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[22]  ( .D(\DP/RegNPC2/N25 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[22] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[23]  ( .D(\DP/RegALU2/N26 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[23] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[23]  ( .D(\DP/RegA1/N26 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[23] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[23]  ( .D(\PC/N26 ), .CK(n635), .Q(\DP/NPC1[23] )
         );
  DFF_X1 \DP/RegNPC1/DOUT_reg[23]  ( .D(\DP/RegNPC1/N26 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[23] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[23]  ( .D(\DP/RegNPC2/N26 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[23] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[24]  ( .D(\DP/RegALU2/N27 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[24] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[24]  ( .D(\DP/RegA1/N27 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[24] ) );
  DFF_X1 \PC/DOUT_reg[24]  ( .D(\PC/N27 ), .CK(n635), .Q(w_PC_OUT[24]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[24]  ( .D(\PC/N27 ), .CK(\DP/RegNPC/net7068 ), 
        .Q(\DP/NPC1[24] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[24]  ( .D(\DP/RegNPC2/N27 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[24] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[25]  ( .D(\DP/RegALU2/N28 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[25] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[25]  ( .D(\DP/RegA1/N28 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[25] ) );
  DFF_X1 \PC/DOUT_reg[25]  ( .D(\PC/N28 ), .CK(\DP/RegNPC/net7068 ), .Q(
        w_PC_OUT[25]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[25]  ( .D(\PC/N28 ), .CK(n635), .Q(\DP/NPC1[25] )
         );
  DFF_X1 \DP/RegNPC2/DOUT_reg[25]  ( .D(\DP/RegNPC2/N28 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[25] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[26]  ( .D(\DP/RegALU2/N29 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[26] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[26]  ( .D(\DP/RegA1/N29 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[26] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[26]  ( .D(\DP/RegNPC2/N29 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[26] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[27]  ( .D(\DP/RegALU2/N30 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[27] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[27]  ( .D(\DP/RegA1/N30 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[27] ) );
  DFF_X1 \PC/DOUT_reg[27]  ( .D(\PC/N30 ), .CK(n635), .Q(w_PC_OUT[27]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[27]  ( .D(\PC/N30 ), .CK(\DP/RegNPC/net7068 ), 
        .Q(\DP/NPC1[27] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[27]  ( .D(\DP/RegNPC2/N30 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[27] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[28]  ( .D(\DP/RegALU2/N31 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[28] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[28]  ( .D(\DP/RegA1/N31 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[28] ) );
  DFF_X1 \PC/DOUT_reg[28]  ( .D(\PC/N31 ), .CK(\DP/RegNPC/net7068 ), .Q(
        w_PC_OUT[28]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[28]  ( .D(\PC/N31 ), .CK(n635), .Q(\DP/NPC1[28] )
         );
  DFF_X1 \DP/RegNPC2/DOUT_reg[28]  ( .D(\DP/RegNPC2/N31 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[28] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[29]  ( .D(\DP/RegALU2/N32 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[29] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[29]  ( .D(\DP/RegA1/N32 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[29] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[29]  ( .D(\PC/N32 ), .CK(\DP/RegNPC/net7068 ), 
        .Q(\DP/NPC1[29] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[29]  ( .D(\DP/RegNPC1/N32 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[29] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[29]  ( .D(\DP/RegNPC2/N32 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[29] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[30]  ( .D(\DP/RegALU1/N33 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[30] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[30]  ( .D(\DP/RegALU2/N33 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[30] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[30]  ( .D(\DP/RegA1/N33 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/RegA1_out[30] ) );
  DFF_X1 \PC/DOUT_reg[30]  ( .D(\PC/N33 ), .CK(n635), .Q(w_PC_OUT[30]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[30]  ( .D(\PC/N33 ), .CK(\DP/RegNPC/net7068 ), 
        .Q(\DP/NPC1[30] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[30]  ( .D(\DP/RegNPC2/N33 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[30] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[31]  ( .D(\DP/RegALU1/N34 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[31] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[31]  ( .D(\DP/RegALU2/N34 ), .CK(
        \DP/RegALU2/net7068 ), .Q(\DP/RegALU2_out[31] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[31]  ( .D(\DP/RegNPC2/N34 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[31] ) );
  AND2_X1 U1179 ( .A1(RST), .A2(\DP/RES[31] ), .ZN(\DP/RegALU1/N34 ) );
  AND2_X1 U1180 ( .A1(RST), .A2(\DP/RES[19] ), .ZN(\DP/RegALU1/N22 ) );
  AND2_X1 U1181 ( .A1(RST), .A2(\DP/RES[17] ), .ZN(\DP/RegALU1/N20 ) );
  AND2_X1 U1182 ( .A1(\DP/RES[0] ), .A2(RST), .ZN(\DP/RegALU1/N3 ) );
  AND2_X1 U1183 ( .A1(RST), .A2(\DP/RES[8] ), .ZN(\DP/RegALU1/N11 ) );
  AND2_X1 U1184 ( .A1(n1043), .A2(n1317), .ZN(n580) );
  NOR2_X1 U1185 ( .A1(n744), .A2(n745), .ZN(n581) );
  NOR2_X1 U1186 ( .A1(n747), .A2(n581), .ZN(n582) );
  OAI222_X1 U1187 ( .A1(n640), .A2(n580), .B1(n759), .B2(n582), .C1(n749), 
        .C2(n748), .ZN(\CU/N88 ) );
  NOR2_X2 U1188 ( .A1(n640), .A2(n682), .ZN(n1056) );
  NOR2_X2 U1189 ( .A1(\DP/FwdD ), .A2(n1223), .ZN(n1257) );
  OAI21_X2 U1190 ( .B1(n1225), .B2(n1224), .A(n1267), .ZN(n1256) );
  NAND2_X1 U1192 ( .A1(n1071), .A2(n1070), .ZN(n1087) );
  AND2_X1 U1193 ( .A1(RST), .A2(n1068), .ZN(n1088) );
  NAND3_X1 U1194 ( .A1(n1058), .A2(\DP/LOAD8[7] ), .A3(w_SIGN_LD), .ZN(n1071)
         );
  OAI21_X1 U1195 ( .B1(n1069), .B2(n1068), .A(RST), .ZN(n1067) );
  AND2_X1 U1196 ( .A1(RST), .A2(IROM_DATA[1]), .ZN(\IR/N4 ) );
  AND2_X1 U1197 ( .A1(RST), .A2(IROM_DATA[2]), .ZN(\IR/N5 ) );
  AND2_X1 U1198 ( .A1(RST), .A2(IROM_DATA[3]), .ZN(\IR/N6 ) );
  AND2_X1 U1199 ( .A1(RST), .A2(IROM_DATA[4]), .ZN(\IR/N7 ) );
  AND2_X1 U1200 ( .A1(RST), .A2(IROM_DATA[5]), .ZN(\IR/N8 ) );
  AND2_X1 U1201 ( .A1(RST), .A2(IROM_DATA[6]), .ZN(\IR/N9 ) );
  AND2_X1 U1202 ( .A1(RST), .A2(IROM_DATA[7]), .ZN(\IR/N10 ) );
  AND2_X1 U1203 ( .A1(RST), .A2(IROM_DATA[8]), .ZN(\IR/N11 ) );
  AND2_X1 U1204 ( .A1(RST), .A2(IROM_DATA[9]), .ZN(\IR/N12 ) );
  AND2_X1 U1205 ( .A1(RST), .A2(IROM_DATA[10]), .ZN(\IR/N13 ) );
  AND2_X1 U1206 ( .A1(RST), .A2(IROM_DATA[11]), .ZN(\IR/N14 ) );
  AND2_X1 U1207 ( .A1(RST), .A2(IROM_DATA[12]), .ZN(\IR/N15 ) );
  AND2_X1 U1208 ( .A1(RST), .A2(IROM_DATA[13]), .ZN(\IR/N16 ) );
  AND2_X1 U1209 ( .A1(RST), .A2(IROM_DATA[14]), .ZN(\IR/N17 ) );
  AND2_X1 U1210 ( .A1(RST), .A2(IROM_DATA[15]), .ZN(\IR/N18 ) );
  AND2_X1 U1211 ( .A1(RST), .A2(IROM_DATA[16]), .ZN(\IR/N19 ) );
  AND2_X1 U1212 ( .A1(RST), .A2(IROM_DATA[17]), .ZN(\IR/N20 ) );
  AND2_X1 U1213 ( .A1(RST), .A2(IROM_DATA[18]), .ZN(\IR/N21 ) );
  AND2_X1 U1214 ( .A1(RST), .A2(IROM_DATA[19]), .ZN(\IR/N22 ) );
  AND2_X1 U1215 ( .A1(RST), .A2(IROM_DATA[20]), .ZN(\IR/N23 ) );
  AND2_X1 U1216 ( .A1(RST), .A2(IROM_DATA[21]), .ZN(\IR/N24 ) );
  AND2_X1 U1217 ( .A1(RST), .A2(IROM_DATA[22]), .ZN(\IR/N25 ) );
  AND2_X1 U1218 ( .A1(RST), .A2(IROM_DATA[23]), .ZN(\IR/N26 ) );
  AND2_X1 U1219 ( .A1(RST), .A2(IROM_DATA[24]), .ZN(\IR/N27 ) );
  AND2_X1 U1220 ( .A1(RST), .A2(IROM_DATA[25]), .ZN(\IR/N28 ) );
  AND2_X1 U1221 ( .A1(RST), .A2(IROM_DATA[26]), .ZN(\IR/N29 ) );
  AND2_X1 U1222 ( .A1(RST), .A2(IROM_DATA[27]), .ZN(\IR/N30 ) );
  AND2_X1 U1223 ( .A1(RST), .A2(IROM_DATA[28]), .ZN(\IR/N31 ) );
  AND2_X1 U1224 ( .A1(RST), .A2(IROM_DATA[29]), .ZN(\IR/N32 ) );
  AND2_X1 U1225 ( .A1(RST), .A2(IROM_DATA[30]), .ZN(\IR/N33 ) );
  AND2_X1 U1226 ( .A1(RST), .A2(IROM_DATA[31]), .ZN(\IR/N34 ) );
  OR2_X1 U1227 ( .A1(n640), .A2(n1039), .ZN(n1052) );
  AND2_X1 U1228 ( .A1(RST), .A2(n676), .ZN(\CU/N82 ) );
  INV_X1 U1229 ( .A(RST), .ZN(n640) );
  INV_X1 U1230 ( .A(RST), .ZN(n641) );
  OR2_X1 U1235 ( .A1(n641), .A2(n655), .ZN(n657) );
  AND2_X1 U1237 ( .A1(RST), .A2(IROM_DATA[0]), .ZN(\IR/N3 ) );
  AND2_X1 U1238 ( .A1(RST), .A2(\DP/RegALU1_out[14] ), .ZN(\DP/RegALU2/N17 )
         );
  AND2_X1 U1239 ( .A1(RST), .A2(\DP/RegALU1_out[15] ), .ZN(\DP/RegALU2/N18 )
         );
  AND2_X1 U1240 ( .A1(RST), .A2(\DP/RegALU1_out[16] ), .ZN(\DP/RegALU2/N19 )
         );
  AND2_X1 U1241 ( .A1(RST), .A2(\DP/RegALU1_out[17] ), .ZN(\DP/RegALU2/N20 )
         );
  AND2_X1 U1242 ( .A1(RST), .A2(\DP/RegALU1_out[18] ), .ZN(\DP/RegALU2/N21 )
         );
  AND2_X1 U1243 ( .A1(RST), .A2(\DP/RegALU1_out[19] ), .ZN(\DP/RegALU2/N22 )
         );
  AND2_X1 U1244 ( .A1(RST), .A2(\DP/RegALU1_out[20] ), .ZN(\DP/RegALU2/N23 )
         );
  AND2_X1 U1245 ( .A1(RST), .A2(\DP/RegALU1_out[21] ), .ZN(\DP/RegALU2/N24 )
         );
  AND2_X1 U1246 ( .A1(RST), .A2(\DP/RegALU1_out[29] ), .ZN(\DP/RegALU2/N32 )
         );
  AND2_X1 U1247 ( .A1(RST), .A2(\DP/RegALU1_out[28] ), .ZN(\DP/RegALU2/N31 )
         );
  AND2_X1 U1248 ( .A1(RST), .A2(\DP/RegALU1_out[27] ), .ZN(\DP/RegALU2/N30 )
         );
  AND2_X1 U1249 ( .A1(RST), .A2(\DP/RegALU1_out[30] ), .ZN(\DP/RegALU2/N33 )
         );
  AND2_X1 U1250 ( .A1(RST), .A2(\DP/RegALU1_out[26] ), .ZN(\DP/RegALU2/N29 )
         );
  AND2_X1 U1251 ( .A1(RST), .A2(\DP/RegALU1_out[25] ), .ZN(\DP/RegALU2/N28 )
         );
  AND2_X1 U1252 ( .A1(RST), .A2(\DP/RegALU1_out[24] ), .ZN(\DP/RegALU2/N27 )
         );
  AND2_X1 U1253 ( .A1(RST), .A2(\DP/RegALU1_out[23] ), .ZN(\DP/RegALU2/N26 )
         );
  AND2_X1 U1254 ( .A1(RST), .A2(\DP/RegALU1_out[22] ), .ZN(\DP/RegALU2/N25 )
         );
  AND2_X1 U1255 ( .A1(RST), .A2(\DP/RegALU1_out[31] ), .ZN(\DP/RegALU2/N34 )
         );
  AND2_X1 U1264 ( .A1(RST), .A2(DRAM_ADDR[0]), .ZN(\DP/RegALU2/N3 ) );
  AND2_X1 U1265 ( .A1(RST), .A2(DRAM_ADDR[1]), .ZN(\DP/RegALU2/N4 ) );
  AND2_X1 U1266 ( .A1(RST), .A2(DRAM_ADDR[2]), .ZN(\DP/RegALU2/N5 ) );
  AND2_X1 U1267 ( .A1(RST), .A2(DRAM_ADDR[3]), .ZN(\DP/RegALU2/N6 ) );
  AND2_X1 U1268 ( .A1(RST), .A2(DRAM_ADDR[4]), .ZN(\DP/RegALU2/N7 ) );
  AND2_X1 U1270 ( .A1(RST), .A2(\DP/RegALU1_out[13] ), .ZN(\DP/RegALU2/N16 )
         );
  AND2_X1 U1271 ( .A1(RST), .A2(\DP/RegALU1_out[12] ), .ZN(\DP/RegALU2/N15 )
         );
  BUF_X1 U1272 ( .A(n892), .Z(n622) );
  BUF_X1 U1273 ( .A(n893), .Z(n623) );
  AND2_X1 U1275 ( .A1(RST), .A2(DRAM_ADDR[11]), .ZN(\DP/RegALU2/N14 ) );
  BUF_X1 U1276 ( .A(n894), .Z(n625) );
  NOR2_X1 U1277 ( .A1(n835), .A2(n609), .ZN(n894) );
  NOR2_X1 U1278 ( .A1(w_MuxB_SEL), .A2(n835), .ZN(n892) );
  BUF_X1 U1279 ( .A(n893), .Z(n624) );
  NOR3_X1 U1280 ( .A1(n75), .A2(\DP/FwdB[1] ), .A3(\DP/FwdB[0] ), .ZN(n893) );
  BUF_X1 U1281 ( .A(n897), .Z(n626) );
  NAND3_X1 U1282 ( .A1(\DP/FwdB[1] ), .A2(n75), .A3(n605), .ZN(n897) );
  AND2_X1 U1284 ( .A1(RST), .A2(DRAM_ADDR[10]), .ZN(\DP/RegALU2/N13 ) );
  AND2_X1 U1286 ( .A1(RST), .A2(DRAM_ADDR[9]), .ZN(\DP/RegALU2/N12 ) );
  AND2_X1 U1287 ( .A1(RST), .A2(DRAM_ADDR[8]), .ZN(\DP/RegALU2/N11 ) );
  INV_X1 U1288 ( .A(n591), .ZN(n633) );
  AND2_X1 U1290 ( .A1(RST), .A2(DRAM_ADDR[7]), .ZN(\DP/RegALU2/N10 ) );
  BUF_X1 U1291 ( .A(n1009), .Z(n629) );
  AND2_X1 U1292 ( .A1(RST), .A2(DRAM_ADDR[6]), .ZN(\DP/RegALU2/N9 ) );
  BUF_X1 U1293 ( .A(n829), .Z(n618) );
  BUF_X1 U1294 ( .A(n1195), .Z(n631) );
  AND3_X1 U1295 ( .A1(RST), .A2(\DP/OUTCOME ), .A3(\DP/JREG ), .ZN(n1195) );
  BUF_X1 U1296 ( .A(n1196), .Z(n632) );
  NOR2_X1 U1297 ( .A1(\DP/JREG ), .A2(n607), .ZN(n1196) );
  INV_X1 U1298 ( .A(n591), .ZN(n634) );
  OR2_X1 U1299 ( .A1(n640), .A2(\DP/OUTCOME ), .ZN(n591) );
  BUF_X1 U1302 ( .A(n831), .Z(n620) );
  NOR2_X1 U1303 ( .A1(w_MuxA_SEL), .A2(n765), .ZN(n831) );
  BUF_X1 U1304 ( .A(n830), .Z(n619) );
  NOR2_X1 U1305 ( .A1(n608), .A2(n765), .ZN(n830) );
  AND3_X1 U1306 ( .A1(n76), .A2(\DP/FwdA[2] ), .A3(n69), .ZN(n829) );
  BUF_X1 U1307 ( .A(n834), .Z(n621) );
  INV_X1 U1308 ( .A(n824), .ZN(n834) );
  NOR3_X1 U1309 ( .A1(\DP/FwdA[2] ), .A2(n69), .A3(n588), .ZN(n824) );
  AND2_X1 U1310 ( .A1(RST), .A2(DRAM_ADDR[5]), .ZN(\DP/RegALU2/N8 ) );
  AND2_X1 U1312 ( .A1(RST), .A2(n975), .ZN(n1009) );
  BUF_X1 U1313 ( .A(n1011), .Z(n630) );
  OR2_X1 U1314 ( .A1(n641), .A2(n974), .ZN(n1011) );
  OAI21_X1 U1318 ( .B1(\DP/JL2 ), .B2(n1237), .A(n954), .ZN(\DP/RF_DATA[21] )
         );
  OAI21_X1 U1320 ( .B1(n1492), .B2(n1247), .A(n959), .ZN(\DP/RF_DATA[26] ) );
  OAI21_X1 U1321 ( .B1(\DP/JL2 ), .B2(n1231), .A(n950), .ZN(\DP/RF_DATA[18] )
         );
  OAI21_X1 U1322 ( .B1(\DP/JL2 ), .B2(n1243), .A(n957), .ZN(\DP/RF_DATA[24] )
         );
  OAI21_X1 U1323 ( .B1(n1492), .B2(n1239), .A(n955), .ZN(\DP/RF_DATA[22] ) );
  INV_X1 U1326 ( .A(n1203), .ZN(n36) );
  INV_X1 U1328 ( .A(n1204), .ZN(n34) );
  INV_X1 U1329 ( .A(n1206), .ZN(n37) );
  INV_X1 U1334 ( .A(n1047), .ZN(n38) );
  INV_X1 U1336 ( .A(n1049), .ZN(n41) );
  OR2_X1 U1337 ( .A1(n1488), .A2(\DP/RD3[3] ), .ZN(\DP/RF_ADDR[3] ) );
  INV_X1 U1338 ( .A(n1051), .ZN(n42) );
  INV_X1 U1340 ( .A(n1280), .ZN(n40) );
  OR2_X1 U1341 ( .A1(n1488), .A2(\DP/RD3[2] ), .ZN(\DP/RF_ADDR[2] ) );
  INV_X1 U1342 ( .A(n1822), .ZN(n39) );
  OR2_X1 U1343 ( .A1(\DP/JL2 ), .A2(\DP/RD3[1] ), .ZN(\DP/RF_ADDR[1] ) );
  BUF_X1 U1345 ( .A(\DP/RegNPC/net7068 ), .Z(n635) );
  OR2_X1 U1348 ( .A1(n589), .A2(n1223), .ZN(n1259) );
  OR2_X1 U1360 ( .A1(n656), .A2(n662), .ZN(n12) );
  INV_X1 U1362 ( .A(n1495), .ZN(n682) );
  NOR2_X1 U1388 ( .A1(n1484), .A2(n62), .ZN(n652) );
  NAND2_X1 U1395 ( .A1(n1327), .A2(n1451), .ZN(n713) );
  NOR2_X1 U1396 ( .A1(n1333), .A2(n713), .ZN(n752) );
  NAND2_X1 U1398 ( .A1(n1041), .A2(n666), .ZN(n702) );
  NAND2_X1 U1405 ( .A1(n1419), .A2(n1432), .ZN(n694) );
  NAND3_X1 U1406 ( .A1(n1041), .A2(n1451), .A3(n1375), .ZN(n653) );
  AOI21_X1 U1408 ( .B1(n694), .B2(n710), .A(n739), .ZN(n1043) );
  INV_X1 U1411 ( .A(n1830), .ZN(n1201) );
  AOI21_X1 U1412 ( .B1(n1202), .B2(n1201), .A(n640), .ZN(\CU/N55 ) );
  INV_X1 U1413 ( .A(\CU/N55 ), .ZN(n654) );
  NAND2_X1 U1414 ( .A1(n654), .A2(n12), .ZN(\CU/N42 ) );
  NOR2_X1 U1415 ( .A1(n640), .A2(n1354), .ZN(\CU/N45 ) );
  NOR2_X1 U1416 ( .A1(n656), .A2(n657), .ZN(\CU/N46 ) );
  NOR2_X1 U1417 ( .A1(n1549), .A2(n657), .ZN(\CU/N47 ) );
  NOR2_X1 U1418 ( .A1(n661), .A2(n657), .ZN(\CU/N48 ) );
  NOR3_X1 U1419 ( .A1(n1299), .A2(n1578), .A3(n657), .ZN(\CU/N49 ) );
  NAND3_X1 U1420 ( .A1(n1464), .A2(n1712), .A3(RST), .ZN(n659) );
  NOR2_X1 U1421 ( .A1(n690), .A2(n659), .ZN(\CU/N50 ) );
  NOR2_X1 U1422 ( .A1(n1549), .A2(n659), .ZN(\CU/N51 ) );
  NOR2_X1 U1423 ( .A1(n661), .A2(n659), .ZN(\CU/N52 ) );
  NOR2_X1 U1425 ( .A1(n640), .A2(n1368), .ZN(\CU/N56 ) );
  AOI21_X1 U1426 ( .B1(n1201), .B2(n1368), .A(n640), .ZN(\CU/N54 ) );
  AND2_X1 U1428 ( .A1(RST), .A2(n1352), .ZN(\CU/N58 ) );
  NOR3_X1 U1430 ( .A1(n663), .A2(n1547), .A3(n662), .ZN(\CU/N60 ) );
  NAND3_X1 U1433 ( .A1(n1201), .A2(n1039), .A3(n1368), .ZN(n668) );
  NOR2_X1 U1435 ( .A1(n641), .A2(n1297), .ZN(\CU/N61 ) );
  NOR2_X1 U1440 ( .A1(n972), .A2(n640), .ZN(\CU/N62 ) );
  NOR2_X1 U1444 ( .A1(n1296), .A2(n641), .ZN(\CU/N63 ) );
  AND2_X1 U1445 ( .A1(RST), .A2(w_RF_WE_EX), .ZN(\CU/N64 ) );
  AND2_X1 U1446 ( .A1(RST), .A2(\CU/cw1[1] ), .ZN(\CU/N65 ) );
  AND2_X1 U1447 ( .A1(RST), .A2(\CU/cw1[2] ), .ZN(\CU/N66 ) );
  AND2_X1 U1448 ( .A1(RST), .A2(\CU/cw1[3] ), .ZN(\CU/N67 ) );
  AND2_X1 U1449 ( .A1(RST), .A2(\CU/cw1[4] ), .ZN(\CU/N68 ) );
  AND2_X1 U1450 ( .A1(RST), .A2(\CU/cw1[5] ), .ZN(\CU/N69 ) );
  AND2_X1 U1451 ( .A1(RST), .A2(\CU/cw1[6] ), .ZN(\CU/N70 ) );
  AND2_X1 U1452 ( .A1(RST), .A2(\CU/cw1[7] ), .ZN(\CU/N71 ) );
  AND2_X1 U1453 ( .A1(RST), .A2(\CU/cw1[8] ), .ZN(\CU/N72 ) );
  AND2_X1 U1454 ( .A1(RST), .A2(\CU/cw1[9] ), .ZN(\CU/N73 ) );
  AND2_X1 U1455 ( .A1(RST), .A2(\CU/cw1[10] ), .ZN(\CU/N74 ) );
  AND2_X1 U1456 ( .A1(RST), .A2(\CU/cw1[11] ), .ZN(\CU/N75 ) );
  AND2_X1 U1457 ( .A1(RST), .A2(\CU/cw1[12] ), .ZN(\CU/N76 ) );
  AND2_X1 U1458 ( .A1(RST), .A2(\CU/cw1[13] ), .ZN(\CU/N77 ) );
  AND2_X1 U1459 ( .A1(RST), .A2(\CU/cw1[14] ), .ZN(\CU/N78 ) );
  NOR2_X1 U1460 ( .A1(n641), .A2(n601), .ZN(\CU/N79 ) );
  AND2_X1 U1461 ( .A1(RST), .A2(\CU/cw2[1] ), .ZN(\CU/N80 ) );
  AND2_X1 U1462 ( .A1(RST), .A2(\CU/cw2[2] ), .ZN(\CU/N81 ) );
  INV_X1 U1465 ( .A(n1472), .ZN(n683) );
  NAND3_X1 U1466 ( .A1(n1544), .A2(IR_OUT[5]), .A3(n595), .ZN(n715) );
  NOR3_X1 U1467 ( .A1(n683), .A2(n1053), .A3(n1314), .ZN(n737) );
  NOR2_X1 U1468 ( .A1(n1472), .A2(n1313), .ZN(n717) );
  NAND2_X1 U1469 ( .A1(n717), .A2(n1053), .ZN(n757) );
  NOR2_X1 U1470 ( .A1(n1472), .A2(n1053), .ZN(n731) );
  NAND2_X1 U1472 ( .A1(n736), .A2(n1658), .ZN(n724) );
  INV_X1 U1473 ( .A(n724), .ZN(n735) );
  NAND3_X1 U1474 ( .A1(n1311), .A2(n735), .A3(n1446), .ZN(n677) );
  OR2_X1 U1476 ( .A1(n1313), .A2(n718), .ZN(n744) );
  INV_X1 U1477 ( .A(n1329), .ZN(n679) );
  NOR3_X1 U1478 ( .A1(n1053), .A2(n679), .A3(n683), .ZN(n722) );
  INV_X1 U1479 ( .A(n722), .ZN(n749) );
  OAI22_X1 U1480 ( .A1(n716), .A2(n744), .B1(n724), .B2(n749), .ZN(n680) );
  AOI211_X1 U1481 ( .C1(n1312), .C2(n736), .A(n747), .B(n680), .ZN(n701) );
  NAND2_X1 U1483 ( .A1(RST), .A2(n755), .ZN(n759) );
  AND2_X1 U1484 ( .A1(IR_OUT[5]), .A2(n1056), .ZN(\DP/RegIMM/N8 ) );
  AND4_X1 U1485 ( .A1(n1053), .A2(n683), .A3(IR_OUT[4]), .A4(n755), .ZN(n684)
         );
  NAND2_X1 U1486 ( .A1(\DP/RegIMM/N8 ), .A2(n684), .ZN(n723) );
  NAND3_X1 U1488 ( .A1(n694), .A2(n1538), .A3(RST), .ZN(n728) );
  INV_X1 U1489 ( .A(n728), .ZN(n686) );
  NOR4_X1 U1490 ( .A1(n760), .A2(n686), .A3(\CU/N82 ), .A4(\CU/N54 ), .ZN(n700) );
  AOI21_X1 U1491 ( .B1(n1482), .B2(n1457), .A(n1843), .ZN(n692) );
  NOR2_X1 U1493 ( .A1(n693), .A2(n1470), .ZN(n695) );
  OAI21_X1 U1495 ( .B1(n1299), .B2(n702), .A(n696), .ZN(n698) );
  OAI21_X1 U1496 ( .B1(n706), .B2(n698), .A(RST), .ZN(n699) );
  OAI211_X1 U1497 ( .C1(n701), .C2(n759), .A(n699), .B(n700), .ZN(\CU/N85 ) );
  INV_X1 U1498 ( .A(n736), .ZN(n730) );
  NAND3_X1 U1500 ( .A1(n730), .A2(n755), .A3(\DP/RegIMM/N4 ), .ZN(n748) );
  NOR3_X1 U1502 ( .A1(n704), .A2(n1549), .A3(n1463), .ZN(n707) );
  NAND3_X1 U1504 ( .A1(n1823), .A2(n62), .A3(n1543), .ZN(n711) );
  OAI211_X1 U1505 ( .C1(n1545), .C2(n1380), .A(n712), .B(n711), .ZN(n727) );
  NAND3_X1 U1507 ( .A1(IR_OUT[4]), .A2(IR_OUT[5]), .A3(n731), .ZN(n758) );
  NOR2_X1 U1508 ( .A1(n717), .A2(n737), .ZN(n719) );
  AOI21_X1 U1514 ( .B1(n757), .B2(n749), .A(n730), .ZN(n734) );
  INV_X1 U1515 ( .A(n731), .ZN(n745) );
  OAI22_X1 U1516 ( .A1(n732), .A2(n758), .B1(n745), .B2(n744), .ZN(n733) );
  NOR2_X1 U1518 ( .A1(n641), .A2(n736), .ZN(\DP/RegIMM/N3 ) );
  INV_X1 U1520 ( .A(n738), .ZN(n740) );
  OAI21_X1 U1521 ( .B1(n740), .B2(n739), .A(RST), .ZN(n741) );
  OAI211_X1 U1522 ( .C1(n743), .C2(n759), .A(n742), .B(n741), .ZN(\CU/N87 ) );
  INV_X1 U1523 ( .A(n1432), .ZN(n753) );
  AOI211_X1 U1524 ( .C1(n754), .C2(n753), .A(n1548), .B(n751), .ZN(n764) );
  NAND2_X1 U1525 ( .A1(n755), .A2(\DP/RegIMM/N3 ), .ZN(n756) );
  OAI22_X1 U1526 ( .A1(n759), .A2(n758), .B1(n757), .B2(n756), .ZN(n761) );
  OAI21_X1 U1528 ( .B1(n764), .B2(n641), .A(n763), .ZN(\CU/N89 ) );
  MUX2_X1 U1529 ( .A(\DP/RegLMD_out[0] ), .B(\DP/RegALU2_out[0] ), .S(n583), 
        .Z(n942) );
  AOI22_X1 U1530 ( .A1(n829), .A2(DRAM_ADDR[0]), .B1(n824), .B2(n942), .ZN(
        n767) );
  NAND3_X1 U1531 ( .A1(n588), .A2(n77), .A3(n69), .ZN(n765) );
  AOI22_X1 U1532 ( .A1(\DP/RegA_out[0] ), .A2(n619), .B1(\DP/NPC2[0] ), .B2(
        n831), .ZN(n766) );
  NAND2_X1 U1533 ( .A1(n767), .A2(n766), .ZN(\DP/A[0] ) );
  AOI22_X1 U1535 ( .A1(\DP/RegA_out[10] ), .A2(n830), .B1(DRAM_ADDR[10]), .B2(
        n618), .ZN(n769) );
  NAND2_X1 U1536 ( .A1(n620), .A2(\DP/NPC2[10] ), .ZN(n768) );
  OAI211_X1 U1537 ( .C1(n1501), .C2(n834), .A(n769), .B(n768), .ZN(\DP/A[10] )
         );
  AOI22_X1 U1538 ( .A1(n1494), .A2(\DP/RegLMD_out[11] ), .B1(
        \DP/RegALU2_out[11] ), .B2(n583), .ZN(n1214) );
  AOI22_X1 U1539 ( .A1(\DP/RegA_out[11] ), .A2(n619), .B1(DRAM_ADDR[11]), .B2(
        n618), .ZN(n771) );
  NAND2_X1 U1540 ( .A1(n620), .A2(\DP/NPC2[11] ), .ZN(n770) );
  OAI211_X1 U1541 ( .C1(n1214), .C2(n621), .A(n771), .B(n770), .ZN(\DP/A[11] )
         );
  AOI22_X1 U1542 ( .A1(n639), .A2(\DP/RegLMD_out[12] ), .B1(
        \DP/RegALU2_out[12] ), .B2(n583), .ZN(n1216) );
  AOI22_X1 U1543 ( .A1(\DP/RegA_out[12] ), .A2(n830), .B1(\DP/RegALU1_out[12] ), .B2(n829), .ZN(n773) );
  NAND2_X1 U1544 ( .A1(n620), .A2(\DP/NPC2[12] ), .ZN(n772) );
  OAI211_X1 U1545 ( .C1(n1216), .C2(n834), .A(n773), .B(n772), .ZN(\DP/A[12] )
         );
  AOI22_X1 U1546 ( .A1(n1494), .A2(\DP/RegLMD_out[13] ), .B1(
        \DP/RegALU2_out[13] ), .B2(n583), .ZN(n1218) );
  AOI22_X1 U1547 ( .A1(\DP/RegALU1_out[13] ), .A2(n829), .B1(\DP/RegA_out[13] ), .B2(n619), .ZN(n775) );
  NAND2_X1 U1548 ( .A1(n620), .A2(\DP/NPC2[13] ), .ZN(n774) );
  OAI211_X1 U1549 ( .C1(n1218), .C2(n621), .A(n775), .B(n774), .ZN(\DP/A[13] )
         );
  AOI22_X1 U1551 ( .A1(\DP/RegALU1_out[14] ), .A2(n829), .B1(\DP/RegA_out[14] ), .B2(n619), .ZN(n777) );
  NAND2_X1 U1552 ( .A1(n620), .A2(\DP/NPC2[14] ), .ZN(n776) );
  OAI211_X1 U1553 ( .C1(n1462), .C2(n834), .A(n777), .B(n776), .ZN(\DP/A[14] )
         );
  AOI22_X1 U1554 ( .A1(\DP/RegALU1_out[15] ), .A2(n829), .B1(\DP/RegA_out[15] ), .B2(n619), .ZN(n779) );
  AOI22_X1 U1555 ( .A1(n1494), .A2(\DP/RegLMD_out[15] ), .B1(
        \DP/RegALU2_out[15] ), .B2(n583), .ZN(n985) );
  INV_X1 U1556 ( .A(n985), .ZN(n1221) );
  AOI22_X1 U1557 ( .A1(\DP/NPC2[15] ), .A2(n831), .B1(n824), .B2(n1221), .ZN(
        n778) );
  NAND2_X1 U1558 ( .A1(n779), .A2(n778), .ZN(\DP/A[15] ) );
  AOI22_X1 U1559 ( .A1(n1494), .A2(\DP/RegLMD_out[16] ), .B1(
        \DP/RegALU2_out[16] ), .B2(n583), .ZN(n1227) );
  AOI22_X1 U1560 ( .A1(\DP/RegALU1_out[16] ), .A2(n618), .B1(\DP/RegA_out[16] ), .B2(n619), .ZN(n781) );
  NAND2_X1 U1561 ( .A1(n620), .A2(\DP/NPC2[16] ), .ZN(n780) );
  OAI211_X1 U1562 ( .C1(n1227), .C2(n621), .A(n781), .B(n780), .ZN(\DP/A[16] )
         );
  AOI22_X1 U1563 ( .A1(n1494), .A2(\DP/RegLMD_out[17] ), .B1(
        \DP/RegALU2_out[17] ), .B2(n638), .ZN(n1229) );
  AOI22_X1 U1564 ( .A1(\DP/RegALU1_out[17] ), .A2(n618), .B1(\DP/RegA_out[17] ), .B2(n619), .ZN(n783) );
  NAND2_X1 U1565 ( .A1(n620), .A2(\DP/NPC2[17] ), .ZN(n782) );
  OAI211_X1 U1566 ( .C1(n1361), .C2(n834), .A(n783), .B(n782), .ZN(\DP/A[17] )
         );
  AOI22_X1 U1567 ( .A1(n639), .A2(\DP/RegLMD_out[18] ), .B1(
        \DP/RegALU2_out[18] ), .B2(n638), .ZN(n1231) );
  AOI22_X1 U1568 ( .A1(\DP/RegALU1_out[18] ), .A2(n829), .B1(\DP/RegA_out[18] ), .B2(n619), .ZN(n785) );
  NAND2_X1 U1569 ( .A1(n620), .A2(\DP/NPC2[18] ), .ZN(n784) );
  OAI211_X1 U1570 ( .C1(n1336), .C2(n621), .A(n785), .B(n784), .ZN(\DP/A[18] )
         );
  AOI22_X1 U1571 ( .A1(n1494), .A2(\DP/RegLMD_out[19] ), .B1(
        \DP/RegALU2_out[19] ), .B2(n638), .ZN(n1233) );
  AOI22_X1 U1572 ( .A1(\DP/RegALU1_out[19] ), .A2(n618), .B1(\DP/RegA_out[19] ), .B2(n619), .ZN(n787) );
  NAND2_X1 U1573 ( .A1(n620), .A2(\DP/NPC2[19] ), .ZN(n786) );
  OAI211_X1 U1574 ( .C1(n1233), .C2(n834), .A(n787), .B(n786), .ZN(\DP/A[19] )
         );
  AOI22_X1 U1575 ( .A1(n1364), .A2(\DP/RegLMD_out[1] ), .B1(
        \DP/RegALU2_out[1] ), .B2(n638), .ZN(n1272) );
  AOI22_X1 U1576 ( .A1(\DP/RegA_out[1] ), .A2(n830), .B1(DRAM_ADDR[1]), .B2(
        n829), .ZN(n789) );
  NAND2_X1 U1577 ( .A1(n831), .A2(\DP/NPC2[1] ), .ZN(n788) );
  OAI211_X1 U1578 ( .C1(n1272), .C2(n834), .A(n789), .B(n788), .ZN(\DP/A[1] )
         );
  AOI22_X1 U1579 ( .A1(n639), .A2(\DP/RegLMD_out[20] ), .B1(
        \DP/RegALU2_out[20] ), .B2(n638), .ZN(n1235) );
  AOI22_X1 U1580 ( .A1(\DP/RegALU1_out[20] ), .A2(n829), .B1(\DP/RegA_out[20] ), .B2(n619), .ZN(n791) );
  NAND2_X1 U1581 ( .A1(n831), .A2(\DP/NPC2[20] ), .ZN(n790) );
  OAI211_X1 U1582 ( .C1(n1454), .C2(n834), .A(n791), .B(n790), .ZN(\DP/A[20] )
         );
  AOI22_X1 U1583 ( .A1(n1494), .A2(\DP/RegLMD_out[21] ), .B1(
        \DP/RegALU2_out[21] ), .B2(n638), .ZN(n1237) );
  AOI22_X1 U1584 ( .A1(\DP/RegALU1_out[21] ), .A2(n829), .B1(\DP/RegA_out[21] ), .B2(n619), .ZN(n793) );
  NAND2_X1 U1585 ( .A1(n620), .A2(\DP/NPC2[21] ), .ZN(n792) );
  OAI211_X1 U1586 ( .C1(n1319), .C2(n834), .A(n793), .B(n792), .ZN(\DP/A[21] )
         );
  AOI22_X1 U1587 ( .A1(n639), .A2(\DP/RegLMD_out[22] ), .B1(
        \DP/RegALU2_out[22] ), .B2(n638), .ZN(n1239) );
  AOI22_X1 U1588 ( .A1(\DP/RegALU1_out[22] ), .A2(n829), .B1(\DP/RegA_out[22] ), .B2(n619), .ZN(n795) );
  NAND2_X1 U1589 ( .A1(n620), .A2(\DP/NPC2[22] ), .ZN(n794) );
  OAI211_X1 U1590 ( .C1(n1292), .C2(n621), .A(n795), .B(n794), .ZN(\DP/A[22] )
         );
  AOI22_X1 U1591 ( .A1(n1494), .A2(\DP/RegLMD_out[23] ), .B1(
        \DP/RegALU2_out[23] ), .B2(n638), .ZN(n1241) );
  AOI22_X1 U1592 ( .A1(\DP/RegALU1_out[23] ), .A2(n829), .B1(\DP/RegA_out[23] ), .B2(n830), .ZN(n797) );
  NAND2_X1 U1593 ( .A1(n620), .A2(\DP/NPC2[23] ), .ZN(n796) );
  OAI211_X1 U1594 ( .C1(n1433), .C2(n834), .A(n797), .B(n796), .ZN(\DP/A[23] )
         );
  AOI22_X1 U1595 ( .A1(n1494), .A2(\DP/RegLMD_out[24] ), .B1(
        \DP/RegALU2_out[24] ), .B2(n638), .ZN(n1243) );
  AOI22_X1 U1596 ( .A1(\DP/RegALU1_out[24] ), .A2(n829), .B1(\DP/RegA_out[24] ), .B2(n619), .ZN(n799) );
  NAND2_X1 U1597 ( .A1(n620), .A2(\DP/NPC2[24] ), .ZN(n798) );
  OAI211_X1 U1598 ( .C1(n1318), .C2(n621), .A(n799), .B(n798), .ZN(\DP/A[24] )
         );
  AOI22_X1 U1599 ( .A1(n639), .A2(\DP/RegLMD_out[25] ), .B1(
        \DP/RegALU2_out[25] ), .B2(n638), .ZN(n1245) );
  AOI22_X1 U1600 ( .A1(\DP/RegALU1_out[25] ), .A2(n829), .B1(\DP/RegA_out[25] ), .B2(n619), .ZN(n801) );
  NAND2_X1 U1601 ( .A1(n620), .A2(\DP/NPC2[25] ), .ZN(n800) );
  OAI211_X1 U1602 ( .C1(n1453), .C2(n834), .A(n801), .B(n800), .ZN(\DP/A[25] )
         );
  AOI22_X1 U1603 ( .A1(n639), .A2(\DP/RegLMD_out[26] ), .B1(
        \DP/RegALU2_out[26] ), .B2(n638), .ZN(n1247) );
  AOI22_X1 U1604 ( .A1(\DP/RegALU1_out[26] ), .A2(n829), .B1(\DP/RegA_out[26] ), .B2(n619), .ZN(n803) );
  NAND2_X1 U1605 ( .A1(n620), .A2(\DP/NPC2[26] ), .ZN(n802) );
  OAI211_X1 U1606 ( .C1(n1247), .C2(n621), .A(n803), .B(n802), .ZN(\DP/A[26] )
         );
  AOI22_X1 U1607 ( .A1(n1364), .A2(\DP/RegLMD_out[27] ), .B1(
        \DP/RegALU2_out[27] ), .B2(n638), .ZN(n1249) );
  AOI22_X1 U1608 ( .A1(\DP/RegALU1_out[27] ), .A2(n618), .B1(\DP/RegA_out[27] ), .B2(n619), .ZN(n805) );
  NAND2_X1 U1609 ( .A1(n620), .A2(\DP/NPC2[27] ), .ZN(n804) );
  OAI211_X1 U1610 ( .C1(n1458), .C2(n834), .A(n805), .B(n804), .ZN(\DP/A[27] )
         );
  AOI22_X1 U1612 ( .A1(\DP/RegALU1_out[28] ), .A2(n829), .B1(\DP/RegA_out[28] ), .B2(n619), .ZN(n807) );
  NAND2_X1 U1613 ( .A1(n620), .A2(\DP/NPC2[28] ), .ZN(n806) );
  OAI211_X1 U1614 ( .C1(n1305), .C2(n621), .A(n807), .B(n806), .ZN(\DP/A[28] )
         );
  AOI22_X1 U1615 ( .A1(n1494), .A2(\DP/RegLMD_out[29] ), .B1(
        \DP/RegALU2_out[29] ), .B2(n583), .ZN(n1253) );
  AOI22_X1 U1616 ( .A1(\DP/RegALU1_out[29] ), .A2(n618), .B1(\DP/RegA_out[29] ), .B2(n619), .ZN(n809) );
  NAND2_X1 U1617 ( .A1(n620), .A2(\DP/NPC2[29] ), .ZN(n808) );
  OAI211_X1 U1618 ( .C1(n1253), .C2(n834), .A(n809), .B(n808), .ZN(\DP/A[29] )
         );
  AOI22_X1 U1620 ( .A1(\DP/RegA_out[2] ), .A2(n830), .B1(DRAM_ADDR[2]), .B2(
        n618), .ZN(n811) );
  NAND2_X1 U1621 ( .A1(n831), .A2(\DP/NPC2[2] ), .ZN(n810) );
  AOI22_X1 U1623 ( .A1(n1494), .A2(\DP/RegLMD_out[30] ), .B1(
        \DP/RegALU2_out[30] ), .B2(n583), .ZN(n1255) );
  AOI22_X1 U1624 ( .A1(\DP/RegALU1_out[30] ), .A2(n829), .B1(\DP/RegA_out[30] ), .B2(n619), .ZN(n813) );
  NAND2_X1 U1625 ( .A1(n831), .A2(\DP/NPC2[30] ), .ZN(n812) );
  OAI211_X1 U1626 ( .C1(n1255), .C2(n834), .A(n813), .B(n812), .ZN(\DP/A[30] )
         );
  AOI22_X1 U1628 ( .A1(\DP/RegALU1_out[31] ), .A2(n618), .B1(\DP/RegA_out[31] ), .B2(n619), .ZN(n815) );
  NAND2_X1 U1629 ( .A1(n831), .A2(\DP/NPC2[31] ), .ZN(n814) );
  OAI211_X1 U1630 ( .C1(n1356), .C2(n621), .A(n815), .B(n814), .ZN(\DP/A[31] )
         );
  AOI22_X1 U1631 ( .A1(n639), .A2(\DP/RegLMD_out[3] ), .B1(\DP/RegALU2_out[3] ), .B2(n638), .ZN(n1274) );
  AOI22_X1 U1632 ( .A1(\DP/RegA_out[3] ), .A2(n830), .B1(DRAM_ADDR[3]), .B2(
        n618), .ZN(n817) );
  NAND2_X1 U1633 ( .A1(n831), .A2(\DP/NPC2[3] ), .ZN(n816) );
  OAI211_X1 U1634 ( .C1(n1449), .C2(n834), .A(n817), .B(n816), .ZN(\DP/A[3] )
         );
  AOI22_X1 U1635 ( .A1(n1494), .A2(\DP/RegLMD_out[4] ), .B1(
        \DP/RegALU2_out[4] ), .B2(n583), .ZN(n1275) );
  AOI22_X1 U1636 ( .A1(\DP/RegA_out[4] ), .A2(n830), .B1(DRAM_ADDR[4]), .B2(
        n618), .ZN(n819) );
  NAND2_X1 U1637 ( .A1(n620), .A2(\DP/NPC2[4] ), .ZN(n818) );
  OAI211_X1 U1638 ( .C1(n1367), .C2(n621), .A(n819), .B(n818), .ZN(\DP/A[4] )
         );
  AOI22_X1 U1639 ( .A1(n639), .A2(\DP/RegLMD_out[5] ), .B1(\DP/RegALU2_out[5] ), .B2(n638), .ZN(n1276) );
  AOI22_X1 U1640 ( .A1(\DP/RegA_out[5] ), .A2(n830), .B1(DRAM_ADDR[5]), .B2(
        n618), .ZN(n821) );
  NAND2_X1 U1641 ( .A1(n831), .A2(\DP/NPC2[5] ), .ZN(n820) );
  OAI211_X1 U1642 ( .C1(n1415), .C2(n621), .A(n821), .B(n820), .ZN(\DP/A[5] )
         );
  AOI22_X1 U1644 ( .A1(\DP/RegA_out[6] ), .A2(n830), .B1(DRAM_ADDR[6]), .B2(
        n618), .ZN(n823) );
  NAND2_X1 U1645 ( .A1(n620), .A2(\DP/NPC2[6] ), .ZN(n822) );
  AOI22_X1 U1647 ( .A1(\DP/RegA_out[7] ), .A2(n830), .B1(DRAM_ADDR[7]), .B2(
        n618), .ZN(n826) );
  MUX2_X1 U1648 ( .A(\DP/RegLMD_out[7] ), .B(\DP/RegALU2_out[7] ), .S(n583), 
        .Z(n1210) );
  AOI22_X1 U1649 ( .A1(\DP/NPC2[7] ), .A2(n831), .B1(n824), .B2(n1210), .ZN(
        n825) );
  NAND2_X1 U1650 ( .A1(n826), .A2(n825), .ZN(\DP/A[7] ) );
  AOI22_X1 U1651 ( .A1(n639), .A2(\DP/RegLMD_out[8] ), .B1(\DP/RegALU2_out[8] ), .B2(n583), .ZN(n1265) );
  AOI22_X1 U1652 ( .A1(\DP/RegA_out[8] ), .A2(n619), .B1(DRAM_ADDR[8]), .B2(
        n618), .ZN(n828) );
  NAND2_X1 U1653 ( .A1(n831), .A2(\DP/NPC2[8] ), .ZN(n827) );
  OAI211_X1 U1654 ( .C1(n1471), .C2(n621), .A(n828), .B(n827), .ZN(\DP/A[8] )
         );
  AOI22_X1 U1655 ( .A1(n639), .A2(\DP/RegLMD_out[9] ), .B1(\DP/RegALU2_out[9] ), .B2(n638), .ZN(n1270) );
  AOI22_X1 U1656 ( .A1(\DP/RegA_out[9] ), .A2(n830), .B1(DRAM_ADDR[9]), .B2(
        n618), .ZN(n833) );
  NAND2_X1 U1657 ( .A1(n620), .A2(\DP/NPC2[9] ), .ZN(n832) );
  OAI211_X1 U1658 ( .C1(n1270), .C2(n621), .A(n833), .B(n832), .ZN(\DP/A[9] )
         );
  INV_X1 U1659 ( .A(n942), .ZN(n1271) );
  NAND3_X1 U1660 ( .A1(n75), .A2(\DP/FwdB[0] ), .A3(n604), .ZN(n835) );
  AOI22_X1 U1661 ( .A1(DRAM_ADDR[0]), .A2(n624), .B1(\DP/RegB_out[0] ), .B2(
        n892), .ZN(n837) );
  NAND2_X1 U1662 ( .A1(n625), .A2(\DP/RegIMM_out[0] ), .ZN(n836) );
  OAI211_X1 U1663 ( .C1(n1271), .C2(n626), .A(n837), .B(n836), .ZN(\DP/B[0] )
         );
  AOI22_X1 U1664 ( .A1(DRAM_ADDR[10]), .A2(n623), .B1(n622), .B2(
        \DP/RegB_out[10] ), .ZN(n839) );
  NAND2_X1 U1665 ( .A1(n894), .A2(\DP/RegIMM_out[10] ), .ZN(n838) );
  OAI211_X1 U1666 ( .C1(n1501), .C2(n897), .A(n839), .B(n838), .ZN(\DP/B[10] )
         );
  AOI22_X1 U1667 ( .A1(DRAM_ADDR[11]), .A2(n624), .B1(n892), .B2(
        \DP/RegB_out[11] ), .ZN(n841) );
  NAND2_X1 U1668 ( .A1(n625), .A2(\DP/RegIMM_out[11] ), .ZN(n840) );
  OAI211_X1 U1669 ( .C1(n1214), .C2(n626), .A(n841), .B(n840), .ZN(\DP/B[11] )
         );
  AOI22_X1 U1670 ( .A1(\DP/RegALU1_out[12] ), .A2(n624), .B1(n622), .B2(
        \DP/RegB_out[12] ), .ZN(n843) );
  NAND2_X1 U1671 ( .A1(n894), .A2(\DP/RegIMM_out[12] ), .ZN(n842) );
  OAI211_X1 U1672 ( .C1(n1216), .C2(n897), .A(n843), .B(n842), .ZN(\DP/B[12] )
         );
  AOI22_X1 U1673 ( .A1(\DP/RegALU1_out[13] ), .A2(n624), .B1(n892), .B2(
        \DP/RegB_out[13] ), .ZN(n845) );
  NAND2_X1 U1674 ( .A1(n625), .A2(\DP/RegIMM_out[13] ), .ZN(n844) );
  OAI211_X1 U1675 ( .C1(n1218), .C2(n626), .A(n845), .B(n844), .ZN(\DP/B[13] )
         );
  AOI22_X1 U1676 ( .A1(\DP/RegALU1_out[14] ), .A2(n624), .B1(n622), .B2(
        \DP/RegB_out[14] ), .ZN(n847) );
  NAND2_X1 U1677 ( .A1(n894), .A2(\DP/RegIMM_out[14] ), .ZN(n846) );
  OAI211_X1 U1678 ( .C1(n1462), .C2(n897), .A(n847), .B(n846), .ZN(\DP/B[14] )
         );
  AOI22_X1 U1679 ( .A1(\DP/RegALU1_out[15] ), .A2(n624), .B1(n892), .B2(
        \DP/RegB_out[15] ), .ZN(n849) );
  NAND2_X1 U1680 ( .A1(n625), .A2(\DP/RegIMM_out[15] ), .ZN(n848) );
  OAI211_X1 U1681 ( .C1(n985), .C2(n897), .A(n849), .B(n848), .ZN(\DP/B[15] )
         );
  AOI22_X1 U1682 ( .A1(\DP/RegALU1_out[16] ), .A2(n893), .B1(n892), .B2(
        \DP/RegB_out[16] ), .ZN(n851) );
  NAND2_X1 U1683 ( .A1(n894), .A2(\DP/RegIMM_out[16] ), .ZN(n850) );
  OAI211_X1 U1684 ( .C1(n1227), .C2(n897), .A(n851), .B(n850), .ZN(\DP/B[16] )
         );
  AOI22_X1 U1685 ( .A1(\DP/RegALU1_out[17] ), .A2(n893), .B1(n892), .B2(
        \DP/RegB_out[17] ), .ZN(n853) );
  NAND2_X1 U1686 ( .A1(n625), .A2(\DP/RegIMM_out[17] ), .ZN(n852) );
  OAI211_X1 U1687 ( .C1(n1361), .C2(n897), .A(n853), .B(n852), .ZN(\DP/B[17] )
         );
  AOI22_X1 U1688 ( .A1(\DP/RegALU1_out[18] ), .A2(n893), .B1(n892), .B2(
        \DP/RegB_out[18] ), .ZN(n855) );
  NAND2_X1 U1689 ( .A1(n894), .A2(\DP/RegIMM_out[18] ), .ZN(n854) );
  OAI211_X1 U1690 ( .C1(n1336), .C2(n897), .A(n855), .B(n854), .ZN(\DP/B[18] )
         );
  AOI22_X1 U1691 ( .A1(\DP/RegALU1_out[19] ), .A2(n893), .B1(n892), .B2(
        \DP/RegB_out[19] ), .ZN(n857) );
  NAND2_X1 U1692 ( .A1(n625), .A2(\DP/RegIMM_out[19] ), .ZN(n856) );
  OAI211_X1 U1693 ( .C1(n1233), .C2(n897), .A(n857), .B(n856), .ZN(\DP/B[19] )
         );
  AOI22_X1 U1694 ( .A1(DRAM_ADDR[1]), .A2(n893), .B1(n892), .B2(
        \DP/RegB_out[1] ), .ZN(n859) );
  NAND2_X1 U1695 ( .A1(n894), .A2(\DP/RegIMM_out[1] ), .ZN(n858) );
  OAI211_X1 U1696 ( .C1(n1272), .C2(n897), .A(n859), .B(n858), .ZN(\DP/B[1] )
         );
  AOI22_X1 U1697 ( .A1(\DP/RegALU1_out[20] ), .A2(n623), .B1(n622), .B2(
        \DP/RegB_out[20] ), .ZN(n861) );
  NAND2_X1 U1698 ( .A1(n625), .A2(\DP/RegIMM_out[20] ), .ZN(n860) );
  OAI211_X1 U1699 ( .C1(n1454), .C2(n897), .A(n861), .B(n860), .ZN(\DP/B[20] )
         );
  AOI22_X1 U1700 ( .A1(\DP/RegALU1_out[21] ), .A2(n623), .B1(n622), .B2(
        \DP/RegB_out[21] ), .ZN(n863) );
  NAND2_X1 U1701 ( .A1(n625), .A2(\DP/RegIMM_out[21] ), .ZN(n862) );
  OAI211_X1 U1702 ( .C1(n1319), .C2(n626), .A(n863), .B(n862), .ZN(\DP/B[21] )
         );
  AOI22_X1 U1703 ( .A1(\DP/RegALU1_out[22] ), .A2(n623), .B1(n622), .B2(
        \DP/RegB_out[22] ), .ZN(n865) );
  NAND2_X1 U1704 ( .A1(n625), .A2(\DP/RegIMM_out[22] ), .ZN(n864) );
  OAI211_X1 U1705 ( .C1(n1292), .C2(n897), .A(n865), .B(n864), .ZN(\DP/B[22] )
         );
  AOI22_X1 U1706 ( .A1(\DP/RegALU1_out[23] ), .A2(n623), .B1(n622), .B2(
        \DP/RegB_out[23] ), .ZN(n867) );
  NAND2_X1 U1707 ( .A1(n625), .A2(\DP/RegIMM_out[23] ), .ZN(n866) );
  OAI211_X1 U1708 ( .C1(n1433), .C2(n626), .A(n867), .B(n866), .ZN(\DP/B[23] )
         );
  AOI22_X1 U1709 ( .A1(\DP/RegALU1_out[24] ), .A2(n623), .B1(n622), .B2(
        \DP/RegB_out[24] ), .ZN(n869) );
  NAND2_X1 U1710 ( .A1(n894), .A2(\DP/RegIMM_out[24] ), .ZN(n868) );
  OAI211_X1 U1711 ( .C1(n1318), .C2(n897), .A(n869), .B(n868), .ZN(\DP/B[24] )
         );
  AOI22_X1 U1712 ( .A1(\DP/RegALU1_out[25] ), .A2(n623), .B1(n622), .B2(
        \DP/RegB_out[25] ), .ZN(n870) );
  NAND2_X1 U1713 ( .A1(n625), .A2(\DP/RegIMM_out[31] ), .ZN(n878) );
  OAI211_X1 U1714 ( .C1(n1453), .C2(n626), .A(n870), .B(n878), .ZN(\DP/B[25] )
         );
  AOI22_X1 U1715 ( .A1(\DP/RegALU1_out[26] ), .A2(n623), .B1(n622), .B2(
        \DP/RegB_out[26] ), .ZN(n871) );
  OAI211_X1 U1716 ( .C1(n1247), .C2(n897), .A(n871), .B(n878), .ZN(\DP/B[26] )
         );
  AOI22_X1 U1717 ( .A1(\DP/RegALU1_out[27] ), .A2(n623), .B1(n622), .B2(
        \DP/RegB_out[27] ), .ZN(n872) );
  OAI211_X1 U1718 ( .C1(n1458), .C2(n626), .A(n872), .B(n878), .ZN(\DP/B[27] )
         );
  AOI22_X1 U1719 ( .A1(\DP/RegALU1_out[28] ), .A2(n623), .B1(n892), .B2(
        \DP/RegB_out[28] ), .ZN(n873) );
  OAI211_X1 U1720 ( .C1(n1305), .C2(n897), .A(n873), .B(n878), .ZN(\DP/B[28] )
         );
  AOI22_X1 U1721 ( .A1(\DP/RegALU1_out[29] ), .A2(n623), .B1(n622), .B2(
        \DP/RegB_out[29] ), .ZN(n874) );
  OAI211_X1 U1722 ( .C1(n1253), .C2(n626), .A(n874), .B(n878), .ZN(\DP/B[29] )
         );
  AOI22_X1 U1723 ( .A1(DRAM_ADDR[2]), .A2(n623), .B1(n892), .B2(
        \DP/RegB_out[2] ), .ZN(n876) );
  NAND2_X1 U1724 ( .A1(n894), .A2(\DP/RegIMM_out[2] ), .ZN(n875) );
  AOI22_X1 U1726 ( .A1(\DP/RegALU1_out[30] ), .A2(n623), .B1(n892), .B2(
        \DP/RegB_out[30] ), .ZN(n877) );
  OAI211_X1 U1727 ( .C1(n1255), .C2(n897), .A(n877), .B(n878), .ZN(\DP/B[30] )
         );
  AOI22_X1 U1728 ( .A1(\DP/RegALU1_out[31] ), .A2(n624), .B1(n622), .B2(
        \DP/RegB_out[31] ), .ZN(n879) );
  OAI211_X1 U1729 ( .C1(n1356), .C2(n626), .A(n879), .B(n878), .ZN(\DP/B[31] )
         );
  AOI22_X1 U1730 ( .A1(DRAM_ADDR[3]), .A2(n624), .B1(n622), .B2(
        \DP/RegB_out[3] ), .ZN(n881) );
  NAND2_X1 U1731 ( .A1(n625), .A2(\DP/RegIMM_out[3] ), .ZN(n880) );
  OAI211_X1 U1732 ( .C1(n1449), .C2(n626), .A(n881), .B(n880), .ZN(\DP/B[3] )
         );
  AOI22_X1 U1733 ( .A1(DRAM_ADDR[4]), .A2(n624), .B1(n622), .B2(
        \DP/RegB_out[4] ), .ZN(n883) );
  NAND2_X1 U1734 ( .A1(n894), .A2(\DP/RegIMM_out[4] ), .ZN(n882) );
  OAI211_X1 U1735 ( .C1(n1367), .C2(n626), .A(n883), .B(n882), .ZN(\DP/B[4] )
         );
  AOI22_X1 U1736 ( .A1(DRAM_ADDR[5]), .A2(n624), .B1(n622), .B2(
        \DP/RegB_out[5] ), .ZN(n885) );
  NAND2_X1 U1737 ( .A1(n625), .A2(\DP/RegIMM_out[5] ), .ZN(n884) );
  OAI211_X1 U1738 ( .C1(n1415), .C2(n626), .A(n885), .B(n884), .ZN(\DP/B[5] )
         );
  AOI22_X1 U1739 ( .A1(DRAM_ADDR[6]), .A2(n624), .B1(n622), .B2(
        \DP/RegB_out[6] ), .ZN(n887) );
  NAND2_X1 U1740 ( .A1(n894), .A2(\DP/RegIMM_out[6] ), .ZN(n886) );
  INV_X1 U1742 ( .A(n1210), .ZN(n1263) );
  AOI22_X1 U1743 ( .A1(DRAM_ADDR[7]), .A2(n624), .B1(n622), .B2(
        \DP/RegB_out[7] ), .ZN(n889) );
  NAND2_X1 U1744 ( .A1(n894), .A2(\DP/RegIMM_out[7] ), .ZN(n888) );
  OAI211_X1 U1745 ( .C1(n1263), .C2(n626), .A(n889), .B(n888), .ZN(\DP/B[7] )
         );
  AOI22_X1 U1746 ( .A1(DRAM_ADDR[8]), .A2(n624), .B1(n622), .B2(
        \DP/RegB_out[8] ), .ZN(n891) );
  NAND2_X1 U1747 ( .A1(n625), .A2(\DP/RegIMM_out[8] ), .ZN(n890) );
  OAI211_X1 U1748 ( .C1(n1471), .C2(n626), .A(n891), .B(n890), .ZN(\DP/B[8] )
         );
  AOI22_X1 U1749 ( .A1(DRAM_ADDR[9]), .A2(n624), .B1(n622), .B2(
        \DP/RegB_out[9] ), .ZN(n896) );
  NAND2_X1 U1750 ( .A1(n625), .A2(\DP/RegIMM_out[9] ), .ZN(n895) );
  OAI211_X1 U1751 ( .C1(n1456), .C2(n626), .A(n896), .B(n895), .ZN(\DP/B[9] )
         );
  NAND2_X1 U1752 ( .A1(n59), .A2(n1056), .ZN(\DP/FFDBRANCH/N2 ) );
  NOR2_X1 U1753 ( .A1(n641), .A2(n590), .ZN(\DP/FFDJL1/N3 ) );
  NOR2_X1 U1754 ( .A1(n58), .A2(n641), .ZN(\DP/FFDJREG/N3 ) );
  NAND4_X1 U1759 ( .A1(n1239), .A2(n1237), .A3(n1235), .A4(n1233), .ZN(n902)
         );
  NAND4_X1 U1760 ( .A1(n1247), .A2(n1245), .A3(n1243), .A4(n1433), .ZN(n901)
         );
  NAND4_X1 U1761 ( .A1(n1218), .A2(n1216), .A3(n1214), .A4(n1212), .ZN(n900)
         );
  NAND4_X1 U1762 ( .A1(n1231), .A2(n1229), .A3(n1227), .A4(n1462), .ZN(n899)
         );
  NAND3_X1 U1766 ( .A1(n77), .A2(n76), .A3(\DP/FwdC[1] ), .ZN(n974) );
  NOR4_X1 U1767 ( .A1(\DP/RegA_out[18] ), .A2(\DP/RegA_out[17] ), .A3(
        \DP/RegA_out[16] ), .A4(\DP/RegA_out[15] ), .ZN(n911) );
  NAND4_X1 U1776 ( .A1(n915), .A2(n914), .A3(n913), .A4(n912), .ZN(n916) );
  NOR3_X1 U1777 ( .A1(n76), .A2(\DP/FwdC[1] ), .A3(\DP/FwdA[2] ), .ZN(n975) );
  OAI21_X1 U1778 ( .B1(n917), .B2(n916), .A(n975), .ZN(n929) );
  NOR4_X1 U1784 ( .A1(\DP/RegALU1_out[31] ), .A2(\DP/RegALU1_out[30] ), .A3(
        DRAM_ADDR[2]), .A4(DRAM_ADDR[1]), .ZN(n925) );
  NOR4_X1 U1785 ( .A1(DRAM_ADDR[6]), .A2(DRAM_ADDR[5]), .A3(DRAM_ADDR[4]), 
        .A4(DRAM_ADDR[3]), .ZN(n924) );
  NAND2_X1 U1796 ( .A1(n935), .A2(RST), .ZN(\DP/RegNPC1/N2 ) );
  NAND2_X1 U1798 ( .A1(n1495), .A2(IR_OUT[20]), .ZN(n1208) );
  NAND2_X1 U1799 ( .A1(n1495), .A2(IR_OUT[19]), .ZN(n1206) );
  NAND2_X1 U1800 ( .A1(n1495), .A2(IR_OUT[17]), .ZN(n1204) );
  NAND2_X1 U1801 ( .A1(n1495), .A2(IR_OUT[16]), .ZN(n1203) );
  NOR4_X1 U1802 ( .A1(\DP/RD2[1] ), .A2(\DP/RD2[0] ), .A3(n593), .A4(n584), 
        .ZN(n936) );
  AOI21_X1 U1803 ( .B1(n936), .B2(n585), .A(n601), .ZN(n1020) );
  AOI22_X1 U1808 ( .A1(n1295), .A2(n585), .B1(\DP/RD2[2] ), .B2(n1205), .ZN(
        n940) );
  NAND2_X1 U1809 ( .A1(n941), .A2(n940), .ZN(n1035) );
  NOR2_X1 U1810 ( .A1(n640), .A2(n1035), .ZN(\DP/FFDFD/N3 ) );
  NAND2_X1 U1811 ( .A1(RST), .A2(n590), .ZN(\DP/RegNPC2/N2 ) );
  NAND2_X1 U1812 ( .A1(n1056), .A2(n590), .ZN(\DP/FFDJL2/N2 ) );
  AND2_X1 U1813 ( .A1(RST), .A2(\DP/JL1 ), .ZN(\DP/FFDJL2/N3 ) );
  NAND2_X1 U1814 ( .A1(n58), .A2(n1056), .ZN(\DP/RegA1/N2 ) );
  NAND2_X1 U1816 ( .A1(n1492), .A2(\DP/NPC_out[10] ), .ZN(n943) );
  NAND2_X1 U1818 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[11] ), .ZN(n944) );
  OAI21_X1 U1819 ( .B1(\DP/JL2 ), .B2(n1214), .A(n944), .ZN(\DP/RF_DATA[11] )
         );
  NAND2_X1 U1820 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[12] ), .ZN(n945) );
  OAI21_X1 U1821 ( .B1(n1488), .B2(n1216), .A(n945), .ZN(\DP/RF_DATA[12] ) );
  NAND2_X1 U1822 ( .A1(n1492), .A2(\DP/NPC_out[13] ), .ZN(n946) );
  OAI21_X1 U1823 ( .B1(n1488), .B2(n1218), .A(n946), .ZN(\DP/RF_DATA[13] ) );
  NAND2_X1 U1824 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[14] ), .ZN(n947) );
  MUX2_X1 U1825 ( .A(n1221), .B(\DP/NPC_out[15] ), .S(\DP/JL2 ), .Z(
        \DP/RF_DATA[15] ) );
  NAND2_X1 U1826 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[16] ), .ZN(n948) );
  NAND2_X1 U1829 ( .A1(n1488), .A2(\DP/NPC_out[18] ), .ZN(n950) );
  NAND2_X1 U1830 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[19] ), .ZN(n951) );
  OAI21_X1 U1831 ( .B1(\DP/JL2 ), .B2(n1233), .A(n951), .ZN(\DP/RF_DATA[19] )
         );
  NAND2_X1 U1832 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[1] ), .ZN(n952) );
  OAI21_X1 U1833 ( .B1(\DP/JL2 ), .B2(n1272), .A(n952), .ZN(\DP/RF_DATA[1] )
         );
  NAND2_X1 U1836 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[21] ), .ZN(n954) );
  NAND2_X1 U1837 ( .A1(n1492), .A2(\DP/NPC_out[22] ), .ZN(n955) );
  NAND2_X1 U1838 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[23] ), .ZN(n956) );
  NAND2_X1 U1839 ( .A1(n1488), .A2(\DP/NPC_out[24] ), .ZN(n957) );
  NAND2_X1 U1840 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[25] ), .ZN(n958) );
  NAND2_X1 U1842 ( .A1(n1488), .A2(\DP/NPC_out[26] ), .ZN(n959) );
  NAND2_X1 U1843 ( .A1(n1492), .A2(\DP/NPC_out[27] ), .ZN(n960) );
  NAND2_X1 U1844 ( .A1(n1492), .A2(\DP/NPC_out[28] ), .ZN(n961) );
  NAND2_X1 U1846 ( .A1(n1488), .A2(\DP/NPC_out[29] ), .ZN(n962) );
  OAI21_X1 U1847 ( .B1(\DP/JL2 ), .B2(n1253), .A(n962), .ZN(\DP/RF_DATA[29] )
         );
  NAND2_X1 U1850 ( .A1(n1488), .A2(\DP/NPC_out[31] ), .ZN(n965) );
  NAND2_X1 U1852 ( .A1(n1492), .A2(\DP/NPC_out[3] ), .ZN(n966) );
  OAI21_X1 U1855 ( .B1(n1488), .B2(n1275), .A(n967), .ZN(\DP/RF_DATA[4] ) );
  NAND2_X1 U1858 ( .A1(n1488), .A2(\DP/NPC_out[6] ), .ZN(n969) );
  MUX2_X1 U1859 ( .A(n1210), .B(\DP/NPC_out[7] ), .S(\DP/JL2 ), .Z(
        \DP/RF_DATA[7] ) );
  NAND2_X1 U1860 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[8] ), .ZN(n970) );
  NAND2_X1 U1862 ( .A1(n1492), .A2(\DP/NPC_out[9] ), .ZN(n971) );
  AND2_X1 U1864 ( .A1(RST), .A2(\DP/RegA_in[7] ), .ZN(\DP/RegA/N10 ) );
  AND2_X1 U1865 ( .A1(RST), .A2(\DP/RegA_in[8] ), .ZN(\DP/RegA/N11 ) );
  AND2_X1 U1866 ( .A1(RST), .A2(\DP/RegA_in[9] ), .ZN(\DP/RegA/N12 ) );
  AND2_X1 U1867 ( .A1(RST), .A2(\DP/RegA_in[10] ), .ZN(\DP/RegA/N13 ) );
  AND2_X1 U1868 ( .A1(RST), .A2(\DP/RegA_in[11] ), .ZN(\DP/RegA/N14 ) );
  AND2_X1 U1869 ( .A1(RST), .A2(\DP/RegA_in[12] ), .ZN(\DP/RegA/N15 ) );
  AND2_X1 U1870 ( .A1(RST), .A2(\DP/RegA_in[13] ), .ZN(\DP/RegA/N16 ) );
  AND2_X1 U1871 ( .A1(RST), .A2(\DP/RegA_in[14] ), .ZN(\DP/RegA/N17 ) );
  AND2_X1 U1872 ( .A1(RST), .A2(\DP/RegA_in[15] ), .ZN(\DP/RegA/N18 ) );
  AND2_X1 U1873 ( .A1(RST), .A2(\DP/RegA_in[16] ), .ZN(\DP/RegA/N19 ) );
  AND2_X1 U1875 ( .A1(RST), .A2(\DP/RegA_in[17] ), .ZN(\DP/RegA/N20 ) );
  AND2_X1 U1876 ( .A1(RST), .A2(\DP/RegA_in[18] ), .ZN(\DP/RegA/N21 ) );
  AND2_X1 U1877 ( .A1(RST), .A2(\DP/RegA_in[19] ), .ZN(\DP/RegA/N22 ) );
  AND2_X1 U1878 ( .A1(RST), .A2(\DP/RegA_in[20] ), .ZN(\DP/RegA/N23 ) );
  AND2_X1 U1879 ( .A1(RST), .A2(\DP/RegA_in[21] ), .ZN(\DP/RegA/N24 ) );
  AND2_X1 U1880 ( .A1(RST), .A2(\DP/RegA_in[22] ), .ZN(\DP/RegA/N25 ) );
  AND2_X1 U1881 ( .A1(RST), .A2(\DP/RegA_in[23] ), .ZN(\DP/RegA/N26 ) );
  AND2_X1 U1882 ( .A1(RST), .A2(\DP/RegA_in[24] ), .ZN(\DP/RegA/N27 ) );
  AND2_X1 U1883 ( .A1(RST), .A2(\DP/RegA_in[25] ), .ZN(\DP/RegA/N28 ) );
  AND2_X1 U1884 ( .A1(RST), .A2(\DP/RegA_in[26] ), .ZN(\DP/RegA/N29 ) );
  AND2_X1 U1885 ( .A1(RST), .A2(\DP/RegA_in[0] ), .ZN(\DP/RegA/N3 ) );
  AND2_X1 U1886 ( .A1(RST), .A2(\DP/RegA_in[27] ), .ZN(\DP/RegA/N30 ) );
  AND2_X1 U1887 ( .A1(RST), .A2(\DP/RegA_in[28] ), .ZN(\DP/RegA/N31 ) );
  AND2_X1 U1888 ( .A1(RST), .A2(\DP/RegA_in[29] ), .ZN(\DP/RegA/N32 ) );
  AND2_X1 U1889 ( .A1(RST), .A2(\DP/RegA_in[30] ), .ZN(\DP/RegA/N33 ) );
  AND2_X1 U1890 ( .A1(RST), .A2(\DP/RegA_in[31] ), .ZN(\DP/RegA/N34 ) );
  AND2_X1 U1891 ( .A1(RST), .A2(\DP/RegA_in[1] ), .ZN(\DP/RegA/N4 ) );
  AND2_X1 U1892 ( .A1(RST), .A2(\DP/RegA_in[2] ), .ZN(\DP/RegA/N5 ) );
  AND2_X1 U1893 ( .A1(RST), .A2(\DP/RegA_in[3] ), .ZN(\DP/RegA/N6 ) );
  AND2_X1 U1894 ( .A1(RST), .A2(\DP/RegA_in[4] ), .ZN(\DP/RegA/N7 ) );
  AND2_X1 U1895 ( .A1(RST), .A2(\DP/RegA_in[5] ), .ZN(\DP/RegA/N8 ) );
  AND2_X1 U1896 ( .A1(RST), .A2(\DP/RegA_in[6] ), .ZN(\DP/RegA/N9 ) );
  AOI22_X1 U1897 ( .A1(\DP/RegA_out[7] ), .A2(n629), .B1(n628), .B2(
        \DP/RegALU2/N10 ), .ZN(n976) );
  OAI21_X1 U1898 ( .B1(n1263), .B2(n630), .A(n976), .ZN(\DP/RegA1/N10 ) );
  AOI22_X1 U1899 ( .A1(\DP/RegA_out[8] ), .A2(n1009), .B1(n628), .B2(
        \DP/RegALU2/N11 ), .ZN(n977) );
  OAI21_X1 U1900 ( .B1(n1471), .B2(n1011), .A(n977), .ZN(\DP/RegA1/N11 ) );
  AOI22_X1 U1901 ( .A1(\DP/RegA_out[9] ), .A2(n1009), .B1(n628), .B2(
        \DP/RegALU2/N12 ), .ZN(n978) );
  OAI21_X1 U1902 ( .B1(n1270), .B2(n630), .A(n978), .ZN(\DP/RegA1/N12 ) );
  AOI22_X1 U1903 ( .A1(\DP/RegA_out[10] ), .A2(n1009), .B1(n628), .B2(
        \DP/RegALU2/N13 ), .ZN(n979) );
  OAI21_X1 U1904 ( .B1(n1501), .B2(n1011), .A(n979), .ZN(\DP/RegA1/N13 ) );
  AOI22_X1 U1905 ( .A1(\DP/RegA_out[11] ), .A2(n1009), .B1(n628), .B2(
        \DP/RegALU2/N14 ), .ZN(n980) );
  OAI21_X1 U1906 ( .B1(n1214), .B2(n630), .A(n980), .ZN(\DP/RegA1/N14 ) );
  AOI22_X1 U1907 ( .A1(\DP/RegA_out[12] ), .A2(n1009), .B1(n628), .B2(
        \DP/RegALU2/N15 ), .ZN(n981) );
  OAI21_X1 U1908 ( .B1(n1216), .B2(n1011), .A(n981), .ZN(\DP/RegA1/N15 ) );
  AOI22_X1 U1909 ( .A1(\DP/RegALU2/N16 ), .A2(n1008), .B1(\DP/RegA_out[13] ), 
        .B2(n629), .ZN(n982) );
  OAI21_X1 U1910 ( .B1(n1218), .B2(n1011), .A(n982), .ZN(\DP/RegA1/N16 ) );
  AOI22_X1 U1911 ( .A1(\DP/RegALU2/N17 ), .A2(n1008), .B1(\DP/RegA_out[14] ), 
        .B2(n1009), .ZN(n983) );
  OAI21_X1 U1912 ( .B1(n1462), .B2(n1011), .A(n983), .ZN(\DP/RegA1/N17 ) );
  AOI22_X1 U1913 ( .A1(\DP/RegALU2/N18 ), .A2(n628), .B1(\DP/RegA_out[15] ), 
        .B2(n1009), .ZN(n984) );
  OAI21_X1 U1914 ( .B1(n985), .B2(n1011), .A(n984), .ZN(\DP/RegA1/N18 ) );
  AOI22_X1 U1915 ( .A1(\DP/RegALU2/N19 ), .A2(n1008), .B1(\DP/RegA_out[16] ), 
        .B2(n629), .ZN(n986) );
  OAI21_X1 U1916 ( .B1(n1227), .B2(n1011), .A(n986), .ZN(\DP/RegA1/N19 ) );
  AOI22_X1 U1917 ( .A1(\DP/RegALU2/N20 ), .A2(n1008), .B1(\DP/RegA_out[17] ), 
        .B2(n1009), .ZN(n987) );
  OAI21_X1 U1918 ( .B1(n1361), .B2(n1011), .A(n987), .ZN(\DP/RegA1/N20 ) );
  AOI22_X1 U1919 ( .A1(\DP/RegALU2/N21 ), .A2(n628), .B1(\DP/RegA_out[18] ), 
        .B2(n629), .ZN(n988) );
  OAI21_X1 U1920 ( .B1(n1336), .B2(n1011), .A(n988), .ZN(\DP/RegA1/N21 ) );
  AOI22_X1 U1921 ( .A1(\DP/RegALU2/N22 ), .A2(n628), .B1(\DP/RegA_out[19] ), 
        .B2(n629), .ZN(n989) );
  OAI21_X1 U1922 ( .B1(n1233), .B2(n1011), .A(n989), .ZN(\DP/RegA1/N22 ) );
  AOI22_X1 U1923 ( .A1(\DP/RegALU2/N23 ), .A2(n628), .B1(\DP/RegA_out[20] ), 
        .B2(n1009), .ZN(n990) );
  OAI21_X1 U1924 ( .B1(n1454), .B2(n630), .A(n990), .ZN(\DP/RegA1/N23 ) );
  AOI22_X1 U1925 ( .A1(\DP/RegALU2/N24 ), .A2(n628), .B1(\DP/RegA_out[21] ), 
        .B2(n629), .ZN(n991) );
  OAI21_X1 U1926 ( .B1(n1319), .B2(n1011), .A(n991), .ZN(\DP/RegA1/N24 ) );
  AOI22_X1 U1927 ( .A1(\DP/RegALU2/N25 ), .A2(n628), .B1(\DP/RegA_out[22] ), 
        .B2(n629), .ZN(n992) );
  OAI21_X1 U1928 ( .B1(n1292), .B2(n630), .A(n992), .ZN(\DP/RegA1/N25 ) );
  AOI22_X1 U1929 ( .A1(\DP/RegALU2/N26 ), .A2(n628), .B1(\DP/RegA_out[23] ), 
        .B2(n1009), .ZN(n993) );
  OAI21_X1 U1930 ( .B1(n1433), .B2(n1011), .A(n993), .ZN(\DP/RegA1/N26 ) );
  AOI22_X1 U1931 ( .A1(\DP/RegALU2/N27 ), .A2(n628), .B1(\DP/RegA_out[24] ), 
        .B2(n629), .ZN(n994) );
  OAI21_X1 U1932 ( .B1(n1318), .B2(n630), .A(n994), .ZN(\DP/RegA1/N27 ) );
  AOI22_X1 U1933 ( .A1(\DP/RegALU2/N28 ), .A2(n628), .B1(\DP/RegA_out[25] ), 
        .B2(n1009), .ZN(n995) );
  OAI21_X1 U1934 ( .B1(n1453), .B2(n1011), .A(n995), .ZN(\DP/RegA1/N28 ) );
  AOI22_X1 U1935 ( .A1(\DP/RegALU2/N29 ), .A2(n628), .B1(\DP/RegA_out[26] ), 
        .B2(n629), .ZN(n996) );
  OAI21_X1 U1936 ( .B1(n1247), .B2(n630), .A(n996), .ZN(\DP/RegA1/N29 ) );
  AOI22_X1 U1937 ( .A1(\DP/RegA_out[0] ), .A2(n1009), .B1(n628), .B2(
        \DP/RegALU2/N3 ), .ZN(n997) );
  OAI21_X1 U1938 ( .B1(n1271), .B2(n1011), .A(n997), .ZN(\DP/RegA1/N3 ) );
  AOI22_X1 U1939 ( .A1(\DP/RegALU2/N30 ), .A2(n628), .B1(\DP/RegA_out[27] ), 
        .B2(n629), .ZN(n998) );
  OAI21_X1 U1940 ( .B1(n1458), .B2(n630), .A(n998), .ZN(\DP/RegA1/N30 ) );
  AOI22_X1 U1941 ( .A1(\DP/RegALU2/N31 ), .A2(n628), .B1(\DP/RegA_out[28] ), 
        .B2(n629), .ZN(n999) );
  OAI21_X1 U1942 ( .B1(n1305), .B2(n1011), .A(n999), .ZN(\DP/RegA1/N31 ) );
  AOI22_X1 U1943 ( .A1(\DP/RegALU2/N32 ), .A2(n628), .B1(\DP/RegA_out[29] ), 
        .B2(n629), .ZN(n1000) );
  OAI21_X1 U1944 ( .B1(n1253), .B2(n1011), .A(n1000), .ZN(\DP/RegA1/N32 ) );
  AOI22_X1 U1945 ( .A1(\DP/RegALU2/N33 ), .A2(n628), .B1(\DP/RegA_out[30] ), 
        .B2(n629), .ZN(n1001) );
  OAI21_X1 U1946 ( .B1(n1255), .B2(n630), .A(n1001), .ZN(\DP/RegA1/N33 ) );
  AOI22_X1 U1947 ( .A1(\DP/RegALU2/N34 ), .A2(n628), .B1(\DP/RegA_out[31] ), 
        .B2(n629), .ZN(n1002) );
  OAI21_X1 U1948 ( .B1(n1356), .B2(n630), .A(n1002), .ZN(\DP/RegA1/N34 ) );
  AOI22_X1 U1949 ( .A1(\DP/RegA_out[1] ), .A2(n1009), .B1(n628), .B2(
        \DP/RegALU2/N4 ), .ZN(n1003) );
  OAI21_X1 U1950 ( .B1(n1272), .B2(n630), .A(n1003), .ZN(\DP/RegA1/N4 ) );
  AOI22_X1 U1951 ( .A1(\DP/RegA_out[2] ), .A2(n1009), .B1(n628), .B2(
        \DP/RegALU2/N5 ), .ZN(n1004) );
  AOI22_X1 U1953 ( .A1(\DP/RegA_out[3] ), .A2(n1009), .B1(n628), .B2(
        \DP/RegALU2/N6 ), .ZN(n1005) );
  OAI21_X1 U1954 ( .B1(n1449), .B2(n630), .A(n1005), .ZN(\DP/RegA1/N6 ) );
  AOI22_X1 U1955 ( .A1(\DP/RegA_out[4] ), .A2(n629), .B1(n628), .B2(
        \DP/RegALU2/N7 ), .ZN(n1006) );
  OAI21_X1 U1956 ( .B1(n1367), .B2(n630), .A(n1006), .ZN(\DP/RegA1/N7 ) );
  AOI22_X1 U1957 ( .A1(\DP/RegA_out[5] ), .A2(n1009), .B1(n628), .B2(
        \DP/RegALU2/N8 ), .ZN(n1007) );
  OAI21_X1 U1958 ( .B1(n1415), .B2(n630), .A(n1007), .ZN(\DP/RegA1/N8 ) );
  AOI22_X1 U1959 ( .A1(\DP/RegA_out[6] ), .A2(n629), .B1(n628), .B2(
        \DP/RegALU2/N9 ), .ZN(n1010) );
  AND2_X1 U1961 ( .A1(RST), .A2(\DP/RES[7] ), .ZN(\DP/RegALU1/N10 ) );
  AND2_X1 U1962 ( .A1(RST), .A2(\DP/RES[9] ), .ZN(\DP/RegALU1/N12 ) );
  AND2_X1 U1963 ( .A1(RST), .A2(\DP/RES[10] ), .ZN(\DP/RegALU1/N13 ) );
  AND2_X1 U1964 ( .A1(RST), .A2(\DP/RES[11] ), .ZN(\DP/RegALU1/N14 ) );
  AND2_X1 U1965 ( .A1(RST), .A2(\DP/RES[12] ), .ZN(\DP/RegALU1/N15 ) );
  AND2_X1 U1966 ( .A1(RST), .A2(\DP/RES[13] ), .ZN(\DP/RegALU1/N16 ) );
  AND2_X1 U1967 ( .A1(RST), .A2(\DP/RES[14] ), .ZN(\DP/RegALU1/N17 ) );
  AND2_X1 U1968 ( .A1(RST), .A2(\DP/RES[15] ), .ZN(\DP/RegALU1/N18 ) );
  AND2_X1 U1969 ( .A1(RST), .A2(\DP/RES[16] ), .ZN(\DP/RegALU1/N19 ) );
  OR2_X1 U1970 ( .A1(w_EX_EN), .A2(n640), .ZN(\DP/RegALU1/N2 ) );
  AND2_X1 U1971 ( .A1(RST), .A2(\DP/RES[18] ), .ZN(\DP/RegALU1/N21 ) );
  AND2_X1 U1972 ( .A1(\DP/RES[20] ), .A2(RST), .ZN(\DP/RegALU1/N23 ) );
  AND2_X1 U1973 ( .A1(RST), .A2(\DP/RES[21] ), .ZN(\DP/RegALU1/N24 ) );
  AND2_X1 U1974 ( .A1(RST), .A2(\DP/RES[22] ), .ZN(\DP/RegALU1/N25 ) );
  AND2_X1 U1975 ( .A1(RST), .A2(\DP/RES[23] ), .ZN(\DP/RegALU1/N26 ) );
  AND2_X1 U1976 ( .A1(RST), .A2(\DP/RES[24] ), .ZN(\DP/RegALU1/N27 ) );
  AND2_X1 U1977 ( .A1(RST), .A2(\DP/RES[25] ), .ZN(\DP/RegALU1/N28 ) );
  AND2_X1 U1978 ( .A1(RST), .A2(\DP/RES[26] ), .ZN(\DP/RegALU1/N29 ) );
  AND2_X1 U1979 ( .A1(RST), .A2(\DP/RES[27] ), .ZN(\DP/RegALU1/N30 ) );
  AND2_X1 U1980 ( .A1(RST), .A2(\DP/RES[28] ), .ZN(\DP/RegALU1/N31 ) );
  AND2_X1 U1981 ( .A1(\DP/RES[29] ), .A2(RST), .ZN(\DP/RegALU1/N32 ) );
  AND2_X1 U1982 ( .A1(RST), .A2(\DP/RES[30] ), .ZN(\DP/RegALU1/N33 ) );
  AND2_X1 U1983 ( .A1(RST), .A2(\DP/RES[1] ), .ZN(\DP/RegALU1/N4 ) );
  AND2_X1 U1984 ( .A1(\DP/RES[2] ), .A2(RST), .ZN(\DP/RegALU1/N5 ) );
  AND2_X1 U1985 ( .A1(RST), .A2(\DP/RES[3] ), .ZN(\DP/RegALU1/N6 ) );
  AND2_X1 U1986 ( .A1(RST), .A2(\DP/RES[4] ), .ZN(\DP/RegALU1/N7 ) );
  AND2_X1 U1987 ( .A1(RST), .A2(\DP/RES[5] ), .ZN(\DP/RegALU1/N8 ) );
  AND2_X1 U1988 ( .A1(\DP/RES[6] ), .A2(RST), .ZN(\DP/RegALU1/N9 ) );
  OR2_X1 U1989 ( .A1(w_RegALU2_LATCH_EN), .A2(n641), .ZN(\DP/RegALU2/N2 ) );
  AND2_X1 U1990 ( .A1(RST), .A2(\DP/RegB_in[7] ), .ZN(\DP/RegB/N10 ) );
  AND2_X1 U1991 ( .A1(RST), .A2(\DP/RegB_in[8] ), .ZN(\DP/RegB/N11 ) );
  AND2_X1 U1992 ( .A1(RST), .A2(\DP/RegB_in[9] ), .ZN(\DP/RegB/N12 ) );
  AND2_X1 U1993 ( .A1(RST), .A2(\DP/RegB_in[10] ), .ZN(\DP/RegB/N13 ) );
  AND2_X1 U1994 ( .A1(RST), .A2(\DP/RegB_in[11] ), .ZN(\DP/RegB/N14 ) );
  AND2_X1 U1995 ( .A1(RST), .A2(\DP/RegB_in[12] ), .ZN(\DP/RegB/N15 ) );
  AND2_X1 U1996 ( .A1(RST), .A2(\DP/RegB_in[13] ), .ZN(\DP/RegB/N16 ) );
  AND2_X1 U1997 ( .A1(RST), .A2(\DP/RegB_in[14] ), .ZN(\DP/RegB/N17 ) );
  AND2_X1 U1998 ( .A1(RST), .A2(\DP/RegB_in[15] ), .ZN(\DP/RegB/N18 ) );
  AND2_X1 U1999 ( .A1(RST), .A2(\DP/RegB_in[16] ), .ZN(\DP/RegB/N19 ) );
  OR2_X1 U2000 ( .A1(n641), .A2(w_RF_RD2), .ZN(\DP/RegB/N2 ) );
  AND2_X1 U2001 ( .A1(RST), .A2(\DP/RegB_in[17] ), .ZN(\DP/RegB/N20 ) );
  AND2_X1 U2002 ( .A1(RST), .A2(\DP/RegB_in[18] ), .ZN(\DP/RegB/N21 ) );
  AND2_X1 U2003 ( .A1(RST), .A2(\DP/RegB_in[19] ), .ZN(\DP/RegB/N22 ) );
  AND2_X1 U2004 ( .A1(RST), .A2(\DP/RegB_in[20] ), .ZN(\DP/RegB/N23 ) );
  AND2_X1 U2005 ( .A1(RST), .A2(\DP/RegB_in[21] ), .ZN(\DP/RegB/N24 ) );
  AND2_X1 U2006 ( .A1(RST), .A2(\DP/RegB_in[22] ), .ZN(\DP/RegB/N25 ) );
  AND2_X1 U2007 ( .A1(RST), .A2(\DP/RegB_in[23] ), .ZN(\DP/RegB/N26 ) );
  AND2_X1 U2008 ( .A1(RST), .A2(\DP/RegB_in[24] ), .ZN(\DP/RegB/N27 ) );
  AND2_X1 U2009 ( .A1(RST), .A2(\DP/RegB_in[25] ), .ZN(\DP/RegB/N28 ) );
  AND2_X1 U2010 ( .A1(RST), .A2(\DP/RegB_in[26] ), .ZN(\DP/RegB/N29 ) );
  AND2_X1 U2011 ( .A1(RST), .A2(\DP/RegB_in[0] ), .ZN(\DP/RegB/N3 ) );
  AND2_X1 U2012 ( .A1(RST), .A2(\DP/RegB_in[27] ), .ZN(\DP/RegB/N30 ) );
  AND2_X1 U2013 ( .A1(RST), .A2(\DP/RegB_in[28] ), .ZN(\DP/RegB/N31 ) );
  AND2_X1 U2014 ( .A1(RST), .A2(\DP/RegB_in[29] ), .ZN(\DP/RegB/N32 ) );
  AND2_X1 U2015 ( .A1(RST), .A2(\DP/RegB_in[30] ), .ZN(\DP/RegB/N33 ) );
  AND2_X1 U2016 ( .A1(RST), .A2(\DP/RegB_in[31] ), .ZN(\DP/RegB/N34 ) );
  AND2_X1 U2017 ( .A1(RST), .A2(\DP/RegB_in[1] ), .ZN(\DP/RegB/N4 ) );
  AND2_X1 U2018 ( .A1(RST), .A2(\DP/RegB_in[2] ), .ZN(\DP/RegB/N5 ) );
  AND2_X1 U2019 ( .A1(RST), .A2(\DP/RegB_in[3] ), .ZN(\DP/RegB/N6 ) );
  AND2_X1 U2020 ( .A1(RST), .A2(\DP/RegB_in[4] ), .ZN(\DP/RegB/N7 ) );
  AND2_X1 U2021 ( .A1(RST), .A2(\DP/RegB_in[5] ), .ZN(\DP/RegB/N8 ) );
  AND2_X1 U2022 ( .A1(RST), .A2(\DP/RegB_in[6] ), .ZN(\DP/RegB/N9 ) );
  NAND2_X1 U2023 ( .A1(n1544), .A2(IR_OUT[24]), .ZN(n1049) );
  NAND2_X1 U2024 ( .A1(n1544), .A2(IR_OUT[21]), .ZN(n1047) );
  NAND2_X1 U2025 ( .A1(n1544), .A2(IR_OUT[22]), .ZN(n1048) );
  NAND2_X1 U2026 ( .A1(n1544), .A2(IR_OUT[25]), .ZN(n1051) );
  OR4_X1 U2027 ( .A1(\DP/RD1[1] ), .A2(\DP/RD1[0] ), .A3(\DP/RD1[4] ), .A4(
        \DP/RD1[3] ), .ZN(n1012) );
  OAI21_X1 U2028 ( .B1(\DP/RD1[2] ), .B2(n1012), .A(w_RF_WE_EX), .ZN(n1033) );
  OAI22_X1 U2029 ( .A1(n1047), .A2(\DP/RD1[0] ), .B1(n1049), .B2(\DP/RD1[3] ), 
        .ZN(n1013) );
  AOI221_X1 U2030 ( .B1(n1047), .B2(\DP/RD1[0] ), .C1(\DP/RD1[3] ), .C2(n1049), 
        .A(n1013), .ZN(n1018) );
  NAND2_X1 U2031 ( .A1(n1544), .A2(IR_OUT[23]), .ZN(n1280) );
  AOI22_X1 U2032 ( .A1(n1280), .A2(\DP/RD1[2] ), .B1(n1048), .B2(\DP/RD1[1] ), 
        .ZN(n1015) );
  NOR2_X1 U2036 ( .A1(n1033), .A2(n1019), .ZN(n1028) );
  OAI221_X1 U2038 ( .B1(n41), .B2(n72), .C1(n1049), .C2(n584), .A(n1020), .ZN(
        n1025) );
  AOI22_X1 U2039 ( .A1(n42), .A2(n73), .B1(n1048), .B2(\DP/RD2[1] ), .ZN(n1021) );
  OAI221_X1 U2040 ( .B1(n42), .B2(n73), .C1(n1822), .C2(\DP/RD2[1] ), .A(n1021), .ZN(n1024) );
  AOI22_X1 U2041 ( .A1(n1280), .A2(\DP/RD2[2] ), .B1(n1047), .B2(\DP/RD2[0] ), 
        .ZN(n1022) );
  OAI221_X1 U2042 ( .B1(n1280), .B2(\DP/RD2[2] ), .C1(n1047), .C2(\DP/RD2[0] ), 
        .A(n1022), .ZN(n1023) );
  NOR3_X1 U2044 ( .A1(n1027), .A2(n1028), .A3(n640), .ZN(\DP/RegFC/N3 ) );
  AND2_X1 U2045 ( .A1(RST), .A2(n1027), .ZN(\DP/RegFC/N4 ) );
  AND2_X1 U2046 ( .A1(RST), .A2(n1028), .ZN(\DP/RegFC/N5 ) );
  OAI22_X1 U2047 ( .A1(n1203), .A2(\DP/RD1[0] ), .B1(n1206), .B2(\DP/RD1[3] ), 
        .ZN(n1029) );
  AOI221_X1 U2048 ( .B1(n1203), .B2(\DP/RD1[0] ), .C1(\DP/RD1[3] ), .C2(n1206), 
        .A(n1029), .ZN(n1030) );
  OAI221_X1 U2049 ( .B1(n32), .B2(n597), .C1(n1205), .C2(\DP/RD1[2] ), .A(
        n1030), .ZN(n1031) );
  NOR2_X1 U2052 ( .A1(n1034), .A2(n1033), .ZN(n1038) );
  INV_X1 U2053 ( .A(n1034), .ZN(n1036) );
  NOR2_X1 U2054 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR3_X1 U2055 ( .A1(n1037), .A2(n1038), .A3(n640), .ZN(\DP/RegFB/N3 ) );
  AND2_X1 U2058 ( .A1(IR_OUT[7]), .A2(n1056), .ZN(\DP/RegIMM/N10 ) );
  AND2_X1 U2059 ( .A1(IR_OUT[8]), .A2(n1056), .ZN(\DP/RegIMM/N11 ) );
  INV_X1 U2060 ( .A(n1056), .ZN(n1055) );
  NOR2_X1 U2061 ( .A1(n600), .A2(n1055), .ZN(\DP/RegIMM/N12 ) );
  AND2_X1 U2062 ( .A1(IR_OUT[10]), .A2(n1056), .ZN(\DP/RegIMM/N13 ) );
  NAND2_X1 U2063 ( .A1(n1056), .A2(IR_OUT[11]), .ZN(n190) );
  NAND2_X1 U2064 ( .A1(n1056), .A2(IR_OUT[12]), .ZN(n188) );
  NAND2_X1 U2065 ( .A1(n1056), .A2(IR_OUT[13]), .ZN(n186) );
  NAND2_X1 U2066 ( .A1(n1056), .A2(IR_OUT[14]), .ZN(n184) );
  NAND2_X1 U2067 ( .A1(n1056), .A2(IR_OUT[15]), .ZN(n181) );
  OAI211_X1 U2068 ( .C1(n586), .C2(n592), .A(n1823), .B(n1581), .ZN(n1044) );
  NAND4_X1 U2069 ( .A1(n1043), .A2(n1044), .A3(n1201), .A4(n1368), .ZN(n1045)
         );
  OAI21_X1 U2071 ( .B1(n1203), .B2(n1052), .A(n1050), .ZN(\DP/RegIMM/N19 ) );
  NAND2_X1 U2072 ( .A1(n1046), .A2(RST), .ZN(\DP/RegIMM/N2 ) );
  OAI21_X1 U2073 ( .B1(n1052), .B2(n1452), .A(n1050), .ZN(\DP/RegIMM/N20 ) );
  OAI21_X1 U2074 ( .B1(n1052), .B2(n1205), .A(n1050), .ZN(\DP/RegIMM/N21 ) );
  OAI21_X1 U2075 ( .B1(n1052), .B2(n1206), .A(n1050), .ZN(\DP/RegIMM/N22 ) );
  OAI21_X1 U2076 ( .B1(n1052), .B2(n1301), .A(n1050), .ZN(\DP/RegIMM/N23 ) );
  OAI21_X1 U2077 ( .B1(n1052), .B2(n1047), .A(n1050), .ZN(\DP/RegIMM/N24 ) );
  OAI21_X1 U2078 ( .B1(n1052), .B2(n1822), .A(n1050), .ZN(\DP/RegIMM/N25 ) );
  OAI21_X1 U2079 ( .B1(n1052), .B2(n1280), .A(n1050), .ZN(\DP/RegIMM/N26 ) );
  OAI21_X1 U2080 ( .B1(n1052), .B2(n1049), .A(n1050), .ZN(\DP/RegIMM/N27 ) );
  OAI21_X1 U2081 ( .B1(n1052), .B2(n1051), .A(n1050), .ZN(\DP/RegIMM/N34 ) );
  NOR2_X1 U2082 ( .A1(n640), .A2(n1053), .ZN(\DP/RegIMM/N5 ) );
  NOR2_X1 U2083 ( .A1(n641), .A2(n1472), .ZN(\DP/RegIMM/N6 ) );
  NOR2_X1 U2084 ( .A1(n595), .A2(n1055), .ZN(\DP/RegIMM/N7 ) );
  AND2_X1 U2085 ( .A1(IR_OUT[6]), .A2(n1056), .ZN(\DP/RegIMM/N9 ) );
  NAND4_X1 U2086 ( .A1(n53), .A2(RST), .A3(w_LOAD_SIZE[2]), .A4(n587), .ZN(
        n1057) );
  NOR3_X1 U2087 ( .A1(w_LOAD_SIZE[2]), .A2(n602), .A3(n587), .ZN(n1069) );
  NOR3_X1 U2088 ( .A1(n53), .A2(w_LOAD_SIZE[2]), .A3(w_LOAD_SIZE[1]), .ZN(
        n1068) );
  NAND2_X1 U2089 ( .A1(n1057), .A2(n1067), .ZN(n1090) );
  AND2_X1 U2090 ( .A1(\DP/LOAD8[7] ), .A2(n1090), .ZN(\DP/RegLMD/N10 ) );
  INV_X1 U2091 ( .A(\DP/LOAD16[8] ), .ZN(n1059) );
  INV_X1 U2092 ( .A(n1057), .ZN(n1058) );
  OAI21_X1 U2093 ( .B1(n1067), .B2(n1059), .A(n1071), .ZN(\DP/RegLMD/N11 ) );
  INV_X1 U2094 ( .A(\DP/LOAD16[9] ), .ZN(n1060) );
  OAI21_X1 U2095 ( .B1(n1067), .B2(n1060), .A(n1071), .ZN(\DP/RegLMD/N12 ) );
  INV_X1 U2096 ( .A(\DP/LOAD16[10] ), .ZN(n1061) );
  OAI21_X1 U2097 ( .B1(n1067), .B2(n1061), .A(n1071), .ZN(\DP/RegLMD/N13 ) );
  INV_X1 U2098 ( .A(\DP/LOAD16[11] ), .ZN(n1062) );
  OAI21_X1 U2099 ( .B1(n1067), .B2(n1062), .A(n1071), .ZN(\DP/RegLMD/N14 ) );
  INV_X1 U2100 ( .A(\DP/LOAD16[12] ), .ZN(n1063) );
  OAI21_X1 U2101 ( .B1(n1067), .B2(n1063), .A(n1071), .ZN(\DP/RegLMD/N15 ) );
  INV_X1 U2102 ( .A(\DP/LOAD16[13] ), .ZN(n1064) );
  OAI21_X1 U2103 ( .B1(n1067), .B2(n1064), .A(n1071), .ZN(\DP/RegLMD/N16 ) );
  INV_X1 U2104 ( .A(\DP/LOAD16[14] ), .ZN(n1065) );
  OAI21_X1 U2105 ( .B1(n1067), .B2(n1065), .A(n1071), .ZN(\DP/RegLMD/N17 ) );
  INV_X1 U2106 ( .A(\DP/LOAD16[15] ), .ZN(n1066) );
  OAI21_X1 U2107 ( .B1(n1067), .B2(n1066), .A(n1071), .ZN(\DP/RegLMD/N18 ) );
  NAND4_X1 U2108 ( .A1(RST), .A2(n1069), .A3(w_SIGN_LD), .A4(\DP/LOAD16[15] ), 
        .ZN(n1070) );
  AOI21_X1 U2109 ( .B1(n1088), .B2(DRAM_DATA_IN[16]), .A(n1087), .ZN(n1072) );
  INV_X1 U2110 ( .A(n1072), .ZN(\DP/RegLMD/N19 ) );
  OR2_X1 U2111 ( .A1(w_RegLMD_LATCH_EN), .A2(n640), .ZN(\DP/RegLMD/N2 ) );
  AOI21_X1 U2112 ( .B1(n1088), .B2(DRAM_DATA_IN[17]), .A(n1087), .ZN(n1073) );
  INV_X1 U2113 ( .A(n1073), .ZN(\DP/RegLMD/N20 ) );
  AOI21_X1 U2114 ( .B1(n1088), .B2(DRAM_DATA_IN[18]), .A(n1087), .ZN(n1074) );
  INV_X1 U2115 ( .A(n1074), .ZN(\DP/RegLMD/N21 ) );
  AOI21_X1 U2116 ( .B1(n1088), .B2(DRAM_DATA_IN[19]), .A(n1087), .ZN(n1075) );
  INV_X1 U2117 ( .A(n1075), .ZN(\DP/RegLMD/N22 ) );
  AOI21_X1 U2118 ( .B1(n1088), .B2(DRAM_DATA_IN[20]), .A(n1087), .ZN(n1076) );
  INV_X1 U2119 ( .A(n1076), .ZN(\DP/RegLMD/N23 ) );
  AOI21_X1 U2120 ( .B1(n1088), .B2(DRAM_DATA_IN[21]), .A(n1087), .ZN(n1077) );
  AOI21_X1 U2122 ( .B1(n1088), .B2(DRAM_DATA_IN[22]), .A(n1087), .ZN(n1078) );
  INV_X1 U2123 ( .A(n1078), .ZN(\DP/RegLMD/N25 ) );
  AOI21_X1 U2124 ( .B1(n1088), .B2(DRAM_DATA_IN[23]), .A(n1087), .ZN(n1079) );
  INV_X1 U2125 ( .A(n1079), .ZN(\DP/RegLMD/N26 ) );
  AOI21_X1 U2126 ( .B1(n1088), .B2(DRAM_DATA_IN[24]), .A(n1087), .ZN(n1080) );
  INV_X1 U2127 ( .A(n1080), .ZN(\DP/RegLMD/N27 ) );
  AOI21_X1 U2128 ( .B1(n1088), .B2(DRAM_DATA_IN[25]), .A(n1087), .ZN(n1081) );
  INV_X1 U2129 ( .A(n1081), .ZN(\DP/RegLMD/N28 ) );
  AOI21_X1 U2130 ( .B1(n1088), .B2(DRAM_DATA_IN[26]), .A(n1087), .ZN(n1082) );
  INV_X1 U2131 ( .A(n1082), .ZN(\DP/RegLMD/N29 ) );
  AND2_X1 U2132 ( .A1(\DP/LOAD8[0] ), .A2(n1090), .ZN(\DP/RegLMD/N3 ) );
  AOI21_X1 U2133 ( .B1(n1088), .B2(DRAM_DATA_IN[27]), .A(n1087), .ZN(n1083) );
  INV_X1 U2134 ( .A(n1083), .ZN(\DP/RegLMD/N30 ) );
  AOI21_X1 U2135 ( .B1(n1088), .B2(DRAM_DATA_IN[28]), .A(n1087), .ZN(n1084) );
  INV_X1 U2136 ( .A(n1084), .ZN(\DP/RegLMD/N31 ) );
  AOI21_X1 U2137 ( .B1(n1088), .B2(DRAM_DATA_IN[29]), .A(n1087), .ZN(n1085) );
  INV_X1 U2138 ( .A(n1085), .ZN(\DP/RegLMD/N32 ) );
  AOI21_X1 U2139 ( .B1(n1088), .B2(DRAM_DATA_IN[30]), .A(n1087), .ZN(n1086) );
  INV_X1 U2140 ( .A(n1086), .ZN(\DP/RegLMD/N33 ) );
  AOI21_X1 U2141 ( .B1(n1088), .B2(DRAM_DATA_IN[31]), .A(n1087), .ZN(n1089) );
  INV_X1 U2142 ( .A(n1089), .ZN(\DP/RegLMD/N34 ) );
  AND2_X1 U2143 ( .A1(\DP/LOAD8[1] ), .A2(n1090), .ZN(\DP/RegLMD/N4 ) );
  AND2_X1 U2144 ( .A1(\DP/LOAD8[2] ), .A2(n1090), .ZN(\DP/RegLMD/N5 ) );
  AND2_X1 U2145 ( .A1(\DP/LOAD8[3] ), .A2(n1090), .ZN(\DP/RegLMD/N6 ) );
  AND2_X1 U2146 ( .A1(\DP/LOAD8[4] ), .A2(n1090), .ZN(\DP/RegLMD/N7 ) );
  AND2_X1 U2147 ( .A1(\DP/LOAD8[5] ), .A2(n1090), .ZN(\DP/RegLMD/N8 ) );
  AND2_X1 U2148 ( .A1(\DP/LOAD8[6] ), .A2(n1090), .ZN(\DP/RegLMD/N9 ) );
  AND2_X1 U2149 ( .A1(RST), .A2(\DP/RegB_out[7] ), .ZN(\DP/RegME/N10 ) );
  AND2_X1 U2150 ( .A1(RST), .A2(\DP/RegB_out[8] ), .ZN(\DP/RegME/N11 ) );
  AND2_X1 U2151 ( .A1(RST), .A2(\DP/RegB_out[9] ), .ZN(\DP/RegME/N12 ) );
  AND2_X1 U2152 ( .A1(RST), .A2(\DP/RegB_out[10] ), .ZN(\DP/RegME/N13 ) );
  AND2_X1 U2153 ( .A1(RST), .A2(\DP/RegB_out[11] ), .ZN(\DP/RegME/N14 ) );
  AND2_X1 U2154 ( .A1(RST), .A2(\DP/RegB_out[12] ), .ZN(\DP/RegME/N15 ) );
  AND2_X1 U2155 ( .A1(RST), .A2(\DP/RegB_out[13] ), .ZN(\DP/RegME/N16 ) );
  AND2_X1 U2156 ( .A1(RST), .A2(\DP/RegB_out[14] ), .ZN(\DP/RegME/N17 ) );
  AND2_X1 U2157 ( .A1(RST), .A2(\DP/RegB_out[15] ), .ZN(\DP/RegME/N18 ) );
  AND2_X1 U2158 ( .A1(RST), .A2(\DP/RegB_out[16] ), .ZN(\DP/RegME/N19 ) );
  OR2_X1 U2159 ( .A1(w_RegME_LATCH_EN), .A2(n640), .ZN(\DP/RegME/N2 ) );
  AND2_X1 U2160 ( .A1(RST), .A2(\DP/RegB_out[17] ), .ZN(\DP/RegME/N20 ) );
  AND2_X1 U2161 ( .A1(RST), .A2(\DP/RegB_out[18] ), .ZN(\DP/RegME/N21 ) );
  AND2_X1 U2162 ( .A1(RST), .A2(\DP/RegB_out[19] ), .ZN(\DP/RegME/N22 ) );
  AND2_X1 U2163 ( .A1(RST), .A2(\DP/RegB_out[20] ), .ZN(\DP/RegME/N23 ) );
  AND2_X1 U2164 ( .A1(RST), .A2(\DP/RegB_out[21] ), .ZN(\DP/RegME/N24 ) );
  AND2_X1 U2165 ( .A1(RST), .A2(\DP/RegB_out[22] ), .ZN(\DP/RegME/N25 ) );
  AND2_X1 U2166 ( .A1(RST), .A2(\DP/RegB_out[23] ), .ZN(\DP/RegME/N26 ) );
  AND2_X1 U2167 ( .A1(RST), .A2(\DP/RegB_out[24] ), .ZN(\DP/RegME/N27 ) );
  AND2_X1 U2168 ( .A1(RST), .A2(\DP/RegB_out[25] ), .ZN(\DP/RegME/N28 ) );
  AND2_X1 U2169 ( .A1(RST), .A2(\DP/RegB_out[26] ), .ZN(\DP/RegME/N29 ) );
  AND2_X1 U2170 ( .A1(RST), .A2(\DP/RegB_out[0] ), .ZN(\DP/RegME/N3 ) );
  AND2_X1 U2171 ( .A1(RST), .A2(\DP/RegB_out[27] ), .ZN(\DP/RegME/N30 ) );
  AND2_X1 U2172 ( .A1(RST), .A2(\DP/RegB_out[28] ), .ZN(\DP/RegME/N31 ) );
  AND2_X1 U2173 ( .A1(RST), .A2(\DP/RegB_out[29] ), .ZN(\DP/RegME/N32 ) );
  AND2_X1 U2174 ( .A1(RST), .A2(\DP/RegB_out[30] ), .ZN(\DP/RegME/N33 ) );
  AND2_X1 U2175 ( .A1(RST), .A2(\DP/RegB_out[31] ), .ZN(\DP/RegME/N34 ) );
  AND2_X1 U2176 ( .A1(RST), .A2(\DP/RegB_out[1] ), .ZN(\DP/RegME/N4 ) );
  AND2_X1 U2177 ( .A1(RST), .A2(\DP/RegB_out[2] ), .ZN(\DP/RegME/N5 ) );
  AND2_X1 U2178 ( .A1(RST), .A2(\DP/RegB_out[3] ), .ZN(\DP/RegME/N6 ) );
  AND2_X1 U2179 ( .A1(RST), .A2(\DP/RegB_out[4] ), .ZN(\DP/RegME/N7 ) );
  AND2_X1 U2180 ( .A1(RST), .A2(\DP/RegB_out[5] ), .ZN(\DP/RegME/N8 ) );
  AND2_X1 U2181 ( .A1(RST), .A2(\DP/RegB_out[6] ), .ZN(\DP/RegME/N9 ) );
  OAI21_X1 U2188 ( .B1(n1091), .B2(IROM_ADDR[7]), .A(n633), .ZN(n1093) );
  AOI22_X1 U2189 ( .A1(n632), .A2(\DP/RegALU2/N10 ), .B1(n631), .B2(
        \DP/RegA1_out[7] ), .ZN(n1092) );
  OAI21_X1 U2190 ( .B1(n1094), .B2(n1093), .A(n1092), .ZN(\PC/N10 ) );
  AOI22_X1 U2191 ( .A1(n1196), .A2(\DP/RegALU2/N11 ), .B1(n1195), .B2(
        \DP/RegA1_out[8] ), .ZN(n1096) );
  OAI211_X1 U2193 ( .C1(n1094), .C2(IROM_ADDR[8]), .A(n634), .B(n1097), .ZN(
        n1095) );
  NAND2_X1 U2194 ( .A1(n1096), .A2(n1095), .ZN(\PC/N11 ) );
  OAI21_X1 U2196 ( .B1(n1098), .B2(IROM_ADDR[9]), .A(n633), .ZN(n1100) );
  AOI22_X1 U2197 ( .A1(n632), .A2(\DP/RegALU2/N12 ), .B1(n631), .B2(
        \DP/RegA1_out[9] ), .ZN(n1099) );
  OAI21_X1 U2198 ( .B1(n1101), .B2(n1100), .A(n1099), .ZN(\PC/N12 ) );
  AOI22_X1 U2199 ( .A1(n1196), .A2(\DP/RegALU2/N13 ), .B1(n1195), .B2(
        \DP/RegA1_out[10] ), .ZN(n1103) );
  OAI211_X1 U2201 ( .C1(n1101), .C2(IROM_ADDR[10]), .A(n634), .B(n1104), .ZN(
        n1102) );
  NAND2_X1 U2202 ( .A1(n1103), .A2(n1102), .ZN(\PC/N13 ) );
  OAI21_X1 U2204 ( .B1(n1105), .B2(IROM_ADDR[11]), .A(n633), .ZN(n1107) );
  AOI22_X1 U2205 ( .A1(n632), .A2(\DP/RegALU2/N14 ), .B1(n631), .B2(
        \DP/RegA1_out[11] ), .ZN(n1106) );
  OAI21_X1 U2206 ( .B1(n1108), .B2(n1107), .A(n1106), .ZN(\PC/N14 ) );
  AOI22_X1 U2207 ( .A1(n1196), .A2(\DP/RegALU2/N15 ), .B1(n1195), .B2(
        \DP/RegA1_out[12] ), .ZN(n1110) );
  OAI211_X1 U2209 ( .C1(n1108), .C2(w_PC_OUT[12]), .A(n633), .B(n1111), .ZN(
        n1109) );
  NAND2_X1 U2210 ( .A1(n1110), .A2(n1109), .ZN(\PC/N15 ) );
  OAI21_X1 U2212 ( .B1(n1112), .B2(\DP/NPC1[13] ), .A(n634), .ZN(n1114) );
  AOI22_X1 U2213 ( .A1(n1196), .A2(\DP/RegALU2/N16 ), .B1(n1195), .B2(
        \DP/RegA1_out[13] ), .ZN(n1113) );
  OAI21_X1 U2214 ( .B1(n1115), .B2(n1114), .A(n1113), .ZN(\PC/N16 ) );
  AOI22_X1 U2215 ( .A1(n1196), .A2(\DP/RegALU2/N17 ), .B1(n1195), .B2(
        \DP/RegA1_out[14] ), .ZN(n1117) );
  OAI211_X1 U2217 ( .C1(n1115), .C2(\DP/NPC1[14] ), .A(n633), .B(n1323), .ZN(
        n1116) );
  NAND2_X1 U2218 ( .A1(n1117), .A2(n1116), .ZN(\PC/N17 ) );
  OAI21_X1 U2220 ( .B1(n1119), .B2(\DP/NPC1[15] ), .A(n634), .ZN(n1121) );
  AOI22_X1 U2221 ( .A1(n1196), .A2(\DP/RegALU2/N18 ), .B1(n1195), .B2(
        \DP/RegA1_out[15] ), .ZN(n1120) );
  OAI21_X1 U2222 ( .B1(n1324), .B2(n1121), .A(n1120), .ZN(\PC/N18 ) );
  AOI22_X1 U2223 ( .A1(n1196), .A2(\DP/RegALU2/N19 ), .B1(n1195), .B2(
        \DP/RegA1_out[16] ), .ZN(n1124) );
  OAI211_X1 U2225 ( .C1(n1324), .C2(\DP/NPC1[16] ), .A(n633), .B(n1125), .ZN(
        n1123) );
  NAND2_X1 U2226 ( .A1(n1124), .A2(n1123), .ZN(\PC/N19 ) );
  OR2_X1 U2227 ( .A1(w_IF_EN), .A2(n641), .ZN(\PC/N2 ) );
  OAI21_X1 U2229 ( .B1(n1126), .B2(w_PC_OUT[17]), .A(n634), .ZN(n1128) );
  AOI22_X1 U2230 ( .A1(n1196), .A2(\DP/RegALU2/N20 ), .B1(n1195), .B2(
        \DP/RegA1_out[17] ), .ZN(n1127) );
  OAI21_X1 U2231 ( .B1(n1129), .B2(n1128), .A(n1127), .ZN(\PC/N20 ) );
  AOI22_X1 U2232 ( .A1(n1196), .A2(\DP/RegALU2/N21 ), .B1(n1195), .B2(
        \DP/RegA1_out[18] ), .ZN(n1131) );
  OAI211_X1 U2234 ( .C1(n1129), .C2(w_PC_OUT[18]), .A(n633), .B(n1132), .ZN(
        n1130) );
  NAND2_X1 U2235 ( .A1(n1131), .A2(n1130), .ZN(\PC/N21 ) );
  OAI21_X1 U2237 ( .B1(n1133), .B2(\DP/NPC1[19] ), .A(n634), .ZN(n1135) );
  AOI22_X1 U2238 ( .A1(n632), .A2(\DP/RegALU2/N22 ), .B1(n1195), .B2(
        \DP/RegA1_out[19] ), .ZN(n1134) );
  OAI21_X1 U2239 ( .B1(n1136), .B2(n1135), .A(n1134), .ZN(\PC/N22 ) );
  AOI22_X1 U2240 ( .A1(n632), .A2(\DP/RegALU2/N23 ), .B1(n631), .B2(
        \DP/RegA1_out[20] ), .ZN(n1138) );
  OAI211_X1 U2242 ( .C1(n1136), .C2(\DP/NPC1[20] ), .A(n633), .B(n1139), .ZN(
        n1137) );
  NAND2_X1 U2243 ( .A1(n1138), .A2(n1137), .ZN(\PC/N23 ) );
  OAI21_X1 U2245 ( .B1(n1140), .B2(w_PC_OUT[21]), .A(n634), .ZN(n1142) );
  AOI22_X1 U2246 ( .A1(n632), .A2(\DP/RegALU2/N24 ), .B1(n1195), .B2(
        \DP/RegA1_out[21] ), .ZN(n1141) );
  OAI21_X1 U2247 ( .B1(n1143), .B2(n1142), .A(n1141), .ZN(\PC/N24 ) );
  AOI22_X1 U2248 ( .A1(n632), .A2(\DP/RegALU2/N25 ), .B1(n631), .B2(
        \DP/RegA1_out[22] ), .ZN(n1145) );
  OAI211_X1 U2250 ( .C1(n1143), .C2(\DP/NPC1[22] ), .A(n633), .B(n1146), .ZN(
        n1144) );
  NAND2_X1 U2251 ( .A1(n1145), .A2(n1144), .ZN(\PC/N25 ) );
  OAI21_X1 U2253 ( .B1(n1359), .B2(\DP/NPC1[23] ), .A(n634), .ZN(n1149) );
  AOI22_X1 U2254 ( .A1(n632), .A2(\DP/RegALU2/N26 ), .B1(n1195), .B2(
        \DP/RegA1_out[23] ), .ZN(n1148) );
  OAI21_X1 U2255 ( .B1(n1150), .B2(n1149), .A(n1148), .ZN(\PC/N26 ) );
  AOI22_X1 U2256 ( .A1(n632), .A2(\DP/RegALU2/N27 ), .B1(n631), .B2(
        \DP/RegA1_out[24] ), .ZN(n1152) );
  OAI211_X1 U2258 ( .C1(n1150), .C2(w_PC_OUT[24]), .A(n633), .B(n1153), .ZN(
        n1151) );
  NAND2_X1 U2259 ( .A1(n1152), .A2(n1151), .ZN(\PC/N27 ) );
  OAI21_X1 U2261 ( .B1(n1154), .B2(w_PC_OUT[25]), .A(n633), .ZN(n1156) );
  AOI22_X1 U2262 ( .A1(n632), .A2(\DP/RegALU2/N28 ), .B1(n1195), .B2(
        \DP/RegA1_out[25] ), .ZN(n1155) );
  OAI21_X1 U2263 ( .B1(n1156), .B2(n1157), .A(n1155), .ZN(\PC/N28 ) );
  AOI22_X1 U2264 ( .A1(n632), .A2(\DP/RegALU2/N29 ), .B1(n631), .B2(
        \DP/RegA1_out[26] ), .ZN(n1159) );
  NAND2_X1 U2267 ( .A1(n1158), .A2(n1159), .ZN(\PC/N29 ) );
  AOI22_X1 U2268 ( .A1(n632), .A2(\DP/RegALU2/N3 ), .B1(n1195), .B2(
        \DP/RegA1_out[0] ), .ZN(n1160) );
  OAI21_X1 U2269 ( .B1(IROM_ADDR[0]), .B2(n591), .A(n1160), .ZN(\PC/N3 ) );
  AOI22_X1 U2272 ( .A1(n632), .A2(\DP/RegALU2/N30 ), .B1(n631), .B2(
        \DP/RegA1_out[27] ), .ZN(n1163) );
  OAI21_X1 U2273 ( .B1(n1165), .B2(n1164), .A(n1163), .ZN(\PC/N30 ) );
  AOI22_X1 U2274 ( .A1(n1196), .A2(\DP/RegALU2/N31 ), .B1(n1195), .B2(
        \DP/RegA1_out[28] ), .ZN(n1167) );
  AOI22_X1 U2280 ( .A1(n1196), .A2(\DP/RegALU2/N32 ), .B1(n1195), .B2(
        \DP/RegA1_out[29] ), .ZN(n1170) );
  OAI21_X1 U2281 ( .B1(n1172), .B2(n1171), .A(n1170), .ZN(\PC/N32 ) );
  AOI22_X1 U2284 ( .A1(n632), .A2(\DP/RegALU2/N33 ), .B1(n631), .B2(
        \DP/RegA1_out[30] ), .ZN(n1173) );
  AOI22_X1 U2287 ( .A1(n632), .A2(\DP/RegALU2/N34 ), .B1(n631), .B2(
        \DP/RegA1_out[31] ), .ZN(n1176) );
  OAI21_X1 U2288 ( .B1(n1177), .B2(n591), .A(n1176), .ZN(\PC/N34 ) );
  AOI22_X1 U2289 ( .A1(n632), .A2(\DP/RegALU2/N4 ), .B1(n631), .B2(
        \DP/RegA1_out[1] ), .ZN(n1179) );
  NAND2_X1 U2290 ( .A1(IROM_ADDR[0]), .A2(\DP/NPC1[1] ), .ZN(n1180) );
  OAI211_X1 U2291 ( .C1(IROM_ADDR[0]), .C2(\DP/NPC1[1] ), .A(n634), .B(n1180), 
        .ZN(n1178) );
  NAND2_X1 U2292 ( .A1(n1179), .A2(n1178), .ZN(\PC/N4 ) );
  AOI22_X1 U2293 ( .A1(n632), .A2(\DP/RegALU2/N5 ), .B1(n631), .B2(
        \DP/RegA1_out[2] ), .ZN(n1184) );
  INV_X1 U2294 ( .A(n1180), .ZN(n1182) );
  OAI211_X1 U2295 ( .C1(n1182), .C2(\DP/NPC1[2] ), .A(n634), .B(n1181), .ZN(
        n1183) );
  NAND2_X1 U2296 ( .A1(n1184), .A2(n1183), .ZN(\PC/N5 ) );
  OAI21_X1 U2297 ( .B1(n1185), .B2(\DP/NPC1[3] ), .A(n633), .ZN(n1187) );
  AOI22_X1 U2298 ( .A1(n632), .A2(\DP/RegALU2/N6 ), .B1(n631), .B2(
        \DP/RegA1_out[3] ), .ZN(n1186) );
  OAI21_X1 U2299 ( .B1(n1189), .B2(n1187), .A(n1186), .ZN(\PC/N6 ) );
  AOI22_X1 U2300 ( .A1(n632), .A2(\DP/RegALU2/N7 ), .B1(n631), .B2(
        \DP/RegA1_out[4] ), .ZN(n1191) );
  OAI211_X1 U2301 ( .C1(n1189), .C2(\DP/NPC1[4] ), .A(n634), .B(n1188), .ZN(
        n1190) );
  NAND2_X1 U2302 ( .A1(n1191), .A2(n1190), .ZN(\PC/N7 ) );
  OAI21_X1 U2303 ( .B1(n1192), .B2(IROM_ADDR[5]), .A(n634), .ZN(n1194) );
  AOI22_X1 U2304 ( .A1(n632), .A2(\DP/RegALU2/N8 ), .B1(n631), .B2(
        \DP/RegA1_out[5] ), .ZN(n1193) );
  OAI21_X1 U2305 ( .B1(n1198), .B2(n1194), .A(n1193), .ZN(\PC/N8 ) );
  AOI22_X1 U2306 ( .A1(n632), .A2(\DP/RegALU2/N9 ), .B1(n631), .B2(
        \DP/RegA1_out[6] ), .ZN(n1200) );
  OAI211_X1 U2307 ( .C1(n1198), .C2(\DP/NPC1[6] ), .A(n633), .B(n1197), .ZN(
        n1199) );
  NAND2_X1 U2308 ( .A1(n1200), .A2(n1199), .ZN(\PC/N9 ) );
  AND2_X1 U2309 ( .A1(RST), .A2(\DP/NPC1[7] ), .ZN(\DP/RegNPC1/N10 ) );
  AND2_X1 U2310 ( .A1(RST), .A2(\DP/NPC1[8] ), .ZN(\DP/RegNPC1/N11 ) );
  AND2_X1 U2311 ( .A1(RST), .A2(\DP/NPC1[9] ), .ZN(\DP/RegNPC1/N12 ) );
  AND2_X1 U2312 ( .A1(RST), .A2(\DP/NPC1[10] ), .ZN(\DP/RegNPC1/N13 ) );
  AND2_X1 U2313 ( .A1(RST), .A2(\DP/NPC1[11] ), .ZN(\DP/RegNPC1/N14 ) );
  AND2_X1 U2314 ( .A1(RST), .A2(\DP/NPC1[12] ), .ZN(\DP/RegNPC1/N15 ) );
  AND2_X1 U2315 ( .A1(RST), .A2(\DP/NPC1[13] ), .ZN(\DP/RegNPC1/N16 ) );
  AND2_X1 U2316 ( .A1(RST), .A2(\DP/NPC1[14] ), .ZN(\DP/RegNPC1/N17 ) );
  AND2_X1 U2317 ( .A1(RST), .A2(\DP/NPC1[15] ), .ZN(\DP/RegNPC1/N18 ) );
  AND2_X1 U2318 ( .A1(RST), .A2(\DP/NPC1[16] ), .ZN(\DP/RegNPC1/N19 ) );
  AND2_X1 U2319 ( .A1(RST), .A2(\DP/NPC1[17] ), .ZN(\DP/RegNPC1/N20 ) );
  AND2_X1 U2320 ( .A1(RST), .A2(\DP/NPC1[18] ), .ZN(\DP/RegNPC1/N21 ) );
  AND2_X1 U2321 ( .A1(RST), .A2(\DP/NPC1[19] ), .ZN(\DP/RegNPC1/N22 ) );
  AND2_X1 U2322 ( .A1(RST), .A2(\DP/NPC1[20] ), .ZN(\DP/RegNPC1/N23 ) );
  AND2_X1 U2323 ( .A1(RST), .A2(w_PC_OUT[21]), .ZN(\DP/RegNPC1/N24 ) );
  AND2_X1 U2324 ( .A1(RST), .A2(\DP/NPC1[22] ), .ZN(\DP/RegNPC1/N25 ) );
  AND2_X1 U2325 ( .A1(RST), .A2(\DP/NPC1[23] ), .ZN(\DP/RegNPC1/N26 ) );
  AND2_X1 U2326 ( .A1(RST), .A2(\DP/NPC1[24] ), .ZN(\DP/RegNPC1/N27 ) );
  AND2_X1 U2327 ( .A1(RST), .A2(\DP/NPC1[25] ), .ZN(\DP/RegNPC1/N28 ) );
  AND2_X1 U2328 ( .A1(RST), .A2(\DP/NPC1[26] ), .ZN(\DP/RegNPC1/N29 ) );
  AND2_X1 U2329 ( .A1(RST), .A2(\DP/NPC1[0] ), .ZN(\DP/RegNPC1/N3 ) );
  AND2_X1 U2330 ( .A1(RST), .A2(\DP/NPC1[27] ), .ZN(\DP/RegNPC1/N30 ) );
  AND2_X1 U2331 ( .A1(RST), .A2(\DP/NPC1[28] ), .ZN(\DP/RegNPC1/N31 ) );
  AND2_X1 U2332 ( .A1(RST), .A2(\DP/NPC1[29] ), .ZN(\DP/RegNPC1/N32 ) );
  AND2_X1 U2333 ( .A1(RST), .A2(\DP/NPC1[30] ), .ZN(\DP/RegNPC1/N33 ) );
  AND2_X1 U2334 ( .A1(RST), .A2(\DP/NPC1[31] ), .ZN(\DP/RegNPC1/N34 ) );
  AND2_X1 U2335 ( .A1(RST), .A2(\DP/NPC1[1] ), .ZN(\DP/RegNPC1/N4 ) );
  AND2_X1 U2336 ( .A1(RST), .A2(\DP/NPC1[2] ), .ZN(\DP/RegNPC1/N5 ) );
  AND2_X1 U2337 ( .A1(RST), .A2(\DP/NPC1[3] ), .ZN(\DP/RegNPC1/N6 ) );
  AND2_X1 U2338 ( .A1(RST), .A2(\DP/NPC1[4] ), .ZN(\DP/RegNPC1/N7 ) );
  AND2_X1 U2339 ( .A1(RST), .A2(\DP/NPC1[5] ), .ZN(\DP/RegNPC1/N8 ) );
  AND2_X1 U2340 ( .A1(RST), .A2(\DP/NPC1[6] ), .ZN(\DP/RegNPC1/N9 ) );
  AND2_X1 U2341 ( .A1(RST), .A2(\DP/NPC2[7] ), .ZN(\DP/RegNPC2/N10 ) );
  AND2_X1 U2342 ( .A1(RST), .A2(\DP/NPC2[8] ), .ZN(\DP/RegNPC2/N11 ) );
  AND2_X1 U2343 ( .A1(RST), .A2(\DP/NPC2[9] ), .ZN(\DP/RegNPC2/N12 ) );
  AND2_X1 U2344 ( .A1(RST), .A2(\DP/NPC2[10] ), .ZN(\DP/RegNPC2/N13 ) );
  AND2_X1 U2345 ( .A1(RST), .A2(\DP/NPC2[11] ), .ZN(\DP/RegNPC2/N14 ) );
  AND2_X1 U2346 ( .A1(RST), .A2(\DP/NPC2[12] ), .ZN(\DP/RegNPC2/N15 ) );
  AND2_X1 U2347 ( .A1(RST), .A2(\DP/NPC2[13] ), .ZN(\DP/RegNPC2/N16 ) );
  AND2_X1 U2348 ( .A1(RST), .A2(\DP/NPC2[14] ), .ZN(\DP/RegNPC2/N17 ) );
  AND2_X1 U2349 ( .A1(RST), .A2(\DP/NPC2[15] ), .ZN(\DP/RegNPC2/N18 ) );
  AND2_X1 U2350 ( .A1(RST), .A2(\DP/NPC2[16] ), .ZN(\DP/RegNPC2/N19 ) );
  AND2_X1 U2351 ( .A1(RST), .A2(\DP/NPC2[17] ), .ZN(\DP/RegNPC2/N20 ) );
  AND2_X1 U2352 ( .A1(RST), .A2(\DP/NPC2[18] ), .ZN(\DP/RegNPC2/N21 ) );
  AND2_X1 U2353 ( .A1(RST), .A2(\DP/NPC2[19] ), .ZN(\DP/RegNPC2/N22 ) );
  AND2_X1 U2354 ( .A1(RST), .A2(\DP/NPC2[20] ), .ZN(\DP/RegNPC2/N23 ) );
  AND2_X1 U2355 ( .A1(RST), .A2(\DP/NPC2[21] ), .ZN(\DP/RegNPC2/N24 ) );
  AND2_X1 U2356 ( .A1(RST), .A2(\DP/NPC2[22] ), .ZN(\DP/RegNPC2/N25 ) );
  AND2_X1 U2357 ( .A1(RST), .A2(\DP/NPC2[23] ), .ZN(\DP/RegNPC2/N26 ) );
  AND2_X1 U2358 ( .A1(RST), .A2(\DP/NPC2[24] ), .ZN(\DP/RegNPC2/N27 ) );
  AND2_X1 U2359 ( .A1(RST), .A2(\DP/NPC2[25] ), .ZN(\DP/RegNPC2/N28 ) );
  AND2_X1 U2360 ( .A1(RST), .A2(\DP/NPC2[26] ), .ZN(\DP/RegNPC2/N29 ) );
  AND2_X1 U2361 ( .A1(RST), .A2(\DP/NPC2[0] ), .ZN(\DP/RegNPC2/N3 ) );
  AND2_X1 U2362 ( .A1(RST), .A2(\DP/NPC2[27] ), .ZN(\DP/RegNPC2/N30 ) );
  AND2_X1 U2363 ( .A1(RST), .A2(\DP/NPC2[28] ), .ZN(\DP/RegNPC2/N31 ) );
  AND2_X1 U2364 ( .A1(RST), .A2(\DP/NPC2[29] ), .ZN(\DP/RegNPC2/N32 ) );
  AND2_X1 U2365 ( .A1(RST), .A2(\DP/NPC2[30] ), .ZN(\DP/RegNPC2/N33 ) );
  AND2_X1 U2366 ( .A1(RST), .A2(\DP/NPC2[31] ), .ZN(\DP/RegNPC2/N34 ) );
  AND2_X1 U2367 ( .A1(RST), .A2(\DP/NPC2[1] ), .ZN(\DP/RegNPC2/N4 ) );
  AND2_X1 U2368 ( .A1(RST), .A2(\DP/NPC2[2] ), .ZN(\DP/RegNPC2/N5 ) );
  AND2_X1 U2369 ( .A1(RST), .A2(\DP/NPC2[3] ), .ZN(\DP/RegNPC2/N6 ) );
  AND2_X1 U2370 ( .A1(RST), .A2(\DP/NPC2[4] ), .ZN(\DP/RegNPC2/N7 ) );
  AND2_X1 U2371 ( .A1(RST), .A2(\DP/NPC2[5] ), .ZN(\DP/RegNPC2/N8 ) );
  AND2_X1 U2372 ( .A1(RST), .A2(\DP/NPC2[6] ), .ZN(\DP/RegNPC2/N9 ) );
  AND2_X1 U2373 ( .A1(RST), .A2(\DP/NPC3[7] ), .ZN(\DP/RegNPC3/N10 ) );
  AND2_X1 U2374 ( .A1(RST), .A2(\DP/NPC3[8] ), .ZN(\DP/RegNPC3/N11 ) );
  AND2_X1 U2375 ( .A1(RST), .A2(\DP/NPC3[9] ), .ZN(\DP/RegNPC3/N12 ) );
  AND2_X1 U2376 ( .A1(RST), .A2(\DP/NPC3[10] ), .ZN(\DP/RegNPC3/N13 ) );
  AND2_X1 U2377 ( .A1(RST), .A2(\DP/NPC3[11] ), .ZN(\DP/RegNPC3/N14 ) );
  AND2_X1 U2378 ( .A1(RST), .A2(\DP/NPC3[12] ), .ZN(\DP/RegNPC3/N15 ) );
  AND2_X1 U2379 ( .A1(RST), .A2(\DP/NPC3[13] ), .ZN(\DP/RegNPC3/N16 ) );
  AND2_X1 U2380 ( .A1(RST), .A2(\DP/NPC3[14] ), .ZN(\DP/RegNPC3/N17 ) );
  AND2_X1 U2381 ( .A1(RST), .A2(\DP/NPC3[15] ), .ZN(\DP/RegNPC3/N18 ) );
  AND2_X1 U2382 ( .A1(RST), .A2(\DP/NPC3[16] ), .ZN(\DP/RegNPC3/N19 ) );
  OR2_X1 U2383 ( .A1(\DP/JL1 ), .A2(n640), .ZN(\DP/RegNPC3/N2 ) );
  AND2_X1 U2384 ( .A1(RST), .A2(\DP/NPC3[17] ), .ZN(\DP/RegNPC3/N20 ) );
  AND2_X1 U2385 ( .A1(RST), .A2(\DP/NPC3[18] ), .ZN(\DP/RegNPC3/N21 ) );
  AND2_X1 U2386 ( .A1(RST), .A2(\DP/NPC3[19] ), .ZN(\DP/RegNPC3/N22 ) );
  AND2_X1 U2387 ( .A1(RST), .A2(\DP/NPC3[20] ), .ZN(\DP/RegNPC3/N23 ) );
  AND2_X1 U2388 ( .A1(RST), .A2(\DP/NPC3[21] ), .ZN(\DP/RegNPC3/N24 ) );
  AND2_X1 U2389 ( .A1(RST), .A2(\DP/NPC3[22] ), .ZN(\DP/RegNPC3/N25 ) );
  AND2_X1 U2390 ( .A1(RST), .A2(\DP/NPC3[23] ), .ZN(\DP/RegNPC3/N26 ) );
  AND2_X1 U2391 ( .A1(RST), .A2(\DP/NPC3[24] ), .ZN(\DP/RegNPC3/N27 ) );
  AND2_X1 U2392 ( .A1(RST), .A2(\DP/NPC3[25] ), .ZN(\DP/RegNPC3/N28 ) );
  AND2_X1 U2393 ( .A1(RST), .A2(\DP/NPC3[26] ), .ZN(\DP/RegNPC3/N29 ) );
  AND2_X1 U2394 ( .A1(RST), .A2(\DP/NPC3[0] ), .ZN(\DP/RegNPC3/N3 ) );
  AND2_X1 U2395 ( .A1(RST), .A2(\DP/NPC3[27] ), .ZN(\DP/RegNPC3/N30 ) );
  AND2_X1 U2396 ( .A1(RST), .A2(\DP/NPC3[28] ), .ZN(\DP/RegNPC3/N31 ) );
  AND2_X1 U2397 ( .A1(RST), .A2(\DP/NPC3[29] ), .ZN(\DP/RegNPC3/N32 ) );
  AND2_X1 U2398 ( .A1(RST), .A2(\DP/NPC3[30] ), .ZN(\DP/RegNPC3/N33 ) );
  AND2_X1 U2399 ( .A1(RST), .A2(\DP/NPC3[31] ), .ZN(\DP/RegNPC3/N34 ) );
  AND2_X1 U2400 ( .A1(RST), .A2(\DP/NPC3[1] ), .ZN(\DP/RegNPC3/N4 ) );
  AND2_X1 U2401 ( .A1(RST), .A2(\DP/NPC3[2] ), .ZN(\DP/RegNPC3/N5 ) );
  AND2_X1 U2402 ( .A1(RST), .A2(\DP/NPC3[3] ), .ZN(\DP/RegNPC3/N6 ) );
  AND2_X1 U2403 ( .A1(RST), .A2(\DP/NPC3[4] ), .ZN(\DP/RegNPC3/N7 ) );
  AND2_X1 U2404 ( .A1(RST), .A2(\DP/NPC3[5] ), .ZN(\DP/RegNPC3/N8 ) );
  AND2_X1 U2405 ( .A1(RST), .A2(\DP/NPC3[6] ), .ZN(\DP/RegNPC3/N9 ) );
  NAND3_X1 U2406 ( .A1(n1825), .A2(RST), .A3(n1201), .ZN(\DP/RegRD1/N2 ) );
  OR2_X1 U2413 ( .A1(w_RegRD2_LATCH_EN), .A2(n641), .ZN(\DP/RegRD2/N2 ) );
  NOR2_X1 U2415 ( .A1(n641), .A2(n599), .ZN(\DP/RegRD2/N4 ) );
  NOR2_X1 U2416 ( .A1(n641), .A2(n597), .ZN(\DP/RegRD2/N5 ) );
  AND2_X1 U2417 ( .A1(RST), .A2(\DP/RD1[3] ), .ZN(\DP/RegRD2/N6 ) );
  NOR2_X1 U2418 ( .A1(n641), .A2(n596), .ZN(\DP/RegRD2/N7 ) );
  OR2_X1 U2419 ( .A1(w_RegRD3_LATCH_EN), .A2(n641), .ZN(\DP/RegRD3/N2 ) );
  NOR2_X1 U2420 ( .A1(n640), .A2(n598), .ZN(\DP/RegRD3/N3 ) );
  NOR2_X1 U2421 ( .A1(n640), .A2(n594), .ZN(\DP/RegRD3/N4 ) );
  NOR2_X1 U2422 ( .A1(n640), .A2(n585), .ZN(\DP/RegRD3/N5 ) );
  NOR2_X1 U2423 ( .A1(n72), .A2(n641), .ZN(\DP/RegRD3/N6 ) );
  NOR2_X1 U2424 ( .A1(n73), .A2(n640), .ZN(\DP/RegRD3/N7 ) );
  NAND3_X1 U2425 ( .A1(n57), .A2(w_STORE_SIZE[1]), .A3(n606), .ZN(n1225) );
  NAND3_X1 U2426 ( .A1(n57), .A2(w_STORE_SIZE[0]), .A3(n603), .ZN(n1223) );
  NAND2_X1 U2427 ( .A1(n1225), .A2(n1223), .ZN(n1261) );
  NAND2_X1 U2428 ( .A1(\DP/FwdD ), .A2(n1261), .ZN(n1269) );
  INV_X1 U2429 ( .A(n1261), .ZN(n1222) );
  NOR2_X1 U2430 ( .A1(\DP/FwdD ), .A2(n1222), .ZN(n1266) );
  NAND2_X1 U2431 ( .A1(n1266), .A2(\DP/RegME_out[10] ), .ZN(n1211) );
  NOR3_X1 U2432 ( .A1(w_STORE_SIZE[1]), .A2(n57), .A3(w_STORE_SIZE[0]), .ZN(
        n1262) );
  OAI221_X1 U2433 ( .B1(\DP/FwdD ), .B2(\DP/RegME_out[7] ), .C1(n589), .C2(
        n1210), .A(n1262), .ZN(n1267) );
  OAI211_X1 U2434 ( .C1(n1501), .C2(n1269), .A(n1211), .B(n1267), .ZN(
        DRAM_DATA_OUT[10]) );
  NAND2_X1 U2435 ( .A1(n1266), .A2(\DP/RegME_out[11] ), .ZN(n1213) );
  OAI211_X1 U2436 ( .C1(n1214), .C2(n1269), .A(n1213), .B(n1267), .ZN(
        DRAM_DATA_OUT[11]) );
  NAND2_X1 U2437 ( .A1(n1266), .A2(\DP/RegME_out[12] ), .ZN(n1215) );
  OAI211_X1 U2438 ( .C1(n1216), .C2(n1269), .A(n1215), .B(n1267), .ZN(
        DRAM_DATA_OUT[12]) );
  NAND2_X1 U2439 ( .A1(n1266), .A2(\DP/RegME_out[13] ), .ZN(n1217) );
  OAI211_X1 U2440 ( .C1(n1218), .C2(n1269), .A(n1217), .B(n1267), .ZN(
        DRAM_DATA_OUT[13]) );
  NAND2_X1 U2441 ( .A1(n1266), .A2(\DP/RegME_out[14] ), .ZN(n1219) );
  OAI211_X1 U2442 ( .C1(n1462), .C2(n1269), .A(n1219), .B(n1267), .ZN(
        DRAM_DATA_OUT[14]) );
  AOI22_X1 U2443 ( .A1(\DP/FwdD ), .A2(n1221), .B1(\DP/RegME_out[15] ), .B2(
        n589), .ZN(n1224) );
  OAI21_X1 U2444 ( .B1(n1222), .B2(n1224), .A(n1267), .ZN(DRAM_DATA_OUT[15])
         );
  AOI21_X1 U2445 ( .B1(n1257), .B2(\DP/RegME_out[16] ), .A(n1256), .ZN(n1226)
         );
  OAI21_X1 U2446 ( .B1(n1227), .B2(n1259), .A(n1226), .ZN(DRAM_DATA_OUT[16])
         );
  AOI21_X1 U2447 ( .B1(n1257), .B2(\DP/RegME_out[17] ), .A(n1256), .ZN(n1228)
         );
  OAI21_X1 U2448 ( .B1(n1361), .B2(n1259), .A(n1228), .ZN(DRAM_DATA_OUT[17])
         );
  AOI21_X1 U2449 ( .B1(n1257), .B2(\DP/RegME_out[18] ), .A(n1256), .ZN(n1230)
         );
  OAI21_X1 U2450 ( .B1(n1336), .B2(n1259), .A(n1230), .ZN(DRAM_DATA_OUT[18])
         );
  AOI21_X1 U2451 ( .B1(n1257), .B2(\DP/RegME_out[19] ), .A(n1256), .ZN(n1232)
         );
  OAI21_X1 U2452 ( .B1(n1233), .B2(n1259), .A(n1232), .ZN(DRAM_DATA_OUT[19])
         );
  AOI21_X1 U2453 ( .B1(n1257), .B2(\DP/RegME_out[20] ), .A(n1256), .ZN(n1234)
         );
  OAI21_X1 U2454 ( .B1(n1454), .B2(n1259), .A(n1234), .ZN(DRAM_DATA_OUT[20])
         );
  AOI21_X1 U2455 ( .B1(n1257), .B2(\DP/RegME_out[21] ), .A(n1256), .ZN(n1236)
         );
  OAI21_X1 U2456 ( .B1(n1319), .B2(n1259), .A(n1236), .ZN(DRAM_DATA_OUT[21])
         );
  AOI21_X1 U2457 ( .B1(n1257), .B2(\DP/RegME_out[22] ), .A(n1256), .ZN(n1238)
         );
  OAI21_X1 U2458 ( .B1(n1292), .B2(n1259), .A(n1238), .ZN(DRAM_DATA_OUT[22])
         );
  AOI21_X1 U2459 ( .B1(n1257), .B2(\DP/RegME_out[23] ), .A(n1256), .ZN(n1240)
         );
  OAI21_X1 U2460 ( .B1(n1433), .B2(n1259), .A(n1240), .ZN(DRAM_DATA_OUT[23])
         );
  AOI21_X1 U2461 ( .B1(n1257), .B2(\DP/RegME_out[24] ), .A(n1256), .ZN(n1242)
         );
  OAI21_X1 U2462 ( .B1(n1318), .B2(n1259), .A(n1242), .ZN(DRAM_DATA_OUT[24])
         );
  AOI21_X1 U2463 ( .B1(n1257), .B2(\DP/RegME_out[25] ), .A(n1256), .ZN(n1244)
         );
  OAI21_X1 U2464 ( .B1(n1453), .B2(n1259), .A(n1244), .ZN(DRAM_DATA_OUT[25])
         );
  AOI21_X1 U2465 ( .B1(n1257), .B2(\DP/RegME_out[26] ), .A(n1256), .ZN(n1246)
         );
  OAI21_X1 U2466 ( .B1(n1247), .B2(n1259), .A(n1246), .ZN(DRAM_DATA_OUT[26])
         );
  AOI21_X1 U2467 ( .B1(n1257), .B2(\DP/RegME_out[27] ), .A(n1256), .ZN(n1248)
         );
  OAI21_X1 U2468 ( .B1(n1458), .B2(n1259), .A(n1248), .ZN(DRAM_DATA_OUT[27])
         );
  AOI21_X1 U2469 ( .B1(n1257), .B2(\DP/RegME_out[28] ), .A(n1256), .ZN(n1250)
         );
  OAI21_X1 U2470 ( .B1(n1305), .B2(n1259), .A(n1250), .ZN(DRAM_DATA_OUT[28])
         );
  AOI21_X1 U2471 ( .B1(n1257), .B2(\DP/RegME_out[29] ), .A(n1256), .ZN(n1252)
         );
  OAI21_X1 U2472 ( .B1(n1253), .B2(n1259), .A(n1252), .ZN(DRAM_DATA_OUT[29])
         );
  AOI21_X1 U2473 ( .B1(n1257), .B2(\DP/RegME_out[30] ), .A(n1256), .ZN(n1254)
         );
  OAI21_X1 U2474 ( .B1(n1255), .B2(n1259), .A(n1254), .ZN(DRAM_DATA_OUT[30])
         );
  AOI21_X1 U2475 ( .B1(n1257), .B2(\DP/RegME_out[31] ), .A(n1256), .ZN(n1258)
         );
  OAI21_X1 U2476 ( .B1(n1356), .B2(n1259), .A(n1258), .ZN(DRAM_DATA_OUT[31])
         );
  OAI21_X1 U2477 ( .B1(n1262), .B2(n1261), .A(\DP/FwdD ), .ZN(n1278) );
  OAI21_X1 U2478 ( .B1(n1262), .B2(n1261), .A(n589), .ZN(n1277) );
  OAI22_X1 U2479 ( .A1(n1263), .A2(n1278), .B1(n1277), .B2(n610), .ZN(
        DRAM_DATA_OUT[7]) );
  NAND2_X1 U2480 ( .A1(n1266), .A2(\DP/RegME_out[8] ), .ZN(n1264) );
  OAI211_X1 U2481 ( .C1(n1471), .C2(n1269), .A(n1264), .B(n1267), .ZN(
        DRAM_DATA_OUT[8]) );
  NAND2_X1 U2482 ( .A1(n1266), .A2(\DP/RegME_out[9] ), .ZN(n1268) );
  OAI211_X1 U2483 ( .C1(n1456), .C2(n1269), .A(n1268), .B(n1267), .ZN(
        DRAM_DATA_OUT[9]) );
  OAI22_X1 U2484 ( .A1(n1271), .A2(n1278), .B1(n611), .B2(n1277), .ZN(
        DRAM_DATA_OUT[0]) );
  OAI22_X1 U2485 ( .A1(n1272), .A2(n1278), .B1(n612), .B2(n1277), .ZN(
        DRAM_DATA_OUT[1]) );
  OAI22_X1 U2487 ( .A1(n1449), .A2(n1278), .B1(n614), .B2(n1277), .ZN(
        DRAM_DATA_OUT[3]) );
  OAI22_X1 U2488 ( .A1(n1367), .A2(n1278), .B1(n615), .B2(n1277), .ZN(
        DRAM_DATA_OUT[4]) );
  OAI22_X1 U2489 ( .A1(n1415), .A2(n1278), .B1(n616), .B2(n1277), .ZN(
        DRAM_DATA_OUT[5]) );
  DFF_X1 \CU/cw1_reg[4]  ( .D(n1507), .CK(CLK), .Q(\CU/cw1[4] ) );
  DFF_X1 \CU/cw1_reg[1]  ( .D(n1506), .CK(CLK), .Q(\CU/cw1[1] ) );
  DFF_X1 \CU/cw2_reg[2]  ( .D(\CU/N66 ), .CK(CLK), .Q(\CU/cw2[2] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[0]  ( .D(\DP/RegNPC2/N3 ), .CK(
        \DP/RegNPC2/net7068 ), .Q(\DP/NPC3[0] ) );
  DFF_X2 \CU/cw1_reg[2]  ( .D(\CU/N42 ), .CK(CLK), .Q(\CU/cw1[2] ) );
  DFF_X2 \CU/cw1_reg[0]  ( .D(\CU/N42 ), .CK(CLK), .Q(w_RF_WE_EX) );
  DFF_X2 \DP/RegIMM/DOUT_reg[31]  ( .D(\DP/RegIMM/N34 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[31] ) );
  DFF_X2 \DP/RegIMM/DOUT_reg[24]  ( .D(\DP/RegIMM/N27 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[24] ) );
  DFF_X2 \DP/RegIMM/DOUT_reg[23]  ( .D(\DP/RegIMM/N26 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[23] ) );
  DFF_X2 \DP/RegIMM/DOUT_reg[22]  ( .D(\DP/RegIMM/N25 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[22] ) );
  DFF_X2 \DP/RegIMM/DOUT_reg[21]  ( .D(\DP/RegIMM/N24 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[21] ) );
  DFF_X2 \DP/RegIMM/DOUT_reg[20]  ( .D(\DP/RegIMM/N23 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[20] ) );
  DFF_X2 \DP/RegIMM/DOUT_reg[19]  ( .D(\DP/RegIMM/N22 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[19] ) );
  DFF_X2 \DP/RegIMM/DOUT_reg[18]  ( .D(\DP/RegIMM/N21 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[18] ) );
  DFF_X2 \DP/RegIMM/DOUT_reg[17]  ( .D(\DP/RegIMM/N20 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[17] ) );
  NAND3_X1 U1232 ( .A1(n1466), .A2(n1821), .A3(n1282), .ZN(n1573) );
  INV_X1 U1233 ( .A(n1400), .ZN(n1282) );
  NAND2_X1 U1257 ( .A1(n1495), .A2(n1284), .ZN(n678) );
  NAND2_X1 U1258 ( .A1(n1286), .A2(n1285), .ZN(n1284) );
  INV_X1 U1259 ( .A(IR_OUT[4]), .ZN(n1285) );
  INV_X1 U1260 ( .A(IR_OUT[5]), .ZN(n1286) );
  INV_X1 U1262 ( .A(n1288), .ZN(n1569) );
  OAI21_X1 U1263 ( .B1(n1580), .B2(n665), .A(n1289), .ZN(n1288) );
  NAND2_X1 U1285 ( .A1(n1546), .A2(n688), .ZN(n1580) );
  AND2_X1 U1289 ( .A1(n1484), .A2(n592), .ZN(n688) );
  INV_X1 U1300 ( .A(n1704), .ZN(n1703) );
  NOR2_X1 U1301 ( .A1(n1707), .A2(n1705), .ZN(n1704) );
  NOR2_X2 U1311 ( .A1(n1812), .A2(n1291), .ZN(n1290) );
  INV_X2 U1315 ( .A(n1290), .ZN(n1811) );
  NAND2_X1 U1317 ( .A1(n755), .A2(n1662), .ZN(n742) );
  OR2_X1 U1319 ( .A1(w_RF_RD2), .A2(n1722), .ZN(n1726) );
  BUF_X2 U1325 ( .A(n1493), .Z(n639) );
  CLKBUF_X1 U1327 ( .A(n1239), .Z(n1292) );
  NOR2_X1 U1330 ( .A1(n1294), .A2(n1293), .ZN(n1202) );
  OR2_X1 U1331 ( .A1(n1469), .A2(n1485), .ZN(n1293) );
  NAND2_X1 U1332 ( .A1(n1043), .A2(n1298), .ZN(n1294) );
  INV_X1 U1344 ( .A(n1205), .ZN(n1295) );
  INV_X1 U1346 ( .A(n1205), .ZN(n32) );
  NAND2_X1 U1347 ( .A1(n1544), .A2(IR_OUT[18]), .ZN(n1205) );
  CLKBUF_X1 U1349 ( .A(n935), .Z(n1296) );
  NOR2_X1 U1350 ( .A1(n1645), .A2(n1205), .ZN(n1640) );
  NOR3_X1 U1351 ( .A1(n675), .A2(n674), .A3(n668), .ZN(n1297) );
  NOR3_X1 U1352 ( .A1(n675), .A2(n674), .A3(n668), .ZN(n1046) );
  INV_X1 U1354 ( .A(n1572), .ZN(n1298) );
  CLKBUF_X1 U1355 ( .A(n714), .Z(n1545) );
  INV_X1 U1356 ( .A(n1540), .ZN(n751) );
  OR3_X1 U1357 ( .A1(n752), .A2(n1310), .A3(n648), .ZN(n1469) );
  BUF_X1 U1359 ( .A(n697), .Z(n1299) );
  NAND2_X1 U1363 ( .A1(n966), .A2(n1553), .ZN(\DP/RF_DATA[3] ) );
  CLKBUF_X2 U1364 ( .A(w_MuxWB_SEL), .Z(n1494) );
  BUF_X1 U1365 ( .A(n1333), .Z(n1463) );
  AND2_X1 U1366 ( .A1(n1331), .A2(n1556), .ZN(n1555) );
  NOR2_X1 U1367 ( .A1(n1369), .A2(n1709), .ZN(n1708) );
  NOR2_X1 U1368 ( .A1(n898), .A2(n1366), .ZN(n1300) );
  INV_X1 U1371 ( .A(n35), .ZN(n1301) );
  NAND2_X1 U1372 ( .A1(n941), .A2(n940), .ZN(n1302) );
  NOR2_X1 U1373 ( .A1(n1302), .A2(n1303), .ZN(\DP/RegFB/N4 ) );
  OR2_X1 U1374 ( .A1(n1304), .A2(n1036), .ZN(n1303) );
  INV_X1 U1375 ( .A(RST), .ZN(n1304) );
  INV_X2 U1376 ( .A(\DP/NPC1[15] ), .ZN(n1761) );
  INV_X1 U1377 ( .A(n1761), .ZN(n1750) );
  NAND2_X1 U1378 ( .A1(n1736), .A2(n1775), .ZN(n1735) );
  NAND2_X1 U1379 ( .A1(n1736), .A2(n1701), .ZN(n1700) );
  CLKBUF_X1 U1380 ( .A(n1251), .Z(n1305) );
  NOR2_X1 U1381 ( .A1(n1411), .A2(n1412), .ZN(n1251) );
  INV_X1 U1382 ( .A(n1352), .ZN(n1306) );
  OR2_X1 U1383 ( .A1(n1307), .A2(n674), .ZN(n676) );
  NAND2_X1 U1384 ( .A1(n1306), .A2(n1039), .ZN(n1307) );
  OAI21_X1 U1385 ( .B1(n1276), .B2(\DP/JL2 ), .A(n968), .ZN(\DP/RF_DATA[5] )
         );
  OAI22_X1 U1386 ( .A1(n1654), .A2(n1278), .B1(n617), .B2(n1277), .ZN(
        DRAM_DATA_OUT[6]) );
  OR2_X1 U1387 ( .A1(n1492), .A2(n1654), .ZN(n1646) );
  NOR2_X1 U1390 ( .A1(n630), .A2(n1654), .ZN(n1648) );
  NOR2_X1 U1391 ( .A1(n621), .A2(n1654), .ZN(n1650) );
  NOR2_X1 U1392 ( .A1(n626), .A2(n1654), .ZN(n1653) );
  OR2_X1 U1393 ( .A1(n1097), .A2(n1719), .ZN(n1308) );
  OR2_X2 U1394 ( .A1(n1308), .A2(n1309), .ZN(n1153) );
  OR2_X1 U1397 ( .A1(n1735), .A2(n1732), .ZN(n1309) );
  NOR3_X1 U1399 ( .A1(n704), .A2(n1564), .A3(n665), .ZN(n1310) );
  OAI211_X1 U1400 ( .C1(n1691), .C2(n1678), .A(n1677), .B(n59), .ZN(n1676) );
  NAND2_X1 U1401 ( .A1(n1691), .A2(w_JUMP_EQ), .ZN(n1677) );
  INV_X1 U1402 ( .A(n745), .ZN(n1311) );
  BUF_X1 U1403 ( .A(n737), .Z(n1312) );
  OR2_X1 U1404 ( .A1(n721), .A2(n1529), .ZN(n1528) );
  AOI211_X4 U1407 ( .C1(n1312), .C2(n735), .A(n734), .B(n733), .ZN(n743) );
  NAND3_X1 U1409 ( .A1(n1544), .A2(IR_OUT[5]), .A3(n595), .ZN(n1313) );
  NAND3_X1 U1410 ( .A1(n1544), .A2(IR_OUT[5]), .A3(n595), .ZN(n1314) );
  OR2_X1 U1424 ( .A1(n757), .A2(n1664), .ZN(n1315) );
  OR2_X1 U1427 ( .A1(n1274), .A2(n1492), .ZN(n1553) );
  NOR2_X1 U1429 ( .A1(n1645), .A2(n1206), .ZN(n1642) );
  NOR2_X1 U1431 ( .A1(n1206), .A2(n584), .ZN(n1605) );
  AND2_X1 U1432 ( .A1(n1514), .A2(n1518), .ZN(n903) );
  AND2_X1 U1434 ( .A1(n1570), .A2(n653), .ZN(n1316) );
  CLKBUF_X1 U1436 ( .A(n1461), .Z(n1317) );
  CLKBUF_X1 U1437 ( .A(n1243), .Z(n1318) );
  BUF_X1 U1438 ( .A(n1241), .Z(n1433) );
  OR2_X1 U1439 ( .A1(n1241), .A2(n1488), .ZN(n1523) );
  NOR2_X1 U1441 ( .A1(n1742), .A2(n1761), .ZN(n1740) );
  NAND2_X1 U1442 ( .A1(n1762), .A2(n1743), .ZN(n1742) );
  CLKBUF_X1 U1443 ( .A(n1237), .Z(n1319) );
  AND2_X1 U1463 ( .A1(n1499), .A2(n1320), .ZN(n1372) );
  NOR2_X1 U1471 ( .A1(n1724), .A2(n1321), .ZN(n1320) );
  INV_X32 U1475 ( .A(n1373), .ZN(n1321) );
  INV_X4 U1482 ( .A(n641), .ZN(n1373) );
  INV_X1 U1487 ( .A(n1724), .ZN(n1684) );
  OAI21_X1 U1492 ( .B1(n748), .B2(n757), .A(n728), .ZN(n1335) );
  CLKBUF_X1 U1494 ( .A(n723), .Z(n1322) );
  CLKBUF_X1 U1499 ( .A(n1118), .Z(n1323) );
  NOR2_X1 U1501 ( .A1(n1118), .A2(n1761), .ZN(n1324) );
  AND2_X1 U1509 ( .A1(n660), .A2(n586), .ZN(n1327) );
  AND3_X1 U1510 ( .A1(n1353), .A2(n1668), .A3(n1728), .ZN(n1328) );
  CLKBUF_X1 U1511 ( .A(n703), .Z(n1549) );
  NOR2_X1 U1512 ( .A1(n901), .A2(n899), .ZN(n1514) );
  INV_X1 U1517 ( .A(n1697), .ZN(n1802) );
  AOI21_X1 U1519 ( .B1(n761), .B2(n1657), .A(n760), .ZN(n763) );
  NAND3_X2 U1527 ( .A1(IR_OUT[15]), .A2(RST), .A3(n1045), .ZN(n1050) );
  CLKBUF_X1 U1534 ( .A(n1485), .Z(n1343) );
  CLKBUF_X1 U1550 ( .A(n678), .Z(n1329) );
  AND2_X2 U1611 ( .A1(w_PC_OUT[27]), .A2(w_PC_OUT[28]), .ZN(n1817) );
  INV_X1 U1619 ( .A(n1814), .ZN(n1813) );
  OR2_X4 U1622 ( .A1(n1798), .A2(n1800), .ZN(n1797) );
  AND2_X1 U1643 ( .A1(n1330), .A2(n666), .ZN(n1331) );
  NAND2_X1 U1646 ( .A1(n1495), .A2(n1692), .ZN(n1332) );
  NAND2_X1 U1725 ( .A1(n1694), .A2(n1693), .ZN(n1692) );
  OR2_X1 U1741 ( .A1(n645), .A2(n1590), .ZN(n1333) );
  NAND2_X1 U1755 ( .A1(n729), .A2(n1334), .ZN(\CU/N86 ) );
  INV_X2 U1756 ( .A(n1335), .ZN(n1334) );
  CLKBUF_X3 U1757 ( .A(n1231), .Z(n1336) );
  INV_X1 U1758 ( .A(n1337), .ZN(n1027) );
  NAND4_X1 U1763 ( .A1(n1342), .A2(n1341), .A3(n1340), .A4(n1019), .ZN(n1337)
         );
  NAND2_X1 U1764 ( .A1(n1338), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1765 ( .A1(n1016), .A2(n1339), .ZN(n1338) );
  XNOR2_X1 U1768 ( .A(n1051), .B(\DP/RD1[4] ), .ZN(n1339) );
  INV_X1 U1769 ( .A(n1023), .ZN(n1340) );
  INV_X1 U1770 ( .A(n1025), .ZN(n1341) );
  INV_X1 U1771 ( .A(n1024), .ZN(n1342) );
  OR2_X2 U1772 ( .A1(n1344), .A2(n1345), .ZN(\DP/RF_DATA[2] ) );
  NOR2_X1 U1773 ( .A1(n1488), .A2(n1632), .ZN(n1344) );
  AND2_X1 U1774 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[2] ), .ZN(n1345) );
  AND3_X2 U1775 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1711) );
  AND2_X1 U1779 ( .A1(n1276), .A2(n1654), .ZN(n1346) );
  AND4_X1 U1780 ( .A1(n1255), .A2(n1253), .A3(n1251), .A4(n1249), .ZN(n1347)
         );
  AND4_X1 U1781 ( .A1(n1270), .A2(n1265), .A3(n985), .A4(n1260), .ZN(n1348) );
  BUF_X1 U1782 ( .A(n1563), .Z(n1350) );
  AND3_X2 U1783 ( .A1(IROM_ADDR[0]), .A2(\DP/NPC1[1] ), .A3(\DP/NPC1[2] ), 
        .ZN(n1351) );
  INV_X4 U1786 ( .A(n1351), .ZN(n1181) );
  NAND4_X1 U1787 ( .A1(n1609), .A2(n1608), .A3(n1600), .A4(n1599), .ZN(n1598)
         );
  AOI21_X1 U1788 ( .B1(n34), .B2(n594), .A(n1601), .ZN(n1600) );
  NOR2_X1 U1789 ( .A1(n1645), .A2(n1203), .ZN(n1636) );
  OAI21_X1 U1790 ( .B1(n1203), .B2(\DP/RD2[0] ), .A(n1020), .ZN(n1607) );
  NOR2_X1 U1791 ( .A1(n1580), .A2(n1844), .ZN(n1352) );
  CLKBUF_X1 U1794 ( .A(n1825), .Z(n1354) );
  BUF_X2 U1795 ( .A(w_MuxWB_SEL), .Z(n1493) );
  INV_X1 U1797 ( .A(n1133), .ZN(n1132) );
  AND3_X2 U1804 ( .A1(n1324), .A2(n1743), .A3(w_PC_OUT[17]), .ZN(n1129) );
  NAND2_X1 U1805 ( .A1(n1718), .A2(n1717), .ZN(n1716) );
  INV_X1 U1807 ( .A(n1112), .ZN(n1111) );
  AND2_X1 U1817 ( .A1(n1112), .A2(\DP/NPC1[13] ), .ZN(n1115) );
  INV_X1 U1835 ( .A(n1466), .ZN(n681) );
  CLKBUF_X1 U1841 ( .A(n1260), .Z(n1356) );
  OR2_X1 U1845 ( .A1(n1800), .A2(n1357), .ZN(n1358) );
  INV_X1 U1848 ( .A(n1789), .ZN(n1357) );
  NOR4_X1 U1851 ( .A1(n1118), .A2(n1761), .A3(n1752), .A4(n1745), .ZN(n1359)
         );
  NOR4_X1 U1853 ( .A1(n1118), .A2(n1761), .A3(n1752), .A4(n1745), .ZN(n1360)
         );
  NOR4_X1 U1857 ( .A1(n1118), .A2(n1761), .A3(n1752), .A4(n1745), .ZN(n1147)
         );
  CLKBUF_X1 U1861 ( .A(n1229), .Z(n1361) );
  OR2_X1 U1863 ( .A1(n707), .A2(n1555), .ZN(n1554) );
  NAND2_X1 U1874 ( .A1(n1495), .A2(n1587), .ZN(n1586) );
  NAND3_X1 U1952 ( .A1(n908), .A2(n909), .A3(n910), .ZN(n1362) );
  NAND2_X1 U1960 ( .A1(n911), .A2(n1363), .ZN(n917) );
  INV_X1 U2033 ( .A(n1362), .ZN(n1363) );
  AND4_X2 U2034 ( .A1(n1401), .A2(n1402), .A3(n1403), .A4(n1404), .ZN(n910) );
  AND4_X2 U2035 ( .A1(n1382), .A2(n1383), .A3(n1384), .A4(n1385), .ZN(n908) );
  CLKBUF_X1 U2037 ( .A(n1494), .Z(n1364) );
  NOR2_X1 U2043 ( .A1(n1210), .A2(n942), .ZN(n1365) );
  NOR2_X1 U2050 ( .A1(n898), .A2(n1366), .ZN(n904) );
  INV_X1 U2051 ( .A(n1365), .ZN(n1366) );
  INV_X1 U2056 ( .A(n1623), .ZN(n1367) );
  CLKBUF_X1 U2070 ( .A(n1042), .Z(n1368) );
  AOI21_X1 U2121 ( .B1(n1370), .B2(n1371), .A(n1416), .ZN(n1369) );
  AND4_X1 U2182 ( .A1(n925), .A2(n924), .A3(n923), .A4(n922), .ZN(n1370) );
  AND4_X1 U2183 ( .A1(n921), .A2(n920), .A3(n919), .A4(n918), .ZN(n1371) );
  INV_X1 U2184 ( .A(n1416), .ZN(n1008) );
  AND4_X1 U2185 ( .A1(n1390), .A2(n1391), .A3(n1392), .A4(n1393), .ZN(n922) );
  AOI21_X1 U2186 ( .B1(n639), .B2(\DP/RegLMD_out[6] ), .A(n1655), .ZN(n1654)
         );
  NOR2_X1 U2187 ( .A1(n723), .A2(n1657), .ZN(n760) );
  INV_X1 U2192 ( .A(n1328), .ZN(n1581) );
  NAND2_X1 U2195 ( .A1(n1372), .A2(n1685), .ZN(\DP/RegA/N2 ) );
  CLKBUF_X1 U2200 ( .A(n1830), .Z(n1374) );
  AND2_X1 U2203 ( .A1(\DP/RegALU2_out[6] ), .A2(n583), .ZN(n1655) );
  CLKBUF_X1 U2208 ( .A(n660), .Z(n1375) );
  AND4_X1 U2211 ( .A1(n1376), .A2(n1377), .A3(n1378), .A4(n1379), .ZN(n921) );
  INV_X1 U2216 ( .A(n1815), .ZN(n1800) );
  NAND2_X1 U2219 ( .A1(n1815), .A2(w_PC_OUT[30]), .ZN(n1814) );
  CLKBUF_X1 U2224 ( .A(n713), .Z(n1380) );
  AND4_X1 U2233 ( .A1(n1386), .A2(n1387), .A3(n1388), .A4(n1389), .ZN(n923) );
  AND4_X1 U2236 ( .A1(n1394), .A2(n1395), .A3(n1396), .A4(n1397), .ZN(n915) );
  INV_X1 U2244 ( .A(n678), .ZN(n1400) );
  AND4_X1 U2252 ( .A1(n1407), .A2(n1408), .A3(n1409), .A4(n1410), .ZN(n909) );
  AND2_X1 U2257 ( .A1(n639), .A2(\DP/RegLMD_out[28] ), .ZN(n1411) );
  AND2_X1 U2260 ( .A1(\DP/RegALU2_out[28] ), .A2(n583), .ZN(n1412) );
  CLKBUF_X1 U2266 ( .A(n1276), .Z(n1415) );
  INV_X1 U2271 ( .A(n1745), .ZN(n1743) );
  NAND3_X1 U2275 ( .A1(\DP/FwdA[2] ), .A2(n69), .A3(n76), .ZN(n1416) );
  BUF_X2 U2276 ( .A(n1008), .Z(n628) );
  AND2_X1 U2277 ( .A1(n639), .A2(\DP/RegLMD_out[31] ), .ZN(n1417) );
  AND2_X1 U2278 ( .A1(\DP/RegALU2_out[31] ), .A2(n583), .ZN(n1418) );
  NOR2_X2 U2279 ( .A1(n1417), .A2(n1418), .ZN(n1260) );
  NAND2_X1 U2282 ( .A1(n1330), .A2(n1350), .ZN(n1419) );
  INV_X1 U2283 ( .A(n1816), .ZN(n1815) );
  AND4_X1 U2285 ( .A1(n1420), .A2(n1421), .A3(n1422), .A4(n1423), .ZN(n918) );
  AND4_X1 U2286 ( .A1(n1424), .A2(n1425), .A3(n1426), .A4(n1427), .ZN(n912) );
  AND4_X2 U2407 ( .A1(n1428), .A2(n1429), .A3(n1430), .A4(n1431), .ZN(n920) );
  BUF_X1 U2408 ( .A(n750), .Z(n1432) );
  NAND2_X2 U2409 ( .A1(n943), .A2(n1511), .ZN(\DP/RF_DATA[10] ) );
  AND4_X1 U2410 ( .A1(n1434), .A2(n1435), .A3(n1436), .A4(n1437), .ZN(n913) );
  AND4_X1 U2411 ( .A1(n1438), .A2(n1439), .A3(n1440), .A4(n1441), .ZN(n919) );
  AND4_X1 U2412 ( .A1(n1442), .A2(n1443), .A3(n1444), .A4(n1445), .ZN(n914) );
  INV_X1 U2414 ( .A(n679), .ZN(n1446) );
  OR2_X2 U2486 ( .A1(n682), .A2(n1447), .ZN(n736) );
  CLKBUF_X1 U2490 ( .A(n1713), .Z(n1540) );
  INV_X1 U2492 ( .A(n1274), .ZN(n1448) );
  INV_X2 U2493 ( .A(n1448), .ZN(n1449) );
  NAND2_X1 U2494 ( .A1(n1763), .A2(n1760), .ZN(n1759) );
  INV_X1 U2495 ( .A(n1736), .ZN(n1707) );
  NOR2_X1 U2496 ( .A1(n1761), .A2(n1755), .ZN(n1760) );
  OAI21_X1 U2497 ( .B1(n1118), .B2(n1739), .A(n1741), .ZN(n1450) );
  BUF_X1 U2498 ( .A(n652), .Z(n1451) );
  CLKBUF_X1 U2499 ( .A(n1204), .Z(n1452) );
  OR2_X2 U2500 ( .A1(n1716), .A2(n1097), .ZN(n1118) );
  CLKBUF_X1 U2501 ( .A(n1245), .Z(n1453) );
  NAND2_X1 U2502 ( .A1(n1208), .A2(n593), .ZN(n1603) );
  NOR2_X1 U2503 ( .A1(n1645), .A2(n1301), .ZN(n1644) );
  CLKBUF_X1 U2504 ( .A(n1235), .Z(n1454) );
  INV_X1 U2505 ( .A(n1463), .ZN(n1455) );
  CLKBUF_X1 U2506 ( .A(n1270), .Z(n1456) );
  NOR2_X1 U2507 ( .A1(n1104), .A2(n1734), .ZN(n1108) );
  NOR3_X1 U2508 ( .A1(n1104), .A2(n1732), .A3(n1703), .ZN(n1150) );
  INV_X1 U2509 ( .A(n1732), .ZN(n1699) );
  INV_X1 U2510 ( .A(n1732), .ZN(n1701) );
  NAND2_X1 U2511 ( .A1(n719), .A2(n736), .ZN(n1527) );
  CLKBUF_X1 U2512 ( .A(n688), .Z(n1457) );
  NOR2_X1 U2513 ( .A1(n706), .A2(n1554), .ZN(n712) );
  CLKBUF_X1 U2514 ( .A(n1249), .Z(n1458) );
  OAI21_X1 U2516 ( .B1(n1129), .B2(n1128), .A(n1127), .ZN(n1460) );
  INV_X1 U2517 ( .A(n1829), .ZN(n655) );
  AND3_X1 U2518 ( .A1(n1590), .A2(n714), .A3(n62), .ZN(n1476) );
  NAND2_X1 U2519 ( .A1(n687), .A2(n1543), .ZN(n1461) );
  AOI21_X1 U2520 ( .B1(n639), .B2(\DP/RegLMD_out[14] ), .A(n1520), .ZN(n1462)
         );
  CLKBUF_X1 U2521 ( .A(n1455), .Z(n1464) );
  BUF_X1 U2522 ( .A(n1666), .Z(n1465) );
  OAI21_X1 U2523 ( .B1(n1467), .B2(n1468), .A(n1349), .ZN(n1466) );
  OR4_X2 U2524 ( .A1(IR_OUT[10]), .A2(IR_OUT[6]), .A3(IR_OUT[7]), .A4(
        IR_OUT[8]), .ZN(n1467) );
  CLKBUF_X1 U2525 ( .A(\CU/N55 ), .Z(n1486) );
  CLKBUF_X1 U2526 ( .A(n1463), .Z(n1470) );
  CLKBUF_X1 U2527 ( .A(n1265), .Z(n1471) );
  INV_X1 U2528 ( .A(n929), .ZN(n1709) );
  INV_X1 U2529 ( .A(n1740), .ZN(n1739) );
  BUF_X1 U2530 ( .A(n1054), .Z(n1472) );
  NAND2_X1 U2531 ( .A1(n1495), .A2(IR_OUT[3]), .ZN(n1054) );
  AND2_X1 U2532 ( .A1(n1332), .A2(n1686), .ZN(n1473) );
  AND2_X1 U2533 ( .A1(n1041), .A2(n1563), .ZN(n1474) );
  AND2_X1 U2536 ( .A1(n35), .A2(n596), .ZN(n1477) );
  AND2_X1 U2537 ( .A1(n1208), .A2(\DP/RD1[4] ), .ZN(n1478) );
  NOR3_X1 U2538 ( .A1(n1031), .A2(n1478), .A3(n1477), .ZN(n1032) );
  INV_X2 U2539 ( .A(n1208), .ZN(n35) );
  NOR2_X1 U2540 ( .A1(n1181), .A2(n1820), .ZN(n1189) );
  INV_X1 U2541 ( .A(n1181), .ZN(n1185) );
  INV_X1 U2542 ( .A(n1118), .ZN(n1119) );
  NAND2_X1 U2543 ( .A1(n1355), .A2(n1042), .ZN(w_RF_RD2) );
  OR2_X1 U2544 ( .A1(n1280), .A2(\DP/RD1[2] ), .ZN(n1479) );
  OR2_X1 U2545 ( .A1(n1048), .A2(\DP/RD1[1] ), .ZN(n1480) );
  NAND3_X1 U2546 ( .A1(n1479), .A2(n1480), .A3(n1015), .ZN(n1016) );
  OR2_X1 U2547 ( .A1(n739), .A2(n1830), .ZN(n1722) );
  NOR2_X1 U2549 ( .A1(\CU/JUMP3 ), .A2(\CU/JUMP2 ), .ZN(n1729) );
  NAND3_X1 U2550 ( .A1(n1353), .A2(n1668), .A3(n1728), .ZN(n1483) );
  NOR2_X1 U2552 ( .A1(n674), .A2(n1352), .ZN(n973) );
  INV_X1 U2553 ( .A(n1360), .ZN(n1146) );
  NAND2_X1 U2554 ( .A1(n1359), .A2(n1789), .ZN(n1161) );
  AND2_X1 U2555 ( .A1(n1484), .A2(n1669), .ZN(n666) );
  INV_X1 U2556 ( .A(n1689), .ZN(n1669) );
  NAND2_X1 U2557 ( .A1(n1472), .A2(n1053), .ZN(n716) );
  NAND2_X1 U2558 ( .A1(n1122), .A2(\DP/NPC1[16] ), .ZN(n1125) );
  NAND2_X1 U2559 ( .A1(n1041), .A2(n688), .ZN(n750) );
  INV_X1 U2560 ( .A(n1457), .ZN(n693) );
  INV_X1 U2561 ( .A(n1795), .ZN(n1794) );
  NOR2_X1 U2562 ( .A1(n1811), .A2(n1790), .ZN(n1789) );
  INV_X1 U2563 ( .A(w_PC_OUT[25]), .ZN(n1812) );
  AND2_X1 U2564 ( .A1(IR_OUT[27]), .A2(n1728), .ZN(n1576) );
  CLKBUF_X1 U2565 ( .A(n752), .Z(n1548) );
  NOR2_X1 U2566 ( .A1(n715), .A2(n1465), .ZN(n1661) );
  NAND2_X1 U2567 ( .A1(n736), .A2(n1465), .ZN(n732) );
  INV_X1 U2568 ( .A(\DP/NPC1[16] ), .ZN(n1745) );
  INV_X1 U2569 ( .A(\DP/NPC1[16] ), .ZN(n1755) );
  NAND4_X1 U2570 ( .A1(n1461), .A2(n1713), .A3(n1757), .A4(n1758), .ZN(n1485)
         );
  INV_X1 U2571 ( .A(n1582), .ZN(n674) );
  INV_X1 U2572 ( .A(n973), .ZN(n1724) );
  OR2_X1 U2573 ( .A1(n697), .A2(n1592), .ZN(n1579) );
  INV_X1 U2574 ( .A(IROM_ADDR[11]), .ZN(n1734) );
  INV_X1 U2575 ( .A(n1732), .ZN(n1731) );
  AND2_X1 U2576 ( .A1(n1147), .A2(n1776), .ZN(n1165) );
  INV_X2 U2577 ( .A(n1487), .ZN(n1488) );
  NAND3_X1 U2582 ( .A1(n1449), .A2(n1272), .A3(n1620), .ZN(n898) );
  NAND2_X1 U2583 ( .A1(n1514), .A2(n904), .ZN(n1513) );
  OR2_X1 U2585 ( .A1(n34), .A2(n599), .ZN(n1497) );
  OR2_X1 U2586 ( .A1(n1452), .A2(\DP/RD1[1] ), .ZN(n1498) );
  NAND3_X1 U2587 ( .A1(n1032), .A2(n1498), .A3(n1497), .ZN(n1034) );
  OAI21_X1 U2588 ( .B1(n1450), .B2(n1796), .A(n1173), .ZN(n1795) );
  INV_X1 U2589 ( .A(w_PC_OUT[27]), .ZN(n1793) );
  NAND2_X1 U2590 ( .A1(n1784), .A2(n1817), .ZN(n1810) );
  NAND2_X1 U2591 ( .A1(n1817), .A2(\DP/NPC1[29] ), .ZN(n1816) );
  NOR2_X1 U2592 ( .A1(n1469), .A2(n1485), .ZN(n1500) );
  OR2_X1 U2594 ( .A1(n1558), .A2(n1844), .ZN(n662) );
  INV_X1 U2595 ( .A(n1734), .ZN(n1733) );
  CLKBUF_X1 U2596 ( .A(n1212), .Z(n1501) );
  INV_X1 U2597 ( .A(n1824), .ZN(n1727) );
  AND2_X1 U2598 ( .A1(n1824), .A2(n1684), .ZN(n1683) );
  NAND2_X1 U2599 ( .A1(n1669), .A2(n1483), .ZN(n1688) );
  AND2_X1 U2604 ( .A1(n1374), .A2(RST), .ZN(n1506) );
  AND2_X1 U2605 ( .A1(n1374), .A2(RST), .ZN(n1507) );
  INV_X1 U2608 ( .A(n1557), .ZN(n1508) );
  OR2_X1 U2610 ( .A1(n1212), .A2(n1492), .ZN(n1511) );
  AOI22_X1 U2611 ( .A1(n639), .A2(\DP/RegLMD_out[10] ), .B1(n638), .B2(
        \DP/RegALU2_out[10] ), .ZN(n1212) );
  NOR2_X1 U2612 ( .A1(n1512), .A2(n1513), .ZN(n1515) );
  NAND3_X1 U2613 ( .A1(n1711), .A2(n1518), .A3(n1516), .ZN(n1512) );
  NOR2_X1 U2614 ( .A1(n1515), .A2(n1676), .ZN(n1675) );
  INV_X1 U2615 ( .A(n1517), .ZN(n1516) );
  NAND2_X1 U2616 ( .A1(n1673), .A2(n1672), .ZN(n1517) );
  NOR2_X1 U2617 ( .A1(n902), .A2(n900), .ZN(n1518) );
  NAND2_X2 U2618 ( .A1(n1610), .A2(n958), .ZN(\DP/RF_DATA[25] ) );
  NAND2_X1 U2619 ( .A1(n947), .A2(n1519), .ZN(\DP/RF_DATA[14] ) );
  OR2_X1 U2620 ( .A1(n1220), .A2(n1492), .ZN(n1519) );
  AOI21_X1 U2621 ( .B1(n639), .B2(\DP/RegLMD_out[14] ), .A(n1520), .ZN(n1220)
         );
  AND2_X1 U2622 ( .A1(\DP/RegALU2_out[14] ), .A2(n583), .ZN(n1520) );
  NAND2_X2 U2623 ( .A1(n1614), .A2(n953), .ZN(\DP/RF_DATA[20] ) );
  NAND2_X2 U2624 ( .A1(n1612), .A2(n961), .ZN(\DP/RF_DATA[28] ) );
  NAND2_X2 U2625 ( .A1(n1616), .A2(n965), .ZN(\DP/RF_DATA[31] ) );
  NAND2_X2 U2626 ( .A1(n964), .A2(n1522), .ZN(\DP/RF_DATA[30] ) );
  NAND2_X2 U2628 ( .A1(n956), .A2(n1523), .ZN(\DP/RF_DATA[23] ) );
  NAND2_X1 U2629 ( .A1(n1573), .A2(n1473), .ZN(n1575) );
  NAND2_X1 U2630 ( .A1(n1332), .A2(n1686), .ZN(n1634) );
  INV_X1 U2631 ( .A(n1726), .ZN(n1685) );
  NAND2_X1 U2632 ( .A1(n1685), .A2(n1683), .ZN(w_RF_RD1) );
  NOR2_X1 U2633 ( .A1(n1524), .A2(n1526), .ZN(n729) );
  OAI21_X1 U2634 ( .B1(n1525), .B2(n759), .A(n1531), .ZN(n1524) );
  AOI21_X1 U2635 ( .B1(n1527), .B2(n1530), .A(n1528), .ZN(n1525) );
  NOR2_X1 U2636 ( .A1(n1322), .A2(n724), .ZN(n1526) );
  AND2_X1 U2637 ( .A1(n722), .A2(n736), .ZN(n1529) );
  AOI21_X1 U2638 ( .B1(n758), .B2(n730), .A(n1658), .ZN(n1530) );
  NAND2_X1 U2639 ( .A1(n727), .A2(RST), .ZN(n1531) );
  NAND2_X1 U2640 ( .A1(n1476), .A2(n1532), .ZN(n1567) );
  NAND2_X1 U2642 ( .A1(n697), .A2(n656), .ZN(n1532) );
  NAND2_X1 U2643 ( .A1(n710), .A2(n1483), .ZN(n656) );
  NOR2_X1 U2644 ( .A1(n1690), .A2(n660), .ZN(n710) );
  INV_X1 U2645 ( .A(n645), .ZN(n714) );
  BUF_X2 U2646 ( .A(n1550), .Z(n1533) );
  AOI21_X1 U2647 ( .B1(n1535), .B2(n1534), .A(n1544), .ZN(\DP/FFDBRANCH/N3 )
         );
  NOR2_X1 U2648 ( .A1(\DP/FFDJL1/N3 ), .A2(\DP/FFDJREG/N3 ), .ZN(n1534) );
  NAND2_X1 U2649 ( .A1(n933), .A2(RST), .ZN(n1535) );
  AND2_X1 U2650 ( .A1(n1536), .A2(n1561), .ZN(n1559) );
  NOR2_X1 U2651 ( .A1(n1715), .A2(n1537), .ZN(n1536) );
  INV_X1 U2652 ( .A(n1560), .ZN(n1537) );
  BUF_X2 U2653 ( .A(n1327), .Z(n1538) );
  NAND2_X1 U2655 ( .A1(n703), .A2(n1591), .ZN(n1561) );
  BUF_X1 U2656 ( .A(n1350), .Z(n1539) );
  AND2_X2 U2657 ( .A1(n1813), .A2(n1541), .ZN(n1805) );
  AND2_X2 U2658 ( .A1(n1290), .A2(n1542), .ZN(n1541) );
  INV_X2 U2659 ( .A(n1806), .ZN(n1542) );
  BUF_X2 U2660 ( .A(n710), .Z(n1543) );
  NAND2_X1 U2663 ( .A1(n660), .A2(n586), .ZN(n1687) );
  INV_X1 U2664 ( .A(n660), .ZN(n1546) );
  CLKBUF_X3 U2665 ( .A(n1634), .Z(n1550) );
  BUF_X2 U2666 ( .A(n691), .Z(n1547) );
  NOR2_X2 U2669 ( .A1(n1550), .A2(n681), .ZN(n755) );
  NAND2_X2 U2670 ( .A1(n1550), .A2(RST), .ZN(n1645) );
  NOR2_X2 U2671 ( .A1(n1551), .A2(n662), .ZN(\CU/N59 ) );
  NAND2_X2 U2672 ( .A1(n1552), .A2(n1539), .ZN(n1551) );
  INV_X2 U2673 ( .A(n661), .ZN(n1552) );
  AOI22_X1 U2674 ( .A1(n695), .A2(n1543), .B1(n1556), .B2(n694), .ZN(n696) );
  INV_X1 U2675 ( .A(n1547), .ZN(n1556) );
  INV_X1 U2676 ( .A(IR_OUT[26]), .ZN(n1557) );
  INV_X2 U2677 ( .A(RST), .ZN(n1558) );
  NAND3_X1 U2678 ( .A1(n1332), .A2(n666), .A3(n1299), .ZN(n1039) );
  NAND2_X1 U2679 ( .A1(n1559), .A2(n1482), .ZN(n1713) );
  INV_X1 U2680 ( .A(n1565), .ZN(n1560) );
  INV_X2 U2683 ( .A(n586), .ZN(n1564) );
  INV_X2 U2684 ( .A(n1714), .ZN(n1565) );
  NOR2_X1 U2685 ( .A1(n1566), .A2(n1568), .ZN(n1723) );
  NAND4_X1 U2686 ( .A1(n1567), .A2(n1569), .A3(n1582), .A4(n1042), .ZN(n1566)
         );
  NAND2_X1 U2687 ( .A1(n1575), .A2(n1316), .ZN(n1568) );
  NAND2_X1 U2688 ( .A1(n1570), .A2(n653), .ZN(n739) );
  NAND3_X1 U2689 ( .A1(n1041), .A2(n688), .A3(n1571), .ZN(n1570) );
  NAND2_X1 U2690 ( .A1(n1577), .A2(n1578), .ZN(n1582) );
  INV_X1 U2691 ( .A(IR_OUT[26]), .ZN(n1571) );
  INV_X1 U2692 ( .A(n1355), .ZN(n1572) );
  CLKBUF_X1 U2693 ( .A(w_RF_RD2), .Z(n1574) );
  NOR2_X1 U2694 ( .A1(n1579), .A2(n665), .ZN(n1577) );
  INV_X2 U2695 ( .A(n1581), .ZN(n1578) );
  NAND2_X2 U2696 ( .A1(n1192), .A2(n1583), .ZN(n1097) );
  NOR2_X2 U2697 ( .A1(n1680), .A2(n1584), .ZN(n1583) );
  NAND2_X2 U2698 ( .A1(\DP/NPC1[6] ), .A2(IROM_ADDR[5]), .ZN(n1584) );
  AND2_X2 U2699 ( .A1(n1192), .A2(IROM_ADDR[5]), .ZN(n1198) );
  NAND2_X2 U2700 ( .A1(n1198), .A2(\DP/NPC1[6] ), .ZN(n1197) );
  NAND2_X2 U2702 ( .A1(n1544), .A2(IR_OUT[2]), .ZN(n1053) );
  NAND2_X2 U2703 ( .A1(n1589), .A2(n1588), .ZN(n1587) );
  INV_X2 U2704 ( .A(IR_OUT[0]), .ZN(n1588) );
  INV_X2 U2705 ( .A(IR_OUT[2]), .ZN(n1589) );
  INV_X2 U2707 ( .A(n1549), .ZN(n754) );
  INV_X1 U2708 ( .A(n1483), .ZN(n1591) );
  INV_X2 U2709 ( .A(n62), .ZN(n1592) );
  INV_X1 U2710 ( .A(n1469), .ZN(n738) );
  NOR2_X1 U2711 ( .A1(n1594), .A2(n675), .ZN(n935) );
  NAND2_X1 U2712 ( .A1(n1595), .A2(n1596), .ZN(n1594) );
  NOR2_X1 U2713 ( .A1(w_RF_RD2), .A2(n1374), .ZN(n1595) );
  INV_X1 U2714 ( .A(n676), .ZN(n1596) );
  NAND2_X1 U2715 ( .A1(n1500), .A2(n1043), .ZN(n675) );
  INV_X2 U2716 ( .A(n1598), .ZN(n941) );
  NAND2_X2 U2717 ( .A1(n35), .A2(n73), .ZN(n1599) );
  NAND4_X2 U2718 ( .A1(n1606), .A2(n1604), .A3(n1603), .A4(n1602), .ZN(n1601)
         );
  NAND2_X2 U2719 ( .A1(n1204), .A2(\DP/RD2[1] ), .ZN(n1602) );
  INV_X2 U2720 ( .A(n1605), .ZN(n1604) );
  INV_X2 U2721 ( .A(n1607), .ZN(n1606) );
  OR2_X2 U2722 ( .A1(n37), .A2(n72), .ZN(n1608) );
  OR2_X2 U2723 ( .A1(n36), .A2(n598), .ZN(n1609) );
  INV_X1 U2724 ( .A(n1611), .ZN(n1610) );
  NOR2_X1 U2725 ( .A1(n1245), .A2(\DP/JL2 ), .ZN(n1611) );
  INV_X1 U2726 ( .A(n1613), .ZN(n1612) );
  NOR2_X1 U2727 ( .A1(n1251), .A2(\DP/JL2 ), .ZN(n1613) );
  INV_X1 U2728 ( .A(n1615), .ZN(n1614) );
  NOR2_X1 U2729 ( .A1(n1235), .A2(\DP/JL2 ), .ZN(n1615) );
  INV_X1 U2730 ( .A(n1617), .ZN(n1616) );
  NOR2_X1 U2731 ( .A1(n1260), .A2(\DP/JL2 ), .ZN(n1617) );
  CLKBUF_X1 U2732 ( .A(n1632), .Z(n1618) );
  AND2_X2 U2733 ( .A1(n1621), .A2(n1619), .ZN(n1632) );
  INV_X2 U2734 ( .A(n1633), .ZN(n1619) );
  AND2_X1 U2735 ( .A1(n1622), .A2(n1621), .ZN(n1620) );
  NAND2_X1 U2736 ( .A1(n639), .A2(\DP/RegLMD_out[2] ), .ZN(n1621) );
  NOR2_X1 U2737 ( .A1(n1623), .A2(n1633), .ZN(n1622) );
  INV_X1 U2738 ( .A(n1275), .ZN(n1623) );
  OAI22_X2 U2739 ( .A1(n1618), .A2(n1278), .B1(n613), .B2(n1277), .ZN(
        DRAM_DATA_OUT[2]) );
  NAND2_X2 U2740 ( .A1(n876), .A2(n1624), .ZN(\DP/B[2] ) );
  NOR2_X2 U2741 ( .A1(n1626), .A2(n1625), .ZN(n1624) );
  NOR2_X2 U2742 ( .A1(n1618), .A2(n897), .ZN(n1625) );
  INV_X2 U2743 ( .A(n875), .ZN(n1626) );
  NAND2_X2 U2744 ( .A1(n1004), .A2(n1627), .ZN(\DP/RegA1/N5 ) );
  INV_X2 U2745 ( .A(n1628), .ZN(n1627) );
  NOR2_X2 U2746 ( .A1(n630), .A2(n1618), .ZN(n1628) );
  NAND2_X2 U2747 ( .A1(n811), .A2(n1629), .ZN(\DP/A[2] ) );
  NOR2_X2 U2748 ( .A1(n1631), .A2(n1630), .ZN(n1629) );
  INV_X2 U2749 ( .A(n810), .ZN(n1630) );
  NOR2_X2 U2750 ( .A1(n621), .A2(n1618), .ZN(n1631) );
  AND2_X1 U2751 ( .A1(\DP/RegALU2_out[2] ), .A2(n583), .ZN(n1633) );
  OAI21_X2 U2752 ( .B1(n190), .B2(n1533), .A(n1635), .ZN(\DP/RegRD1/N3 ) );
  INV_X2 U2753 ( .A(n1636), .ZN(n1635) );
  OAI21_X2 U2754 ( .B1(n188), .B2(n1533), .A(n1637), .ZN(\DP/RegRD1/N4 ) );
  INV_X2 U2755 ( .A(n1638), .ZN(n1637) );
  NOR2_X2 U2756 ( .A1(n1645), .A2(n1452), .ZN(n1638) );
  OAI21_X2 U2757 ( .B1(n186), .B2(n1533), .A(n1639), .ZN(\DP/RegRD1/N5 ) );
  INV_X2 U2758 ( .A(n1640), .ZN(n1639) );
  OAI21_X2 U2759 ( .B1(n184), .B2(n1533), .A(n1641), .ZN(\DP/RegRD1/N6 ) );
  INV_X2 U2760 ( .A(n1642), .ZN(n1641) );
  OAI21_X2 U2761 ( .B1(n181), .B2(n1533), .A(n1643), .ZN(\DP/RegRD1/N7 ) );
  INV_X2 U2762 ( .A(n1644), .ZN(n1643) );
  NAND2_X2 U2763 ( .A1(n969), .A2(n1646), .ZN(\DP/RF_DATA[6] ) );
  NAND2_X2 U2764 ( .A1(n1010), .A2(n1647), .ZN(\DP/RegA1/N9 ) );
  INV_X2 U2765 ( .A(n1648), .ZN(n1647) );
  NAND2_X2 U2766 ( .A1(n822), .A2(n1649), .ZN(\DP/A[6] ) );
  NOR2_X2 U2767 ( .A1(n1651), .A2(n1650), .ZN(n1649) );
  INV_X2 U2768 ( .A(n823), .ZN(n1651) );
  NAND2_X2 U2769 ( .A1(n887), .A2(n1652), .ZN(\DP/B[6] ) );
  NOR2_X2 U2770 ( .A1(n1656), .A2(n1653), .ZN(n1652) );
  INV_X2 U2771 ( .A(n886), .ZN(n1656) );
  INV_X1 U2772 ( .A(n1465), .ZN(n718) );
  NAND2_X1 U2773 ( .A1(n1495), .A2(IR_OUT[1]), .ZN(n1666) );
  CLKBUF_X1 U2774 ( .A(n1465), .Z(n1657) );
  CLKBUF_X1 U2775 ( .A(n718), .Z(n1658) );
  AND2_X2 U2776 ( .A1(n1658), .A2(n1659), .ZN(\DP/RegIMM/N4 ) );
  INV_X2 U2777 ( .A(n641), .ZN(n1659) );
  INV_X2 U2779 ( .A(n1661), .ZN(n1660) );
  INV_X2 U2780 ( .A(n1663), .ZN(n1662) );
  NAND3_X1 U2781 ( .A1(n737), .A2(\DP/RegIMM/N3 ), .A3(n1657), .ZN(n1663) );
  NAND2_X1 U2782 ( .A1(n677), .A2(n1315), .ZN(n747) );
  NOR2_X1 U2783 ( .A1(n1665), .A2(n1658), .ZN(n1664) );
  INV_X1 U2784 ( .A(n732), .ZN(n1665) );
  INV_X2 U2785 ( .A(n1493), .ZN(n638) );
  NAND2_X1 U2786 ( .A1(n1670), .A2(n1674), .ZN(n1671) );
  NAND3_X1 U2787 ( .A1(n903), .A2(n1300), .A3(n1711), .ZN(n1670) );
  NAND2_X1 U2788 ( .A1(n1675), .A2(n1671), .ZN(n933) );
  INV_X1 U2789 ( .A(w_JUMP_EQ), .ZN(n1672) );
  INV_X1 U2790 ( .A(n1691), .ZN(n1673) );
  AND2_X2 U2791 ( .A1(n1710), .A2(w_JUMP_EQ), .ZN(n1674) );
  OR2_X2 U2792 ( .A1(n1710), .A2(w_JUMP_EQ), .ZN(n1678) );
  NOR2_X2 U2794 ( .A1(n1197), .A2(n1682), .ZN(n1094) );
  NAND2_X2 U2795 ( .A1(n1681), .A2(IROM_ADDR[8]), .ZN(n1680) );
  INV_X2 U2796 ( .A(n1682), .ZN(n1681) );
  INV_X1 U2797 ( .A(n1197), .ZN(n1091) );
  INV_X2 U2798 ( .A(IROM_ADDR[7]), .ZN(n1682) );
  INV_X1 U2799 ( .A(n660), .ZN(n697) );
  NOR2_X1 U2800 ( .A1(n1688), .A2(n1687), .ZN(n1686) );
  INV_X1 U2801 ( .A(n62), .ZN(n1689) );
  INV_X2 U2802 ( .A(n1543), .ZN(n690) );
  INV_X2 U2803 ( .A(IR_OUT[26]), .ZN(n1690) );
  NOR2_X2 U2804 ( .A1(n1104), .A2(n1732), .ZN(n1112) );
  OR2_X2 U2805 ( .A1(n1097), .A2(n1719), .ZN(n1104) );
  INV_X1 U2806 ( .A(n1708), .ZN(n1691) );
  OAI21_X2 U2807 ( .B1(n1265), .B2(n1488), .A(n970), .ZN(\DP/RF_DATA[8] ) );
  INV_X2 U2808 ( .A(n1538), .ZN(n661) );
  INV_X2 U2809 ( .A(IR_OUT[31]), .ZN(n1693) );
  INV_X2 U2810 ( .A(IR_OUT[29]), .ZN(n1694) );
  NOR2_X2 U2811 ( .A1(n1696), .A2(IR_OUT[31]), .ZN(n1695) );
  INV_X2 U2812 ( .A(IR_OUT[29]), .ZN(n1696) );
  NOR2_X1 U2813 ( .A1(n1104), .A2(n1700), .ZN(n1140) );
  NOR2_X2 U2814 ( .A1(n1104), .A2(n1698), .ZN(n1697) );
  NAND2_X2 U2815 ( .A1(n1702), .A2(n1699), .ZN(n1698) );
  NOR2_X2 U2816 ( .A1(n1706), .A2(n1703), .ZN(n1702) );
  INV_X2 U2817 ( .A(n1786), .ZN(n1705) );
  INV_X2 U2818 ( .A(n1803), .ZN(n1706) );
  INV_X2 U2819 ( .A(n1125), .ZN(n1126) );
  INV_X2 U2820 ( .A(n974), .ZN(n1710) );
  CLKBUF_X1 U2821 ( .A(n666), .Z(n1712) );
  INV_X2 U2822 ( .A(n1712), .ZN(n663) );
  NAND4_X1 U2823 ( .A1(n1713), .A2(n1461), .A3(n1757), .A4(n1758), .ZN(n1756)
         );
  INV_X1 U2824 ( .A(n62), .ZN(n1714) );
  NOR2_X1 U2825 ( .A1(n1546), .A2(n1328), .ZN(n1715) );
  INV_X2 U2826 ( .A(n1719), .ZN(n1717) );
  INV_X2 U2827 ( .A(n1730), .ZN(n1718) );
  NOR2_X2 U2828 ( .A1(n1097), .A2(n1721), .ZN(n1101) );
  NAND2_X2 U2829 ( .A1(n1720), .A2(IROM_ADDR[10]), .ZN(n1719) );
  INV_X2 U2830 ( .A(n1721), .ZN(n1720) );
  INV_X1 U2831 ( .A(n1097), .ZN(n1098) );
  INV_X2 U2832 ( .A(IROM_ADDR[9]), .ZN(n1721) );
  NOR2_X2 U2834 ( .A1(n1726), .A2(n1727), .ZN(n972) );
  NAND2_X2 U2835 ( .A1(n1731), .A2(n1738), .ZN(n1730) );
  NAND2_X2 U2836 ( .A1(n1733), .A2(w_PC_OUT[12]), .ZN(n1732) );
  INV_X1 U2837 ( .A(n1104), .ZN(n1105) );
  NOR2_X2 U2838 ( .A1(n1759), .A2(n1737), .ZN(n1736) );
  INV_X2 U2839 ( .A(n1738), .ZN(n1737) );
  AND2_X2 U2840 ( .A1(\DP/NPC1[13] ), .A2(\DP/NPC1[14] ), .ZN(n1738) );
  NOR2_X1 U2841 ( .A1(n1118), .A2(n1761), .ZN(n1122) );
  OAI21_X1 U2842 ( .B1(n1118), .B2(n1739), .A(n1741), .ZN(n1798) );
  INV_X2 U2843 ( .A(n1744), .ZN(n1741) );
  INV_X1 U2844 ( .A(n1799), .ZN(n1744) );
  NOR2_X1 U2845 ( .A1(n1118), .A2(n1747), .ZN(n1809) );
  NOR2_X1 U2846 ( .A1(n1118), .A2(n1746), .ZN(n1133) );
  INV_X2 U2847 ( .A(n1748), .ZN(n1746) );
  NAND2_X2 U2848 ( .A1(n1765), .A2(n1748), .ZN(n1747) );
  NOR2_X2 U2849 ( .A1(n1749), .A2(n1754), .ZN(n1748) );
  NAND2_X2 U2850 ( .A1(n1751), .A2(n1750), .ZN(n1749) );
  INV_X2 U2851 ( .A(n1745), .ZN(n1751) );
  NAND2_X2 U2852 ( .A1(n1766), .A2(n1753), .ZN(n1752) );
  INV_X2 U2853 ( .A(n1754), .ZN(n1753) );
  INV_X2 U2854 ( .A(n1764), .ZN(n1754) );
  NAND2_X1 U2855 ( .A1(n1474), .A2(n1538), .ZN(n1757) );
  AND2_X1 U2856 ( .A1(n702), .A2(n750), .ZN(n1758) );
  AND2_X2 U2857 ( .A1(n1785), .A2(n1763), .ZN(n1762) );
  AND2_X2 U2858 ( .A1(n1768), .A2(n1764), .ZN(n1763) );
  AND2_X2 U2859 ( .A1(w_PC_OUT[17]), .A2(w_PC_OUT[18]), .ZN(n1764) );
  AND2_X2 U2860 ( .A1(n1778), .A2(n1766), .ZN(n1765) );
  INV_X2 U2861 ( .A(n1767), .ZN(n1766) );
  NAND2_X2 U2862 ( .A1(n1768), .A2(n1788), .ZN(n1767) );
  AND2_X2 U2863 ( .A1(n1133), .A2(\DP/NPC1[19] ), .ZN(n1136) );
  AND2_X2 U2864 ( .A1(\DP/NPC1[19] ), .A2(\DP/NPC1[20] ), .ZN(n1768) );
  INV_X2 U2865 ( .A(n1140), .ZN(n1139) );
  OAI21_X2 U2866 ( .B1(n1140), .B2(n1773), .A(n1769), .ZN(n1164) );
  AND2_X2 U2867 ( .A1(n1771), .A2(n1770), .ZN(n1769) );
  OR2_X2 U2868 ( .A1(n1773), .A2(n1788), .ZN(n1770) );
  INV_X2 U2869 ( .A(n1772), .ZN(n1771) );
  OAI21_X2 U2870 ( .B1(n1789), .B2(n1773), .A(n634), .ZN(n1772) );
  INV_X2 U2871 ( .A(n1774), .ZN(n1773) );
  INV_X1 U2872 ( .A(w_PC_OUT[27]), .ZN(n1774) );
  OAI211_X1 U2873 ( .C1(n1157), .C2(\DP/NPC1[26] ), .A(n633), .B(n1161), .ZN(
        n1158) );
  AND2_X2 U2874 ( .A1(n1791), .A2(n1788), .ZN(n1775) );
  NOR2_X1 U2875 ( .A1(n1153), .A2(n1812), .ZN(n1157) );
  OR2_X1 U2876 ( .A1(n1809), .A2(n1792), .ZN(n1780) );
  NOR2_X2 U2877 ( .A1(n1782), .A2(n1777), .ZN(n1776) );
  INV_X2 U2878 ( .A(n1791), .ZN(n1777) );
  NOR2_X2 U2879 ( .A1(n1810), .A2(n1779), .ZN(n1778) );
  INV_X2 U2880 ( .A(n1791), .ZN(n1779) );
  OAI21_X1 U2881 ( .B1(n1781), .B2(n1780), .A(n1167), .ZN(\PC/N31 ) );
  NOR2_X1 U2882 ( .A1(n1165), .A2(w_PC_OUT[28]), .ZN(n1781) );
  NAND2_X1 U2883 ( .A1(n1784), .A2(n1783), .ZN(n1782) );
  INV_X1 U2884 ( .A(n1793), .ZN(n1783) );
  INV_X1 U2885 ( .A(n1811), .ZN(n1784) );
  AND2_X2 U2886 ( .A1(n1805), .A2(n1786), .ZN(n1785) );
  INV_X2 U2887 ( .A(n1787), .ZN(n1786) );
  NAND2_X2 U2888 ( .A1(n1788), .A2(\DP/NPC1[23] ), .ZN(n1787) );
  AND2_X2 U2889 ( .A1(n1140), .A2(w_PC_OUT[21]), .ZN(n1143) );
  AND2_X2 U2890 ( .A1(w_PC_OUT[21]), .A2(\DP/NPC1[22] ), .ZN(n1788) );
  INV_X2 U2891 ( .A(n1791), .ZN(n1790) );
  AND2_X2 U2892 ( .A1(\DP/NPC1[23] ), .A2(w_PC_OUT[24]), .ZN(n1791) );
  INV_X1 U2893 ( .A(n633), .ZN(n1792) );
  NOR2_X1 U2894 ( .A1(n1358), .A2(n1146), .ZN(n1172) );
  OAI21_X1 U2895 ( .B1(n1161), .B2(n1797), .A(n1794), .ZN(\PC/N33 ) );
  INV_X2 U2896 ( .A(w_PC_OUT[30]), .ZN(n1796) );
  INV_X1 U2897 ( .A(n591), .ZN(n1799) );
  OAI211_X1 U2898 ( .C1(n1150), .C2(n1807), .A(n1802), .B(n1801), .ZN(n1177)
         );
  OR2_X1 U2899 ( .A1(n1805), .A2(n1807), .ZN(n1801) );
  INV_X1 U2900 ( .A(n1804), .ZN(n1803) );
  NAND2_X1 U2901 ( .A1(n1805), .A2(n1807), .ZN(n1804) );
  INV_X2 U2902 ( .A(w_PC_OUT[24]), .ZN(n1806) );
  INV_X2 U2903 ( .A(n1808), .ZN(n1807) );
  INV_X2 U2904 ( .A(\DP/NPC1[31] ), .ZN(n1808) );
  OAI21_X2 U2905 ( .B1(n1809), .B2(\DP/NPC1[29] ), .A(n634), .ZN(n1171) );
  INV_X1 U2906 ( .A(n1153), .ZN(n1154) );
  INV_X1 U2907 ( .A(n1188), .ZN(n1192) );
  NAND2_X1 U2908 ( .A1(n1818), .A2(n1351), .ZN(n1188) );
  NOR2_X2 U2909 ( .A1(n1820), .A2(n1819), .ZN(n1818) );
  INV_X2 U2910 ( .A(\DP/NPC1[4] ), .ZN(n1819) );
  INV_X1 U2911 ( .A(\DP/NPC1[3] ), .ZN(n1820) );
  DFF_X1 \DP/RegLMD/DOUT_reg[21]  ( .D(n1840), .CK(\DP/RegLMD/net7068 ), .Q(
        \DP/RegLMD_out[21] ) );
  DFF_X1 \PC/DOUT_reg[5]  ( .D(\PC/N8 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IROM_ADDR[5]) );
  DFF_X1 \PC/DOUT_reg[0]  ( .D(\PC/N3 ), .CK(\DP/RegNPC/net7068 ), .Q(
        IROM_ADDR[0]) );
  AND2_X2 U2654 ( .A1(n1328), .A2(n62), .ZN(n1563) );
  AND3_X1 U1191 ( .A1(n1666), .A2(n1054), .A3(n1586), .ZN(n1821) );
  CLKBUF_X1 U1231 ( .A(n1048), .Z(n1822) );
  CLKBUF_X1 U1274 ( .A(n1330), .Z(n1823) );
  CLKBUF_X1 U1353 ( .A(n1041), .Z(n1330) );
  NOR2_X1 U1358 ( .A1(n716), .A2(n1660), .ZN(n721) );
  INV_X1 U1370 ( .A(n1293), .ZN(n1824) );
  NOR2_X1 U1464 ( .A1(n740), .A2(n1343), .ZN(n1499) );
  NOR2_X1 U1627 ( .A1(n1294), .A2(n1293), .ZN(n1825) );
  CLKBUF_X1 U2600 ( .A(n1476), .Z(n1829) );
  AND2_X1 U2601 ( .A1(n1476), .A2(n1532), .ZN(n1830) );
  AND2_X1 U2914 ( .A1(RST), .A2(\DP/RD1[0] ), .ZN(n1839) );
  INV_X1 U2915 ( .A(n1077), .ZN(n1840) );
  BUF_X1 U1361 ( .A(n1495), .Z(n1349) );
  DFF_X1 \DP/RegNPC/DOUT_reg[1]  ( .D(\PC/N4 ), .CK(\DP/RegNPC/net7068 ), .Q(
        \DP/NPC1[1] ) );
  DFF_X1 \PC/DOUT_reg[21]  ( .D(\PC/N24 ), .CK(\DP/RegNPC/net7068 ), .Q(
        w_PC_OUT[21]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[20]  ( .D(\PC/N23 ), .CK(\DP/RegNPC/net7068 ), 
        .Q(\DP/NPC1[20] ) );
  DFF_X1 \DP/RegFB/DOUT_reg[2]  ( .D(n1846), .CK(\DP/RegNPC1/net7068 ), .QN(
        n75) );
  DFF_X1 \DP/RegIMM/DOUT_reg[16]  ( .D(\DP/RegIMM/N19 ), .CK(
        \DP/RegIMM/net7068 ), .Q(\DP/RegIMM_out[16] ) );
  DFF_X1 \DP/RegRD3/DOUT_reg[1]  ( .D(\DP/RegRD3/N4 ), .CK(\DP/RegRD3/net7086 ), .Q(\DP/RD3[1] ) );
  DFF_X1 \DP/RegRD3/DOUT_reg[0]  ( .D(\DP/RegRD3/N3 ), .CK(\DP/RegRD3/net7086 ), .Q(\DP/RD3[0] ) );
  DFF_X1 \CU/cw3_reg[0]  ( .D(\CU/N79 ), .CK(CLK), .Q(w_RF_WE) );
  DFF_X1 \DP/RegRD3/DOUT_reg[3]  ( .D(\DP/RegRD3/N6 ), .CK(\DP/RegRD3/net7086 ), .Q(\DP/RD3[3] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[31]  ( .D(\DP/RegNPC3/N34 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[31] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[30]  ( .D(\DP/RegNPC3/N33 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[30] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[29]  ( .D(\DP/RegNPC3/N32 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[29] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[28]  ( .D(\DP/RegNPC3/N31 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[28] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[27]  ( .D(\DP/RegNPC3/N30 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[27] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[26]  ( .D(\DP/RegNPC3/N29 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[26] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[25]  ( .D(\DP/RegNPC3/N28 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[25] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[24]  ( .D(\DP/RegNPC3/N27 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[24] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[23]  ( .D(\DP/RegNPC3/N26 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[23] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[22]  ( .D(\DP/RegNPC3/N25 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[22] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[21]  ( .D(\DP/RegNPC3/N24 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[21] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[20]  ( .D(\DP/RegNPC3/N23 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[20] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[19]  ( .D(\DP/RegNPC3/N22 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[19] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[18]  ( .D(\DP/RegNPC3/N21 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[18] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[17]  ( .D(\DP/RegNPC3/N20 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[17] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[16]  ( .D(\DP/RegNPC3/N19 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[16] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[15]  ( .D(\DP/RegNPC3/N18 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[15] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[14]  ( .D(\DP/RegNPC3/N17 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[14] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[13]  ( .D(\DP/RegNPC3/N16 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[13] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[12]  ( .D(\DP/RegNPC3/N15 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[12] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[11]  ( .D(\DP/RegNPC3/N14 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[11] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[10]  ( .D(\DP/RegNPC3/N13 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[10] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[9]  ( .D(\DP/RegNPC3/N12 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[9] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[8]  ( .D(\DP/RegNPC3/N11 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[8] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[7]  ( .D(\DP/RegNPC3/N10 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[7] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[6]  ( .D(\DP/RegNPC3/N9 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[6] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[5]  ( .D(\DP/RegNPC3/N8 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[5] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[4]  ( .D(\DP/RegNPC3/N7 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[4] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[3]  ( .D(\DP/RegNPC3/N6 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[3] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[2]  ( .D(\DP/RegNPC3/N5 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[2] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[1]  ( .D(\DP/RegNPC3/N4 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[1] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[0]  ( .D(\DP/RegNPC3/N3 ), .CK(
        \DP/RegNPC3/net7068 ), .Q(\DP/NPC_out[0] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[30]  ( .D(\DP/RegNPC1/N33 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[30] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[28]  ( .D(\DP/RegNPC1/N31 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[28] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[27]  ( .D(\DP/RegNPC1/N30 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[27] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[25]  ( .D(\DP/RegNPC1/N28 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[25] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[24]  ( .D(\DP/RegNPC1/N27 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[24] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[21]  ( .D(\DP/RegNPC1/N24 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[21] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[18]  ( .D(\DP/RegNPC1/N21 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[18] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[17]  ( .D(\DP/RegNPC1/N20 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[17] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[12]  ( .D(\DP/RegNPC1/N15 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[12] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[11]  ( .D(\DP/RegNPC1/N14 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[11] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[10]  ( .D(\DP/RegNPC1/N13 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[10] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[9]  ( .D(\DP/RegNPC1/N12 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[9] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[8]  ( .D(\DP/RegNPC1/N11 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[8] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[7]  ( .D(\DP/RegNPC1/N10 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[7] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[5]  ( .D(\DP/RegNPC1/N8 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[5] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[0]  ( .D(\DP/RegNPC1/N3 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[0] ) );
  DFF_X1 \CU/cw3_reg[2]  ( .D(\CU/N81 ), .CK(CLK), .QN(n1289) );
  DFF_X1 \CU/cw2_reg[14]  ( .D(\CU/N78 ), .CK(CLK), .Q(DRAM_EN) );
  DFF_X1 \CU/cw2_reg[13]  ( .D(\CU/N77 ), .CK(CLK), .Q(DRAM_RW) );
  DFF_X1 \CU/cw2_reg[9]  ( .D(\CU/N73 ), .CK(CLK), .Q(w_SIGN_LD) );
  DFF_X1 \CU/cw2_reg[8]  ( .D(\CU/N72 ), .CK(CLK), .Q(w_LOAD_SIZE[2]) );
  DFF_X1 \CU/cw2_reg[5]  ( .D(\CU/N69 ), .CK(CLK), .Q(w_RegALU2_LATCH_EN) );
  DFF_X1 \CU/cw2_reg[4]  ( .D(\CU/N68 ), .CK(CLK), .Q(w_RegLMD_LATCH_EN) );
  DFF_X1 \CU/cw2_reg[3]  ( .D(\CU/N67 ), .CK(CLK), .Q(w_RegRD3_LATCH_EN) );
  DFF_X1 \CU/cw2_reg[1]  ( .D(\CU/N65 ), .CK(CLK), .Q(\CU/cw2[1] ) );
  DFF_X1 \DP/RegRD3/DOUT_reg[2]  ( .D(\DP/RegRD3/N5 ), .CK(\DP/RegRD3/net7086 ), .Q(\DP/RD3[2] ) );
  DFF_X1 \DP/FFDJREG/Q_reg  ( .D(\DP/FFDJREG/N3 ), .CK(\DP/RegA1/net7068 ), 
        .Q(\DP/JREG ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[26]  ( .D(\DP/RegNPC1/N29 ), .CK(
        \DP/RegNPC1/net7068 ), .Q(\DP/NPC2[26] ) );
  SDFF_X1 \CU/JUMP2_reg  ( .D(1'b0), .SI(n1510), .SE(RST), .CK(CLK), .Q(
        \CU/JUMP2 ), .QN(n1667) );
  NAND2_X1 U1234 ( .A1(n1495), .A2(IR_OUT[29]), .ZN(n1590) );
  OR2_X1 U1269 ( .A1(n704), .A2(n1564), .ZN(n1851) );
  AND2_X2 U1369 ( .A1(n1667), .A2(IR_OUT[28]), .ZN(n1353) );
  NAND4_X1 U1503 ( .A1(n1667), .A2(n1668), .A3(IR_OUT[28]), .A4(n1728), .ZN(
        n1484) );
  BUF_X1 U1506 ( .A(n1575), .Z(n1355) );
  OAI22_X1 U1513 ( .A1(n692), .A2(n1547), .B1(n690), .B2(n1432), .ZN(n706) );
  BUF_X1 U1792 ( .A(n687), .Z(n1843) );
  INV_X1 U1793 ( .A(n1332), .ZN(n1844) );
  AND2_X1 U2228 ( .A1(RST), .A2(n1038), .ZN(n1846) );
  AND3_X1 U2241 ( .A1(n1847), .A2(n1041), .A3(n1563), .ZN(n648) );
  AND2_X2 U2249 ( .A1(n1495), .A2(n1695), .ZN(n1041) );
  NAND2_X1 U2270 ( .A1(n691), .A2(n703), .ZN(n1847) );
  NAND2_X1 U2515 ( .A1(n660), .A2(IR_OUT[26]), .ZN(n703) );
  NAND2_X1 U2548 ( .A1(n1848), .A2(n1723), .ZN(\DP/RF_EN ) );
  NOR2_X1 U2551 ( .A1(n1849), .A2(n1756), .ZN(n1848) );
  OR3_X2 U2584 ( .A1(n752), .A2(n1850), .A3(n648), .ZN(n1849) );
  NOR2_X1 U2593 ( .A1(n665), .A2(n1851), .ZN(n1850) );
  NAND3_X1 U2606 ( .A1(n691), .A2(n1482), .A3(n666), .ZN(n1042) );
  AND2_X2 U2609 ( .A1(n1349), .A2(n1852), .ZN(n1482) );
  AND2_X2 U2641 ( .A1(IR_OUT[31]), .A2(IR_OUT[29]), .ZN(n1852) );
  NAND2_X2 U2535 ( .A1(n1576), .A2(n1729), .ZN(n660) );
  INV_X2 U1389 ( .A(n652), .ZN(n704) );
  OR2_X1 U1236 ( .A1(n1508), .A2(n660), .ZN(n691) );
  CLKBUF_X1 U1256 ( .A(n1495), .Z(n1544) );
  NAND2_X1 U1261 ( .A1(n1495), .A2(IR_OUT[31]), .ZN(n645) );
  NOR2_X1 U1283 ( .A1(n665), .A2(n704), .ZN(n687) );
  AND2_X2 U1806 ( .A1(n1495), .A2(n1692), .ZN(n665) );
  AND2_X1 U2534 ( .A1(RST), .A2(\CU/JUMP2 ), .ZN(n1853) );
  AND2_X4 U2579 ( .A1(n1854), .A2(n1668), .ZN(n1495) );
  NOR2_X1 U2602 ( .A1(n1510), .A2(\CU/JUMP2 ), .ZN(n1854) );
  DFF_X1 \DP/RegRD2/DOUT_reg[1]  ( .D(\DP/RegRD2/N4 ), .CK(\DP/RegRD2/net7086 ), .Q(\DP/RD2[1] ), .QN(n594) );
  DFF_X1 \DP/RegRD2/DOUT_reg[4]  ( .D(\DP/RegRD2/N7 ), .CK(\DP/RegRD2/net7086 ), .Q(n593), .QN(n73) );
  DFF_X1 \DP/RegRD2/DOUT_reg[2]  ( .D(\DP/RegRD2/N5 ), .CK(\DP/RegRD2/net7086 ), .Q(\DP/RD2[2] ), .QN(n585) );
  DFF_X1 \CU/cw3_reg[1]  ( .D(\CU/N80 ), .CK(CLK), .Q(w_MuxWB_SEL), .QN(n583)
         );
  DFF_X1 \CU/cw2_reg[11]  ( .D(\CU/N75 ), .CK(CLK), .Q(w_STORE_SIZE[1]), .QN(
        n603) );
  DFF_X1 \CU/cw2_reg[10]  ( .D(\CU/N74 ), .CK(CLK), .Q(w_STORE_SIZE[0]), .QN(
        n606) );
  DFF_X1 \CU/cw2_reg[7]  ( .D(\CU/N71 ), .CK(CLK), .Q(w_LOAD_SIZE[1]), .QN(
        n587) );
  DFF_X1 \CU/cw2_reg[6]  ( .D(\CU/N70 ), .CK(CLK), .Q(n602), .QN(n53) );
  DFF_X1 \CU/JUMP3_reg  ( .D(n1853), .CK(CLK), .Q(\CU/JUMP3 ), .QN(n1668) );
  DFF_X1 \DP/RegME/DOUT_reg[7]  ( .D(\DP/RegME/N10 ), .CK(\DP/RegME/net7068 ), 
        .Q(\DP/RegME_out[7] ), .QN(n610) );
  DFF_X1 \DP/RegRD2/DOUT_reg[0]  ( .D(n1839), .CK(\DP/RegRD2/net7086 ), .Q(
        \DP/RD2[0] ), .QN(n598) );
  DFF_X1 \DP/RegRD2/DOUT_reg[3]  ( .D(\DP/RegRD2/N6 ), .CK(\DP/RegRD2/net7086 ), .Q(n584), .QN(n72) );
  DFF_X1 \CU/JUMP1_reg  ( .D(\CU/N82 ), .CK(CLK), .Q(n1510), .QN(n1728) );
  DFF_X1 \DP/RegRD1/DOUT_reg[4]  ( .D(\DP/RegRD1/N7 ), .CK(\DP/RegRD1/net7086 ), .Q(\DP/RD1[4] ), .QN(n596) );
  DFF_X1 \DP/RegRD1/DOUT_reg[2]  ( .D(\DP/RegRD1/N5 ), .CK(\DP/RegRD1/net7086 ), .Q(\DP/RD1[2] ), .QN(n597) );
  DFF_X1 \DP/RegRD1/DOUT_reg[1]  ( .D(\DP/RegRD1/N4 ), .CK(\DP/RegRD1/net7086 ), .Q(\DP/RD1[1] ), .QN(n599) );
  DFF_X1 \DP/RegALU1/DOUT_reg[26]  ( .D(\DP/RegALU1/N29 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[26] ), .QN(n1386) );
  DFF_X1 \DP/RegALU1/DOUT_reg[3]  ( .D(\DP/RegALU1/N6 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[3]) );
  DFF_X1 \CU/cw1_reg[21]  ( .D(\CU/N61 ), .CK(CLK), .Q(w_MuxB_SEL), .QN(n609)
         );
  DFF_X1 \DP/FFDFD/Q_reg  ( .D(\DP/FFDFD/N3 ), .CK(\DP/RegNPC1/net7068 ), .Q(
        \DP/FwdD ), .QN(n589) );
  DFF_X1 \DP/RegALU1/DOUT_reg[28]  ( .D(\DP/RegALU1/N31 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[28] ), .QN(n1391) );
  DFF_X1 \DP/RegALU1/DOUT_reg[0]  ( .D(\DP/RegALU1/N3 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[0]), .QN(n1393) );
  DFF_X1 \DP/RegALU1/DOUT_reg[11]  ( .D(\DP/RegALU1/N14 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[11]), .QN(n1423) );
  DFF_X1 \DP/RegALU1/DOUT_reg[9]  ( .D(\DP/RegALU1/N12 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[9]), .QN(n1439) );
  DFF_X1 \DP/RegALU1/DOUT_reg[7]  ( .D(\DP/RegALU1/N10 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[7]), .QN(n1441) );
  DFF_X1 \DP/RegALU1/DOUT_reg[20]  ( .D(\DP/RegALU1/N23 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[20] ), .QN(n1430) );
  DFF_X1 \DP/RegALU1/DOUT_reg[21]  ( .D(\DP/RegALU1/N24 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[21] ), .QN(n1429) );
  DFF_X1 \DP/RegALU1/DOUT_reg[15]  ( .D(\DP/RegALU1/N18 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[15] ), .QN(n1379) );
  DFF_X1 \DP/RegALU1/DOUT_reg[13]  ( .D(\DP/RegALU1/N16 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[13] ), .QN(n1421) );
  DFF_X1 \DP/RegALU1/DOUT_reg[14]  ( .D(\DP/RegALU1/N17 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[14] ), .QN(n1420) );
  DFF_X1 \DP/RegALU1/DOUT_reg[12]  ( .D(\DP/RegALU1/N15 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[12] ), .QN(n1422) );
  DFF_X1 \DP/RegALU1/DOUT_reg[17]  ( .D(\DP/RegALU1/N20 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[17] ), .QN(n1377) );
  DFF_X1 \DP/RegALU1/DOUT_reg[25]  ( .D(\DP/RegALU1/N28 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[25] ), .QN(n1387) );
  DFF_X1 \DP/RegALU1/DOUT_reg[16]  ( .D(\DP/RegALU1/N19 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[16] ), .QN(n1378) );
  DFF_X1 \DP/RegALU1/DOUT_reg[10]  ( .D(\DP/RegALU1/N13 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[10]), .QN(n1438) );
  DFF_X1 \DP/RegALU1/DOUT_reg[18]  ( .D(\DP/RegALU1/N21 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[18] ), .QN(n1376) );
  DFF_X1 \DP/RegALU1/DOUT_reg[23]  ( .D(\DP/RegALU1/N26 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[23] ), .QN(n1389) );
  DFF_X1 \DP/RegALU1/DOUT_reg[22]  ( .D(\DP/RegALU1/N25 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[22] ), .QN(n1428) );
  DFF_X1 \DP/RegNPC/DOUT_reg[26]  ( .D(\PC/N29 ), .CK(n635), .Q(\DP/NPC1[26] ), 
        .QN(n1291) );
  DFF_X1 \DP/RegALU1/DOUT_reg[27]  ( .D(\DP/RegALU1/N30 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[27] ), .QN(n1392) );
  DFF_X1 \DP/RegALU1/DOUT_reg[8]  ( .D(\DP/RegALU1/N11 ), .CK(
        \DP/RegALU1/net7068 ), .Q(DRAM_ADDR[8]), .QN(n1440) );
  DFF_X1 \DP/RegALU1/DOUT_reg[29]  ( .D(\DP/RegALU1/N32 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[29] ), .QN(n1390) );
  DFF_X1 \DP/RegALU1/DOUT_reg[24]  ( .D(\DP/RegALU1/N27 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[24] ), .QN(n1388) );
  DFF_X1 \DP/RegALU1/DOUT_reg[19]  ( .D(\DP/RegALU1/N22 ), .CK(
        \DP/RegALU1/net7068 ), .Q(\DP/RegALU1_out[19] ), .QN(n1431) );
  DFF_X1 \CU/cw1_reg[22]  ( .D(\CU/N62 ), .CK(CLK), .Q(w_MuxA_SEL), .QN(n608)
         );
  DFF_X1 \DP/FFDBRANCH/Q_reg  ( .D(\DP/FFDBRANCH/N3 ), .CK(
        \DP/FFDBRANCH/net7032 ), .Q(\DP/OUTCOME ), .QN(n607) );
  DFF_X1 \DP/RegFC/DOUT_reg[2]  ( .D(\DP/RegFC/N5 ), .CK(\DP/RegNPC1/net7068 ), 
        .Q(\DP/FwdA[2] ), .QN(n77) );
  DFF_X1 \DP/RegFB/DOUT_reg[1]  ( .D(\DP/RegFB/N4 ), .CK(\DP/RegNPC1/net7068 ), 
        .Q(\DP/FwdB[1] ), .QN(n604) );
  DFF_X1 \DP/RegFC/DOUT_reg[1]  ( .D(\DP/RegFC/N4 ), .CK(\DP/RegNPC1/net7068 ), 
        .Q(\DP/FwdC[1] ), .QN(n69) );
  DFF_X1 \DP/RegFC/DOUT_reg[0]  ( .D(\DP/RegFC/N3 ), .CK(\DP/RegNPC1/net7068 ), 
        .Q(n588), .QN(n76) );
  DFF_X1 \DP/RegFB/DOUT_reg[0]  ( .D(\DP/RegFB/N3 ), .CK(\DP/RegNPC1/net7068 ), 
        .Q(\DP/FwdB[0] ), .QN(n605) );
  DFF_X2 \DP/FFDJL2/Q_reg  ( .D(\DP/FFDJL2/N3 ), .CK(\DP/FFDJL2/net7032 ), .Q(
        \DP/JL2 ), .QN(n1487) );
  CLKBUF_X1 U2578 ( .A(\DP/JL2 ), .Z(n1492) );
  ALU_WIDTH32_RADIX4_OPCODE6 \DP/ALU0  ( .A({\DP/A[31] , \DP/A[30] , 
        \DP/A[29] , \DP/A[28] , \DP/A[27] , \DP/A[26] , \DP/A[25] , \DP/A[24] , 
        \DP/A[23] , \DP/A[22] , \DP/A[21] , \DP/A[20] , \DP/A[19] , \DP/A[18] , 
        \DP/A[17] , \DP/A[16] , \DP/A[15] , \DP/A[14] , \DP/A[13] , \DP/A[12] , 
        \DP/A[11] , \DP/A[10] , \DP/A[9] , \DP/A[8] , \DP/A[7] , \DP/A[6] , 
        \DP/A[5] , \DP/A[4] , \DP/A[3] , \DP/A[2] , \DP/A[1] , \DP/A[0] }), 
        .B({\DP/B[31] , \DP/B[30] , \DP/B[29] , \DP/B[28] , \DP/B[27] , 
        \DP/B[26] , \DP/B[25] , \DP/B[24] , \DP/B[23] , \DP/B[22] , \DP/B[21] , 
        \DP/B[20] , \DP/B[19] , \DP/B[18] , \DP/B[17] , \DP/B[16] , \DP/B[15] , 
        \DP/B[14] , \DP/B[13] , \DP/B[12] , \DP/B[11] , \DP/B[10] , \DP/B[9] , 
        \DP/B[8] , \DP/B[7] , \DP/B[6] , \DP/B[5] , \DP/B[4] , \DP/B[3] , 
        \DP/B[2] , \DP/B[1] , \DP/B[0] }), .OP(w_ALU_OPCODE), .Y({\DP/RES[31] , 
        \DP/RES[30] , \DP/RES[29] , \DP/RES[28] , \DP/RES[27] , \DP/RES[26] , 
        \DP/RES[25] , \DP/RES[24] , \DP/RES[23] , \DP/RES[22] , \DP/RES[21] , 
        \DP/RES[20] , \DP/RES[19] , \DP/RES[18] , \DP/RES[17] , \DP/RES[16] , 
        \DP/RES[15] , \DP/RES[14] , \DP/RES[13] , \DP/RES[12] , \DP/RES[11] , 
        \DP/RES[10] , \DP/RES[9] , \DP/RES[8] , \DP/RES[7] , \DP/RES[6] , 
        \DP/RES[5] , \DP/RES[4] , \DP/RES[3] , \DP/RES[2] , \DP/RES[1] , 
        \DP/RES[0] }) );
  REGISTER_FILE_WIDTH32_LENGTH5 \DP/RF0  ( .CLK(CLK), .RST(RST), .EN(
        \DP/RF_EN ), .RD1(w_RF_RD1), .RD2(n1574), .WR(w_RF_WE), .DATAIN({
        \DP/RF_DATA[31] , \DP/RF_DATA[30] , \DP/RF_DATA[29] , \DP/RF_DATA[28] , 
        \DP/RF_DATA[27] , \DP/RF_DATA[26] , \DP/RF_DATA[25] , \DP/RF_DATA[24] , 
        \DP/RF_DATA[23] , \DP/RF_DATA[22] , \DP/RF_DATA[21] , \DP/RF_DATA[20] , 
        \DP/RF_DATA[19] , \DP/RF_DATA[18] , \DP/RF_DATA[17] , \DP/RF_DATA[16] , 
        \DP/RF_DATA[15] , \DP/RF_DATA[14] , \DP/RF_DATA[13] , \DP/RF_DATA[12] , 
        \DP/RF_DATA[11] , \DP/RF_DATA[10] , \DP/RF_DATA[9] , \DP/RF_DATA[8] , 
        \DP/RF_DATA[7] , \DP/RF_DATA[6] , \DP/RF_DATA[5] , \DP/RF_DATA[4] , 
        \DP/RF_DATA[3] , \DP/RF_DATA[2] , \DP/RF_DATA[1] , \DP/RF_DATA[0] }), 
        .OUT1({\DP/RegA_in[31] , \DP/RegA_in[30] , \DP/RegA_in[29] , 
        \DP/RegA_in[28] , \DP/RegA_in[27] , \DP/RegA_in[26] , \DP/RegA_in[25] , 
        \DP/RegA_in[24] , \DP/RegA_in[23] , \DP/RegA_in[22] , \DP/RegA_in[21] , 
        \DP/RegA_in[20] , \DP/RegA_in[19] , \DP/RegA_in[18] , \DP/RegA_in[17] , 
        \DP/RegA_in[16] , \DP/RegA_in[15] , \DP/RegA_in[14] , \DP/RegA_in[13] , 
        \DP/RegA_in[12] , \DP/RegA_in[11] , \DP/RegA_in[10] , \DP/RegA_in[9] , 
        \DP/RegA_in[8] , \DP/RegA_in[7] , \DP/RegA_in[6] , \DP/RegA_in[5] , 
        \DP/RegA_in[4] , \DP/RegA_in[3] , \DP/RegA_in[2] , \DP/RegA_in[1] , 
        \DP/RegA_in[0] }), .OUT2({\DP/RegB_in[31] , \DP/RegB_in[30] , 
        \DP/RegB_in[29] , \DP/RegB_in[28] , \DP/RegB_in[27] , \DP/RegB_in[26] , 
        \DP/RegB_in[25] , \DP/RegB_in[24] , \DP/RegB_in[23] , \DP/RegB_in[22] , 
        \DP/RegB_in[21] , \DP/RegB_in[20] , \DP/RegB_in[19] , \DP/RegB_in[18] , 
        \DP/RegB_in[17] , \DP/RegB_in[16] , \DP/RegB_in[15] , \DP/RegB_in[14] , 
        \DP/RegB_in[13] , \DP/RegB_in[12] , \DP/RegB_in[11] , \DP/RegB_in[10] , 
        \DP/RegB_in[9] , \DP/RegB_in[8] , \DP/RegB_in[7] , \DP/RegB_in[6] , 
        \DP/RegB_in[5] , \DP/RegB_in[4] , \DP/RegB_in[3] , \DP/RegB_in[2] , 
        \DP/RegB_in[1] , \DP/RegB_in[0] }), .ADD_WR({\DP/RF_ADDR[4] , 
        \DP/RF_ADDR[3] , \DP/RF_ADDR[2] , \DP/RF_ADDR[1] , \DP/RF_ADDR[0] }), 
        .ADD_RD1({n42, n41, n40, n39, n38}), .ADD_RD2({n35, n37, n1295, n34, 
        n36}) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH5_0 \DP/RegRD1/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegRD1/N2 ), .ENCLK(\DP/RegRD1/net7086 ), .TE(1'b0)
         );
  SNPS_CLOCK_GATE_HIGH_FFD_0 \DP/FFDBRANCH/clk_gate_Q_reg  ( .CLK(CLK), .EN(
        \DP/FFDBRANCH/N2 ), .ENCLK(\DP/FFDBRANCH/net7032 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_12 \DP/RegNPC/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\PC/N2 ), .ENCLK(\DP/RegNPC/net7068 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_11 \DP/RegNPC1/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegNPC1/N2 ), .ENCLK(\DP/RegNPC1/net7068 ), .TE(
        1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_10 \DP/RegA/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegA/N2 ), .ENCLK(\DP/RegA/net7068 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_9 \DP/RegB/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegB/N2 ), .ENCLK(\DP/RegB/net7068 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_8 \DP/RegIMM/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegIMM/N2 ), .ENCLK(\DP/RegIMM/net7068 ), .TE(1'b0)
         );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_7 \DP/RegA1/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegA1/N2 ), .ENCLK(\DP/RegA1/net7068 ), .TE(1'b0)
         );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_6 \DP/RegNPC2/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegNPC2/N2 ), .ENCLK(\DP/RegNPC2/net7068 ), .TE(
        1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_5 \DP/RegALU1/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegALU1/N2 ), .ENCLK(\DP/RegALU1/net7068 ), .TE(
        1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_4 \DP/RegME/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegME/N2 ), .ENCLK(\DP/RegME/net7068 ), .TE(1'b0)
         );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH5_2 \DP/RegRD2/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegRD2/N2 ), .ENCLK(\DP/RegRD2/net7086 ), .TE(1'b0)
         );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_3 \DP/RegALU2/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegALU2/N2 ), .ENCLK(\DP/RegALU2/net7068 ), .TE(
        1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_2 \DP/RegLMD/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegLMD/N2 ), .ENCLK(\DP/RegLMD/net7068 ), .TE(1'b0)
         );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH5_1 \DP/RegRD3/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegRD3/N2 ), .ENCLK(\DP/RegRD3/net7086 ), .TE(1'b0)
         );
  SNPS_CLOCK_GATE_HIGH_FFD_2 \DP/FFDJL2/clk_gate_Q_reg  ( .CLK(CLK), .EN(
        \DP/FFDJL2/N2 ), .ENCLK(\DP/FFDJL2/net7032 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_1 \DP/RegNPC3/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegNPC3/N2 ), .ENCLK(\DP/RegNPC3/net7068 ), .TE(
        1'b0) );
  OR2_X2 U1316 ( .A1(\DP/JL2 ), .A2(\DP/RD3[4] ), .ZN(\DP/RF_ADDR[4] ) );
  NAND2_X2 U1324 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[4] ), .ZN(n967) );
  OR2_X2 U1333 ( .A1(\DP/JL2 ), .A2(\DP/RD3[0] ), .ZN(\DP/RF_ADDR[0] ) );
  NAND2_X2 U1335 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[30] ), .ZN(n964) );
  NAND2_X2 U1339 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[5] ), .ZN(n968) );
  NAND2_X2 U1815 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[20] ), .ZN(n953) );
  OR2_X2 U1827 ( .A1(n1255), .A2(\DP/JL2 ), .ZN(n1522) );
  OAI21_X2 U1828 ( .B1(n1227), .B2(\DP/JL2 ), .A(n948), .ZN(\DP/RF_DATA[16] )
         );
  NAND2_X2 U1834 ( .A1(n1856), .A2(n1855), .ZN(\DP/RF_DATA[0] ) );
  NAND2_X2 U1849 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[0] ), .ZN(n1855) );
  NAND2_X2 U1854 ( .A1(n942), .A2(n1861), .ZN(n1856) );
  OAI21_X2 U1856 ( .B1(n1229), .B2(\DP/JL2 ), .A(n1857), .ZN(\DP/RF_DATA[17] )
         );
  NAND2_X2 U2265 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[17] ), .ZN(n1857) );
  NAND2_X2 U2580 ( .A1(n971), .A2(n1858), .ZN(\DP/RF_DATA[9] ) );
  NAND2_X2 U2581 ( .A1(n1859), .A2(n1861), .ZN(n1858) );
  INV_X2 U2603 ( .A(n1270), .ZN(n1859) );
  NAND2_X2 U2607 ( .A1(n960), .A2(n1860), .ZN(\DP/RF_DATA[27] ) );
  NAND2_X2 U2627 ( .A1(n1862), .A2(n1861), .ZN(n1860) );
  INV_X2 U2661 ( .A(\DP/JL2 ), .ZN(n1861) );
  INV_X2 U2662 ( .A(n1249), .ZN(n1862) );
endmodule


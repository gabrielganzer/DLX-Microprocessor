
module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_0 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_1 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_2 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_3 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_4 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_5 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_6 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_7 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_8 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_9 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_10 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_11 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_12 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_13 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_14 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_15 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_16 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_17 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_18 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_19 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_20 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_21 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_22 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_23 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_24 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_25 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_26 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_27 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_28 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_29 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_30 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_31 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_32 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_33 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net234775, n2, n3;
  assign net234775 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net234775), .A2(TE), .ZN(n3) );
endmodule


module REGISTER_FILE_WIDTH32_LENGTH5 ( CLK, RST, EN, RD1, RD2, WR, DATAIN, 
        OUT1, OUT2, ADD_WR, ADD_RD1, ADD_RD2 );
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input CLK, RST, EN, RD1, RD2, WR;
  wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n20327, n5910, n5911, n5912, n5913, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n32665, n32666, n32667, n32668, n32669, n32670,
         n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678,
         n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686,
         n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694,
         n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702,
         n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710,
         n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718,
         n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726,
         n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734,
         n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742,
         n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750,
         n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758,
         n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766,
         n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774,
         n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782,
         n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790,
         n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798,
         n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806,
         n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814,
         n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822,
         n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830,
         n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838,
         n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846,
         n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854,
         n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862,
         n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870,
         n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878,
         n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886,
         n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894,
         n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902,
         n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910,
         n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918,
         n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926,
         n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934,
         n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942,
         n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950,
         n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958,
         n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966,
         n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974,
         n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982,
         n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990,
         n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998,
         n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006,
         n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014,
         n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022,
         n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030,
         n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038,
         n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046,
         n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054,
         n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062,
         n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070,
         n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078,
         n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086,
         n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094,
         n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102,
         n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110,
         n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118,
         n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126,
         n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134,
         n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142,
         n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150,
         n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158,
         n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166,
         n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174,
         n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182,
         n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190,
         n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198,
         n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206,
         n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214,
         n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222,
         n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230,
         n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238,
         n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246,
         n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254,
         n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262,
         n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270,
         n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278,
         n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286,
         n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294,
         n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302,
         n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310,
         n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318,
         n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326,
         n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334,
         n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342,
         n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350,
         n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358,
         n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366,
         n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374,
         n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382,
         n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390,
         n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398,
         n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406,
         n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414,
         n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422,
         n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430,
         n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438,
         n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446,
         n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454,
         n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462,
         n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470,
         n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478,
         n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486,
         n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494,
         n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502,
         n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510,
         n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518,
         n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526,
         n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534,
         n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542,
         n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550,
         n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558,
         n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566,
         n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574,
         n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582,
         n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590,
         n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598,
         n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606,
         n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614,
         n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622,
         n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630,
         n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638,
         n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646,
         n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654,
         n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662,
         n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670,
         n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678,
         n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
         n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694,
         n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702,
         n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710,
         n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718,
         n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726,
         n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734,
         n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
         n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750,
         n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758,
         n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766,
         n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774,
         n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782,
         n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790,
         n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798,
         n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806,
         n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814,
         n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822,
         n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830,
         n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838,
         n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846,
         n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
         n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862,
         n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870,
         n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878,
         n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886,
         n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894,
         n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902,
         n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910,
         n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918,
         n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926,
         n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934,
         n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942,
         n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950,
         n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958,
         n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966,
         n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974,
         n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982,
         n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990,
         n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998,
         n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006,
         n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014,
         n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022,
         n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030,
         n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038,
         n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046,
         n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054,
         n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062,
         n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
         n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078,
         n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086,
         n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094,
         n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102,
         n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110,
         n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118,
         n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126,
         n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134,
         n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142,
         n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150,
         n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158,
         n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166,
         n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174,
         n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182,
         n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190,
         n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198,
         n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206,
         n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214,
         n34215, n34216;

  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n5912), .CK(n5878), .Q(n7464) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n5911), .CK(n5878), .Q(n7496) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n5910), .CK(n5878), .Q(n7528) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n32683), .CK(n5878), .Q(n7560) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n5912), .CK(n5889), .Q(n7452) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n5911), .CK(n5889), .Q(n7484) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n5910), .CK(n5889), .Q(n7516) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n5912), .CK(n5900), .Q(n7450) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n5911), .CK(n5900), .Q(n7482) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n5910), .CK(n5900), .Q(n7514) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n5912), .CK(n5903), .Q(n7455) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n5911), .CK(n5903), .Q(n7487) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n5910), .CK(n5903), .Q(n7519) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n5912), .CK(n5904), .Q(n7457) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n5911), .CK(n5904), .Q(n7489) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n5910), .CK(n5904), .Q(n7521) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n5912), .CK(n5905), .Q(n7462) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n5911), .CK(n5905), .Q(n7494) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n5910), .CK(n5905), .Q(n7526) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n5912), .CK(n5906), .Q(n7436) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n5911), .CK(n5906), .Q(n7468) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n5910), .CK(n5906), .Q(n7500) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n5912), .CK(n5907), .Q(n7460) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n5911), .CK(n5907), .Q(n7492) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n5910), .CK(n5907), .Q(n7524) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n5912), .CK(n5908), .Q(n7456) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n5911), .CK(n5908), .Q(n7488) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n5910), .CK(n5908), .Q(n7520) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n5912), .CK(n5909), .Q(n7449) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n5911), .CK(n5909), .Q(n7481) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n5910), .CK(n5909), .Q(n7513) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n5912), .CK(n5879), .Q(n7451) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n5911), .CK(n5879), .Q(n7483) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n5910), .CK(n5879), .Q(n7515) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n5912), .CK(n5880), .Q(n7439) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n5911), .CK(n5880), .Q(n7471) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n5910), .CK(n5880), .Q(n7503) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n5912), .CK(n5881), .Q(n7441) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n5911), .CK(n5881), .Q(n7473) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n5910), .CK(n5881), .Q(n7505) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n5912), .CK(n5882), .Q(n7463) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n5911), .CK(n5882), .Q(n7495) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n5910), .CK(n5882), .Q(n7527) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n5912), .CK(n5883), .Q(n7438) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n5911), .CK(n5883), .Q(n7470) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n5910), .CK(n5883), .Q(n7502) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n5912), .CK(n5884), .Q(n7437) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n5911), .CK(n5884), .Q(n7469) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n5910), .CK(n5884), .Q(n7501) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n5912), .CK(n5885), .Q(n7453) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n5911), .CK(n5885), .Q(n7485) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n5910), .CK(n5885), .Q(n7517) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n5912), .CK(n5886), .Q(n7442) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n5911), .CK(n5886), .Q(n7474) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n5910), .CK(n5886), .Q(n7506) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n5912), .CK(n5887), .Q(n7461) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n5911), .CK(n5887), .Q(n7493) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n5910), .CK(n5887), .Q(n7525) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n5912), .CK(n5888), .Q(n7440) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n5911), .CK(n5888), .Q(n7472) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n5910), .CK(n5888), .Q(n7504) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n5912), .CK(n5890), .Q(n7433) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n5911), .CK(n5890), .Q(n7465) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n5910), .CK(n5890), .Q(n7497) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n5912), .CK(n5891), .Q(n7435) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n5911), .CK(n5891), .Q(n7467) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n5910), .CK(n5891), .Q(n7499) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n5912), .CK(n5892), .Q(n7454) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n5911), .CK(n5892), .Q(n7486) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n5910), .CK(n5892), .Q(n7518) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n5912), .CK(n5893), .Q(n7448) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n5911), .CK(n5893), .Q(n7480) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n5910), .CK(n5893), .Q(n7512) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n5912), .CK(n5894), .Q(n7458) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n5911), .CK(n5894), .Q(n7490) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n5910), .CK(n5894), .Q(n7522) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n5912), .CK(n5895), .Q(n7443) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n5911), .CK(n5895), .Q(n7475) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n5910), .CK(n5895), .Q(n7507) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n5912), .CK(n5896), .Q(n7447) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n5911), .CK(n5896), .Q(n7479) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n5910), .CK(n5896), .Q(n7511) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n5912), .CK(n5897), .Q(n7459) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n5911), .CK(n5897), .Q(n7491) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n5910), .CK(n5897), .Q(n7523) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n5912), .CK(n5898), .Q(n7434) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n5911), .CK(n5898), .Q(n7466) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n5910), .CK(n5898), .Q(n7498) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n5912), .CK(n5899), .Q(n7446) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n5911), .CK(n5899), .Q(n7478) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n5910), .CK(n5899), .Q(n7510) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n5912), .CK(n5901), .Q(n7444) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n5911), .CK(n5901), .Q(n7476) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n5910), .CK(n5901), .Q(n7508) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n5912), .CK(n5902), .Q(n7445) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n5911), .CK(n5902), .Q(n7477) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n5910), .CK(n5902), .Q(n7509) );
  DFF_X1 \OUT1_reg[31]  ( .D(n5777), .CK(n5809), .Q(OUT1[31]) );
  DFF_X1 \OUT1_reg[29]  ( .D(n5779), .CK(n5809), .Q(OUT1[29]) );
  DFF_X1 \OUT1_reg[28]  ( .D(n5780), .CK(n5809), .Q(OUT1[28]) );
  DFF_X1 \OUT1_reg[27]  ( .D(n5781), .CK(n5809), .Q(OUT1[27]) );
  DFF_X1 \OUT1_reg[26]  ( .D(n5782), .CK(n5809), .Q(OUT1[26]) );
  DFF_X1 \OUT1_reg[25]  ( .D(n5783), .CK(n5809), .Q(OUT1[25]) );
  DFF_X1 \OUT1_reg[24]  ( .D(n5784), .CK(n5809), .Q(OUT1[24]) );
  DFF_X1 \OUT1_reg[23]  ( .D(n5785), .CK(n5809), .Q(OUT1[23]) );
  DFF_X1 \OUT1_reg[22]  ( .D(n5786), .CK(n5809), .Q(OUT1[22]) );
  DFF_X1 \OUT1_reg[21]  ( .D(n5787), .CK(n5809), .Q(OUT1[21]) );
  DFF_X1 \OUT1_reg[20]  ( .D(n5788), .CK(n5809), .Q(OUT1[20]) );
  DFF_X1 \OUT1_reg[19]  ( .D(n5789), .CK(n5809), .Q(OUT1[19]) );
  DFF_X1 \OUT1_reg[18]  ( .D(n5790), .CK(n5809), .Q(OUT1[18]) );
  DFF_X1 \OUT1_reg[17]  ( .D(n5791), .CK(n5809), .Q(OUT1[17]) );
  DFF_X1 \OUT1_reg[16]  ( .D(n5792), .CK(n5809), .Q(OUT1[16]) );
  DFF_X1 \OUT1_reg[15]  ( .D(n5793), .CK(n5809), .Q(OUT1[15]) );
  DFF_X1 \OUT1_reg[14]  ( .D(n5794), .CK(n5809), .Q(OUT1[14]) );
  DFF_X1 \OUT1_reg[13]  ( .D(n5795), .CK(n5809), .Q(OUT1[13]) );
  DFF_X1 \OUT1_reg[12]  ( .D(n5796), .CK(n5809), .Q(OUT1[12]) );
  DFF_X1 \OUT1_reg[11]  ( .D(n5797), .CK(n5809), .Q(OUT1[11]) );
  DFF_X1 \OUT1_reg[10]  ( .D(n5798), .CK(n5809), .Q(OUT1[10]) );
  DFF_X1 \OUT1_reg[9]  ( .D(n5799), .CK(n5809), .Q(OUT1[9]) );
  DFF_X1 \OUT1_reg[8]  ( .D(n5800), .CK(n5809), .Q(OUT1[8]) );
  DFF_X1 \OUT1_reg[7]  ( .D(n5801), .CK(n5809), .Q(OUT1[7]) );
  DFF_X1 \OUT1_reg[6]  ( .D(n5802), .CK(n5809), .Q(OUT1[6]) );
  DFF_X1 \OUT1_reg[5]  ( .D(n5803), .CK(n5809), .Q(OUT1[5]) );
  DFF_X1 \OUT1_reg[4]  ( .D(n5804), .CK(n5809), .Q(OUT1[4]) );
  DFF_X1 \OUT1_reg[3]  ( .D(n5805), .CK(n5809), .Q(OUT1[3]) );
  DFF_X1 \OUT1_reg[2]  ( .D(n5806), .CK(n5809), .Q(OUT1[2]) );
  DFF_X1 \OUT1_reg[1]  ( .D(n5807), .CK(n5809), .Q(OUT1[1]) );
  DFF_X1 \OUT1_reg[0]  ( .D(n5808), .CK(n5809), .Q(OUT1[0]) );
  DFF_X1 \OUT2_reg[31]  ( .D(n5812), .CK(n5844), .Q(OUT2[31]) );
  DFF_X1 \OUT2_reg[30]  ( .D(n5813), .CK(n5844), .Q(OUT2[30]) );
  DFF_X1 \OUT2_reg[29]  ( .D(n5814), .CK(n5844), .Q(OUT2[29]) );
  DFF_X1 \OUT2_reg[28]  ( .D(n5815), .CK(n5844), .Q(OUT2[28]) );
  DFF_X1 \OUT2_reg[27]  ( .D(n5816), .CK(n5844), .Q(OUT2[27]) );
  DFF_X1 \OUT2_reg[26]  ( .D(n5817), .CK(n5844), .Q(OUT2[26]) );
  DFF_X1 \OUT2_reg[25]  ( .D(n5818), .CK(n5844), .Q(OUT2[25]) );
  DFF_X1 \OUT2_reg[24]  ( .D(n5819), .CK(n5844), .Q(OUT2[24]) );
  DFF_X1 \OUT2_reg[23]  ( .D(n5820), .CK(n5844), .Q(OUT2[23]) );
  DFF_X1 \OUT2_reg[22]  ( .D(n5821), .CK(n5844), .Q(OUT2[22]) );
  DFF_X1 \OUT2_reg[21]  ( .D(n5822), .CK(n5844), .Q(OUT2[21]) );
  DFF_X1 \OUT2_reg[20]  ( .D(n5823), .CK(n5844), .Q(OUT2[20]) );
  DFF_X1 \OUT2_reg[19]  ( .D(n5824), .CK(n5844), .Q(OUT2[19]) );
  DFF_X1 \OUT2_reg[18]  ( .D(n5825), .CK(n5844), .Q(OUT2[18]) );
  DFF_X1 \OUT2_reg[17]  ( .D(n5826), .CK(n5844), .Q(OUT2[17]) );
  DFF_X1 \OUT2_reg[16]  ( .D(n5827), .CK(n5844), .Q(OUT2[16]) );
  DFF_X1 \OUT2_reg[15]  ( .D(n5828), .CK(n5844), .Q(OUT2[15]) );
  DFF_X1 \OUT2_reg[14]  ( .D(n5829), .CK(n5844), .Q(OUT2[14]) );
  DFF_X1 \OUT2_reg[13]  ( .D(n5830), .CK(n5844), .Q(OUT2[13]) );
  DFF_X1 \OUT2_reg[12]  ( .D(n5831), .CK(n5844), .Q(OUT2[12]) );
  DFF_X1 \OUT2_reg[11]  ( .D(n5832), .CK(n5844), .Q(OUT2[11]) );
  DFF_X1 \OUT2_reg[10]  ( .D(n5833), .CK(n5844), .Q(OUT2[10]) );
  DFF_X1 \OUT2_reg[9]  ( .D(n5834), .CK(n5844), .Q(OUT2[9]) );
  DFF_X1 \OUT2_reg[8]  ( .D(n5835), .CK(n5844), .Q(OUT2[8]) );
  DFF_X1 \OUT2_reg[7]  ( .D(n5836), .CK(n5844), .Q(OUT2[7]) );
  DFF_X1 \OUT2_reg[6]  ( .D(n5837), .CK(n5844), .Q(OUT2[6]) );
  DFF_X1 \OUT2_reg[5]  ( .D(n5838), .CK(n5844), .Q(OUT2[5]) );
  DFF_X1 \OUT2_reg[4]  ( .D(n5839), .CK(n5844), .Q(OUT2[4]) );
  DFF_X1 \OUT2_reg[3]  ( .D(n5840), .CK(n5844), .Q(OUT2[3]) );
  DFF_X1 \OUT2_reg[2]  ( .D(n5841), .CK(n5844), .Q(OUT2[2]) );
  DFF_X1 \OUT2_reg[1]  ( .D(n5842), .CK(n5844), .Q(OUT2[1]) );
  DFF_X1 \OUT2_reg[0]  ( .D(n5843), .CK(n5844), .Q(OUT2[0]) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_0 \clk_gate_REGISTERS_reg[9]  ( 
        .CLK(CLK), .EN(n1063), .ENCLK(n5909), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_1 \clk_gate_REGISTERS_reg[8]  ( 
        .CLK(CLK), .EN(n1064), .ENCLK(n5908), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_2 \clk_gate_REGISTERS_reg[7]  ( 
        .CLK(CLK), .EN(n1072), .ENCLK(n5907), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_3 \clk_gate_REGISTERS_reg[6]  ( 
        .CLK(CLK), .EN(n1071), .ENCLK(n5906), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_4 \clk_gate_REGISTERS_reg[5]  ( 
        .CLK(CLK), .EN(n1065), .ENCLK(n5905), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_5 \clk_gate_REGISTERS_reg[4]  ( 
        .CLK(CLK), .EN(n1066), .ENCLK(n5904), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_6 \clk_gate_REGISTERS_reg[3]  ( 
        .CLK(CLK), .EN(n1070), .ENCLK(n5903), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_7 \clk_gate_REGISTERS_reg[31]  ( 
        .CLK(CLK), .EN(n1045), .ENCLK(n5902), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_8 \clk_gate_REGISTERS_reg[30]  ( 
        .CLK(CLK), .EN(n1046), .ENCLK(n5901), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_9 \clk_gate_REGISTERS_reg[2]  ( 
        .CLK(CLK), .EN(n1069), .ENCLK(n5900), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_10 \clk_gate_REGISTERS_reg[29]  ( 
        .CLK(CLK), .EN(n1076), .ENCLK(n5899), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_11 \clk_gate_REGISTERS_reg[28]  ( 
        .CLK(CLK), .EN(n1075), .ENCLK(n5898), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_12 \clk_gate_REGISTERS_reg[27]  ( 
        .CLK(CLK), .EN(n1047), .ENCLK(n5897), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_13 \clk_gate_REGISTERS_reg[26]  ( 
        .CLK(CLK), .EN(n1048), .ENCLK(n5896), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_14 \clk_gate_REGISTERS_reg[25]  ( 
        .CLK(CLK), .EN(n1074), .ENCLK(n5895), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_15 \clk_gate_REGISTERS_reg[24]  ( 
        .CLK(CLK), .EN(n1073), .ENCLK(n5894), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_16 \clk_gate_REGISTERS_reg[23]  ( 
        .CLK(CLK), .EN(n1049), .ENCLK(n5893), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_17 \clk_gate_REGISTERS_reg[22]  ( 
        .CLK(CLK), .EN(n1050), .ENCLK(n5892), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_18 \clk_gate_REGISTERS_reg[21]  ( 
        .CLK(CLK), .EN(n1051), .ENCLK(n5891), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_19 \clk_gate_REGISTERS_reg[20]  ( 
        .CLK(CLK), .EN(n1052), .ENCLK(n5890), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_20 \clk_gate_REGISTERS_reg[1]  ( 
        .CLK(CLK), .EN(n1067), .ENCLK(n5889), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_21 \clk_gate_REGISTERS_reg[19]  ( 
        .CLK(CLK), .EN(n1053), .ENCLK(n5888), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_22 \clk_gate_REGISTERS_reg[18]  ( 
        .CLK(CLK), .EN(n1054), .ENCLK(n5887), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_23 \clk_gate_REGISTERS_reg[17]  ( 
        .CLK(CLK), .EN(n1055), .ENCLK(n5886), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_24 \clk_gate_REGISTERS_reg[16]  ( 
        .CLK(CLK), .EN(n1056), .ENCLK(n5885), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_25 \clk_gate_REGISTERS_reg[15]  ( 
        .CLK(CLK), .EN(n1057), .ENCLK(n5884), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_26 \clk_gate_REGISTERS_reg[14]  ( 
        .CLK(CLK), .EN(n1058), .ENCLK(n5883), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_27 \clk_gate_REGISTERS_reg[13]  ( 
        .CLK(CLK), .EN(n1059), .ENCLK(n5882), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_28 \clk_gate_REGISTERS_reg[12]  ( 
        .CLK(CLK), .EN(n1060), .ENCLK(n5881), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_29 \clk_gate_REGISTERS_reg[11]  ( 
        .CLK(CLK), .EN(n1061), .ENCLK(n5880), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_30 \clk_gate_REGISTERS_reg[10]  ( 
        .CLK(CLK), .EN(n1062), .ENCLK(n5879), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_31 \clk_gate_REGISTERS_reg[0]  ( 
        .CLK(CLK), .EN(n1068), .ENCLK(n5878), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_32 clk_gate_OUT2_reg ( 
        .CLK(CLK), .EN(n5845), .ENCLK(n5844), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_33 clk_gate_OUT1_reg ( 
        .CLK(CLK), .EN(n5811), .ENCLK(n5809), .TE(1'b0) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n14143), .CK(n5902), .QN(n8021) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n14143), .CK(n5901), .QN(n8020) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n14143), .CK(n5899), .QN(n8022) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n14143), .CK(n5898), .QN(n8010) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n14143), .CK(n5897), .QN(n8035) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n14143), .CK(n5896), .QN(n8023) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n14143), .CK(n5895), .QN(n8019) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n14143), .CK(n5894), .QN(n8034) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n14143), .CK(n5893), .QN(n8024) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n14143), .CK(n5892), .QN(n8030) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n14143), .CK(n5891), .QN(n8011) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n14143), .CK(n5890), .QN(n8009) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n14143), .CK(n5888), .QN(n8016) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n14143), .CK(n5887), .QN(n8037) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n14143), .CK(n5886), .QN(n8018) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n14143), .CK(n5885), .QN(n8029) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n14143), .CK(n5884), .QN(n8013) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n14143), .CK(n5883), .QN(n8014) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n14143), .CK(n5882), .QN(n8039) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n14143), .CK(n5881), .QN(n8017) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n14143), .CK(n5880), .QN(n8015) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n14143), .CK(n5879), .QN(n8027) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n14143), .CK(n5909), .QN(n8025) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n14143), .CK(n5908), .QN(n8032) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n14143), .CK(n5907), .QN(n8036) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n14143), .CK(n5906), .QN(n8012) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n14143), .CK(n5905), .QN(n8038) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n14143), .CK(n5904), .QN(n8033) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n14143), .CK(n5903), .QN(n8031) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n14143), .CK(n5900), .QN(n8026) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n14143), .CK(n5889), .QN(n8028) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n14143), .CK(n5878), .QN(n8040) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n14145), .CK(n5902), .QN(n8085) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n14145), .CK(n5901), .QN(n8084) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n14145), .CK(n5899), .QN(n8086) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n14145), .CK(n5898), .QN(n8074) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n14145), .CK(n5897), .QN(n8099) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n14145), .CK(n5896), .QN(n8087) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n14145), .CK(n5895), .QN(n8083) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n14145), .CK(n5894), .QN(n8098) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n14145), .CK(n5893), .QN(n8088) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n14145), .CK(n5892), .QN(n8094) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n14145), .CK(n5891), .QN(n8075) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n14145), .CK(n5890), .QN(n8073) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n14145), .CK(n5888), .QN(n8080) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n14145), .CK(n5887), .QN(n8101) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n14145), .CK(n5886), .QN(n8082) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n14145), .CK(n5885), .QN(n8093) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n14145), .CK(n5884), .QN(n8077) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n14145), .CK(n5883), .QN(n8078) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n14145), .CK(n5882), .QN(n8103) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n14145), .CK(n5881), .QN(n8081) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n14145), .CK(n5880), .QN(n8079) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n14145), .CK(n5879), .QN(n8091) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n14145), .CK(n5909), .QN(n8089) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n14145), .CK(n5908), .QN(n8096) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n14145), .CK(n5907), .QN(n8100) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n14145), .CK(n5906), .QN(n8076) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n14145), .CK(n5905), .QN(n8102) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n14145), .CK(n5904), .QN(n8097) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n14145), .CK(n5903), .QN(n8095) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n14145), .CK(n5900), .QN(n8090) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n14145), .CK(n5889), .QN(n8092) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n14145), .CK(n5878), .QN(n8104) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n14141), .CK(n5902), .QN(n7957) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n32726), .CK(n5902), .QN(n8149) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n14141), .CK(n5901), .QN(n7956) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n32726), .CK(n5901), .QN(n8148) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n14141), .CK(n5899), .QN(n7958) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n32726), .CK(n5899), .QN(n8150) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n14141), .CK(n5898), .QN(n7946) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n14147), .CK(n5898), .QN(n8138) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n14141), .CK(n5897), .QN(n7971) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n14147), .CK(n5897), .QN(n8163) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n14141), .CK(n5896), .QN(n7959) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n14147), .CK(n5896), .QN(n8151) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n14141), .CK(n5895), .QN(n7955) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n14147), .CK(n5895), .QN(n8147) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n14141), .CK(n5894), .QN(n7970) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n14147), .CK(n5894), .QN(n8162) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n14141), .CK(n5893), .QN(n7960) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n14147), .CK(n5893), .QN(n8152) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n14141), .CK(n5892), .QN(n7966) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n14147), .CK(n5892), .QN(n8158) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n14141), .CK(n5891), .QN(n7947) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n14147), .CK(n5891), .QN(n8139) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n14141), .CK(n5890), .QN(n7945) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n14147), .CK(n5890), .QN(n8137) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n14141), .CK(n5888), .QN(n7952) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n14147), .CK(n5888), .QN(n8144) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n14141), .CK(n5887), .QN(n7973) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n14147), .CK(n5887), .QN(n8165) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n14141), .CK(n5886), .QN(n7954) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n14147), .CK(n5886), .QN(n8146) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n14141), .CK(n5885), .QN(n7965) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n14147), .CK(n5885), .QN(n8157) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n14141), .CK(n5884), .QN(n7949) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n14147), .CK(n5884), .QN(n8141) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n14141), .CK(n5883), .QN(n7950) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n14147), .CK(n5883), .QN(n8142) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n14141), .CK(n5882), .QN(n7975) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n14147), .CK(n5882), .QN(n8167) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n14141), .CK(n5881), .QN(n7953) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n14147), .CK(n5881), .QN(n8145) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n14141), .CK(n5880), .QN(n7951) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n32726), .CK(n5880), .QN(n8143) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n14141), .CK(n5879), .QN(n7963) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n32726), .CK(n5879), .QN(n8155) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n14141), .CK(n5909), .QN(n7961) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n32726), .CK(n5909), .QN(n8153) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n14141), .CK(n5908), .QN(n7968) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n32726), .CK(n5908), .QN(n8160) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n14141), .CK(n5907), .QN(n7972) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n32726), .CK(n5907), .QN(n8164) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n14141), .CK(n5906), .QN(n7948) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n32726), .CK(n5906), .QN(n8140) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n14141), .CK(n5905), .QN(n7974) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n32726), .CK(n5905), .QN(n8166) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n14141), .CK(n5904), .QN(n7969) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n32726), .CK(n5904), .QN(n8161) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n14141), .CK(n5903), .QN(n7967) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n32726), .CK(n5903), .QN(n8159) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n14141), .CK(n5900), .QN(n7962) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n32726), .CK(n5900), .QN(n8154) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n14141), .CK(n5889), .QN(n7964) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n32726), .CK(n5889), .QN(n8156) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n14141), .CK(n5878), .QN(n7976) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n14147), .CK(n5878), .QN(n8168) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n14142), .CK(n5902), .QN(n7989) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n14144), .CK(n5902), .QN(n8053) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n14142), .CK(n5901), .QN(n7988) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n14144), .CK(n5901), .QN(n8052) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n14142), .CK(n5899), .QN(n7990) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n14144), .CK(n5899), .QN(n8054) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n14142), .CK(n5898), .QN(n7978) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n14144), .CK(n5898), .QN(n8042) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n14142), .CK(n5897), .QN(n8003) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n14144), .CK(n5897), .QN(n8067) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n14142), .CK(n5896), .QN(n7991) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n14144), .CK(n5896), .QN(n8055) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n14142), .CK(n5895), .QN(n7987) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n14144), .CK(n5895), .QN(n8051) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n14142), .CK(n5894), .QN(n8002) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n14144), .CK(n5894), .QN(n8066) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n14142), .CK(n5893), .QN(n7992) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n14144), .CK(n5893), .QN(n8056) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n14142), .CK(n5892), .QN(n7998) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n14144), .CK(n5892), .QN(n8062) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n14142), .CK(n5891), .QN(n7979) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n14144), .CK(n5891), .QN(n8043) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n14142), .CK(n5890), .QN(n7977) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n14144), .CK(n5890), .QN(n8041) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n14142), .CK(n5888), .QN(n7984) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n14144), .CK(n5888), .QN(n8048) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n14142), .CK(n5887), .QN(n8005) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n14144), .CK(n5887), .QN(n8069) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n14142), .CK(n5886), .QN(n7986) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n14144), .CK(n5886), .QN(n8050) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n14142), .CK(n5885), .QN(n7997) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n14144), .CK(n5885), .QN(n8061) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n14142), .CK(n5884), .QN(n7981) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n14144), .CK(n5884), .QN(n8045) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n14142), .CK(n5883), .QN(n7982) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n14144), .CK(n5883), .QN(n8046) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n14142), .CK(n5882), .QN(n8007) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n14144), .CK(n5882), .QN(n8071) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n14142), .CK(n5881), .QN(n7985) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n14144), .CK(n5881), .QN(n8049) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n14142), .CK(n5880), .QN(n7983) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n14144), .CK(n5880), .QN(n8047) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n14142), .CK(n5879), .QN(n7995) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n14144), .CK(n5879), .QN(n8059) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n14142), .CK(n5909), .QN(n7993) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n14144), .CK(n5909), .QN(n8057) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n14142), .CK(n5908), .QN(n8000) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n14144), .CK(n5908), .QN(n8064) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n14142), .CK(n5907), .QN(n8004) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n14144), .CK(n5907), .QN(n8068) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n14142), .CK(n5906), .QN(n7980) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n14144), .CK(n5906), .QN(n8044) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n14142), .CK(n5905), .QN(n8006) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n14144), .CK(n5905), .QN(n8070) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n14142), .CK(n5904), .QN(n8001) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n14144), .CK(n5904), .QN(n8065) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n14142), .CK(n5903), .QN(n7999) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n14144), .CK(n5903), .QN(n8063) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n14142), .CK(n5900), .QN(n7994) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n14144), .CK(n5900), .QN(n8058) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n14142), .CK(n5889), .QN(n7996) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n14144), .CK(n5889), .QN(n8060) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n14142), .CK(n5878), .QN(n8008) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n14144), .CK(n5878), .QN(n8072) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n14140), .CK(n5902), .QN(n7925) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n14140), .CK(n5901), .QN(n7924) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n14140), .CK(n5899), .QN(n7926) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n14140), .CK(n5898), .QN(n7914) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n14140), .CK(n5897), .QN(n7939) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n14140), .CK(n5896), .QN(n7927) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n14140), .CK(n5895), .QN(n7923) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n14140), .CK(n5894), .QN(n7938) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n14140), .CK(n5893), .QN(n7928) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n14140), .CK(n5892), .QN(n7934) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n14140), .CK(n5891), .QN(n7915) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n14140), .CK(n5890), .QN(n7913) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n14140), .CK(n5888), .QN(n7920) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n14140), .CK(n5887), .QN(n7941) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n14140), .CK(n5886), .QN(n7922) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n14140), .CK(n5885), .QN(n7933) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n14140), .CK(n5884), .QN(n7917) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n14140), .CK(n5883), .QN(n7918) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n14140), .CK(n5882), .QN(n7943) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n14140), .CK(n5881), .QN(n7921) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n14140), .CK(n5880), .QN(n7919) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n14140), .CK(n5879), .QN(n7931) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n14140), .CK(n5909), .QN(n7929) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n14140), .CK(n5908), .QN(n7936) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n14140), .CK(n5907), .QN(n7940) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n14140), .CK(n5906), .QN(n7916) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n14140), .CK(n5905), .QN(n7942) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n14140), .CK(n5904), .QN(n7937) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n14140), .CK(n5903), .QN(n7935) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n14140), .CK(n5900), .QN(n7930) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n14140), .CK(n5889), .QN(n7932) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n14140), .CK(n5878), .QN(n7944) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n32727), .CK(n5902), .QN(n8117) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n14146), .CK(n5901), .QN(n8116) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n14146), .CK(n5899), .QN(n8118) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n32727), .CK(n5898), .QN(n8106) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n32727), .CK(n5897), .QN(n8131) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n14146), .CK(n5896), .QN(n8119) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n14146), .CK(n5895), .QN(n8115) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n14146), .CK(n5894), .QN(n8130) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n14146), .CK(n5893), .QN(n8120) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n14146), .CK(n5892), .QN(n8126) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n14146), .CK(n5891), .QN(n8107) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n32727), .CK(n5890), .QN(n8105) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n32727), .CK(n5888), .QN(n8112) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n14146), .CK(n5887), .QN(n8133) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n32727), .CK(n5886), .QN(n8114) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n32727), .CK(n5885), .QN(n8125) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n14146), .CK(n5884), .QN(n8109) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n14146), .CK(n5883), .QN(n8110) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n14146), .CK(n5882), .QN(n8135) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n14146), .CK(n5881), .QN(n8113) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n14146), .CK(n5880), .QN(n8111) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n14146), .CK(n5879), .QN(n8123) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n14146), .CK(n5909), .QN(n8121) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n14146), .CK(n5908), .QN(n8128) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n32727), .CK(n5907), .QN(n8132) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n32727), .CK(n5906), .QN(n8108) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n32727), .CK(n5905), .QN(n8134) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n32727), .CK(n5904), .QN(n8129) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n32727), .CK(n5903), .QN(n8127) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n32727), .CK(n5900), .QN(n8122) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n32727), .CK(n5889), .QN(n8124) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n14146), .CK(n5878), .QN(n8136) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n14148), .CK(n5902), .QN(n8181) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n14148), .CK(n5901), .QN(n8180) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n14148), .CK(n5899), .QN(n8182) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n14148), .CK(n5898), .QN(n8170) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n14148), .CK(n5897), .QN(n8195) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n14148), .CK(n5896), .QN(n8183) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n14148), .CK(n5895), .QN(n8179) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n14148), .CK(n5894), .QN(n8194) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n14148), .CK(n5893), .QN(n8184) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n14148), .CK(n5892), .QN(n8190) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n14148), .CK(n5891), .QN(n8171) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n14148), .CK(n5890), .QN(n8169) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n14148), .CK(n5888), .QN(n8176) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n14148), .CK(n5887), .QN(n8197) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n14148), .CK(n5886), .QN(n8178) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n14148), .CK(n5885), .QN(n8189) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n14148), .CK(n5884), .QN(n8173) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n14148), .CK(n5883), .QN(n8174) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n14148), .CK(n5882), .QN(n8199) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n14148), .CK(n5881), .QN(n8177) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n14148), .CK(n5880), .QN(n8175) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n14148), .CK(n5879), .QN(n8187) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n14148), .CK(n5909), .QN(n8185) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n14148), .CK(n5908), .QN(n8192) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n14148), .CK(n5907), .QN(n8196) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n14148), .CK(n5906), .QN(n8172) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n14148), .CK(n5905), .QN(n8198) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n14148), .CK(n5904), .QN(n8193) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n14148), .CK(n5903), .QN(n8191) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n14148), .CK(n5900), .QN(n8186) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n14148), .CK(n5889), .QN(n8188) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n14148), .CK(n5878), .QN(n8200) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n32728), .CK(n5902), .QN(n7893) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n32728), .CK(n5901), .QN(n7892) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n32728), .CK(n5899), .QN(n7894) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n14139), .CK(n5898), .QN(n7882) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n14139), .CK(n5897), .QN(n7907) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n14139), .CK(n5896), .QN(n7895) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n14139), .CK(n5895), .QN(n7891) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n14139), .CK(n5894), .QN(n7906) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n14139), .CK(n5893), .QN(n7896) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n14139), .CK(n5892), .QN(n7902) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n14139), .CK(n5891), .QN(n7883) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n14139), .CK(n5890), .QN(n7881) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n14139), .CK(n5888), .QN(n7888) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n14139), .CK(n5887), .QN(n7909) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n14139), .CK(n5886), .QN(n7890) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n14139), .CK(n5885), .QN(n7901) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n14139), .CK(n5884), .QN(n7885) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n14139), .CK(n5883), .QN(n7886) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n14139), .CK(n5882), .QN(n7911) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n32728), .CK(n5881), .QN(n7889) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n32728), .CK(n5880), .QN(n7887) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n32728), .CK(n5879), .QN(n7899) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n14139), .CK(n5909), .QN(n7897) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n14139), .CK(n5908), .QN(n7904) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n32728), .CK(n5907), .QN(n7908) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n32728), .CK(n5906), .QN(n7884) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n32728), .CK(n5905), .QN(n7910) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n32728), .CK(n5904), .QN(n7905) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n32728), .CK(n5903), .QN(n7903) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n32728), .CK(n5900), .QN(n7898) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n32728), .CK(n5889), .QN(n7900) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n14139), .CK(n5878), .QN(n7912) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n14138), .CK(n5902), .QN(n7861) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n14138), .CK(n5901), .QN(n7860) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n32729), .CK(n5899), .QN(n7862) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n14138), .CK(n5898), .QN(n7850) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n14138), .CK(n5897), .QN(n7875) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n14138), .CK(n5896), .QN(n7863) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n32729), .CK(n5895), .QN(n7859) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n32729), .CK(n5894), .QN(n7874) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n32729), .CK(n5893), .QN(n7864) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n14138), .CK(n5892), .QN(n7870) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n14138), .CK(n5891), .QN(n7851) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n14138), .CK(n5890), .QN(n7849) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n14138), .CK(n5888), .QN(n7856) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n32729), .CK(n5887), .QN(n7877) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n32729), .CK(n5886), .QN(n7858) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n32729), .CK(n5885), .QN(n7869) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n14138), .CK(n5884), .QN(n7853) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n32729), .CK(n5883), .QN(n7854) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n32729), .CK(n5882), .QN(n7879) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n32729), .CK(n5881), .QN(n7857) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n14138), .CK(n5880), .QN(n7855) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n14138), .CK(n5879), .QN(n7867) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n32729), .CK(n5909), .QN(n7865) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n32729), .CK(n5908), .QN(n7872) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n32729), .CK(n5907), .QN(n7876) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n14138), .CK(n5906), .QN(n7852) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n14138), .CK(n5905), .QN(n7878) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n14138), .CK(n5904), .QN(n7873) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n14138), .CK(n5903), .QN(n7871) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n14138), .CK(n5900), .QN(n7866) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n32729), .CK(n5889), .QN(n7868) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n14138), .CK(n5878), .QN(n7880) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n14154), .CK(n5902), .QN(n8373) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n14154), .CK(n5901), .QN(n8372) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n14154), .CK(n5899), .QN(n8374) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n14154), .CK(n5898), .QN(n8362) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n14154), .CK(n5897), .QN(n8387) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n14154), .CK(n5896), .QN(n8375) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n14154), .CK(n5895), .QN(n8371) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n14154), .CK(n5894), .QN(n8386) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n14154), .CK(n5893), .QN(n8376) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n14154), .CK(n5892), .QN(n8382) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n14154), .CK(n5891), .QN(n8363) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n14154), .CK(n5890), .QN(n8361) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n14154), .CK(n5888), .QN(n8368) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n14154), .CK(n5887), .QN(n8389) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n14154), .CK(n5886), .QN(n8370) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n14154), .CK(n5885), .QN(n8381) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n14154), .CK(n5884), .QN(n8365) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n14154), .CK(n5883), .QN(n8366) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n14154), .CK(n5882), .QN(n8391) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n14154), .CK(n5881), .QN(n8369) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n14154), .CK(n5880), .QN(n8367) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n14154), .CK(n5879), .QN(n8379) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n14154), .CK(n5909), .QN(n8377) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n14154), .CK(n5908), .QN(n8384) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n14154), .CK(n5907), .QN(n8388) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n14154), .CK(n5906), .QN(n8364) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n14154), .CK(n5905), .QN(n8390) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n14154), .CK(n5904), .QN(n8385) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n14154), .CK(n5903), .QN(n8383) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n14154), .CK(n5900), .QN(n8378) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n14154), .CK(n5889), .QN(n8380) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n14154), .CK(n5878), .QN(n8392) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n14155), .CK(n5902), .QN(n8405) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n14155), .CK(n5901), .QN(n8404) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n14155), .CK(n5899), .QN(n8406) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n14155), .CK(n5898), .QN(n8394) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n14155), .CK(n5897), .QN(n8419) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n14155), .CK(n5896), .QN(n8407) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n14155), .CK(n5895), .QN(n8403) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n14155), .CK(n5894), .QN(n8418) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n14155), .CK(n5893), .QN(n8408) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n14155), .CK(n5892), .QN(n8414) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n14155), .CK(n5891), .QN(n8395) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n14155), .CK(n5890), .QN(n8393) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n14155), .CK(n5888), .QN(n8400) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n14155), .CK(n5887), .QN(n8421) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n14155), .CK(n5886), .QN(n8402) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n14155), .CK(n5885), .QN(n8413) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n14155), .CK(n5884), .QN(n8397) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n14155), .CK(n5883), .QN(n8398) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n14155), .CK(n5882), .QN(n8423) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n14155), .CK(n5881), .QN(n8401) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n14155), .CK(n5880), .QN(n8399) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n14155), .CK(n5879), .QN(n8411) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n14155), .CK(n5909), .QN(n8409) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n14155), .CK(n5908), .QN(n8416) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n14155), .CK(n5907), .QN(n8420) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n14155), .CK(n5906), .QN(n8396) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n14155), .CK(n5905), .QN(n8422) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n14155), .CK(n5904), .QN(n8417) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n14155), .CK(n5903), .QN(n8415) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n14155), .CK(n5900), .QN(n8410) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n14155), .CK(n5889), .QN(n8412) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n14155), .CK(n5878), .QN(n8424) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n14149), .CK(n5902), .QN(n8213) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n14149), .CK(n5901), .QN(n8212) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n14149), .CK(n5899), .QN(n8214) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n14149), .CK(n5898), .QN(n8202) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n14149), .CK(n5897), .QN(n8227) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n14149), .CK(n5896), .QN(n8215) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n14149), .CK(n5895), .QN(n8211) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n14149), .CK(n5894), .QN(n8226) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n14149), .CK(n5893), .QN(n8216) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n14149), .CK(n5892), .QN(n8222) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n14149), .CK(n5891), .QN(n8203) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n14149), .CK(n5890), .QN(n8201) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n14149), .CK(n5888), .QN(n8208) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n14149), .CK(n5887), .QN(n8229) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n14149), .CK(n5886), .QN(n8210) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n14149), .CK(n5885), .QN(n8221) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n14149), .CK(n5884), .QN(n8205) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n14149), .CK(n5883), .QN(n8206) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n14149), .CK(n5882), .QN(n8231) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n14149), .CK(n5881), .QN(n8209) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n14149), .CK(n5880), .QN(n8207) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n14149), .CK(n5879), .QN(n8219) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n14149), .CK(n5909), .QN(n8217) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n14149), .CK(n5908), .QN(n8224) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n14149), .CK(n5907), .QN(n8228) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n14149), .CK(n5906), .QN(n8204) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n14149), .CK(n5905), .QN(n8230) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n14149), .CK(n5904), .QN(n8225) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n14149), .CK(n5903), .QN(n8223) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n14149), .CK(n5900), .QN(n8218) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n14149), .CK(n5889), .QN(n8220) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n14149), .CK(n5878), .QN(n8232) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n14151), .CK(n5902), .QN(n8277) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n14153), .CK(n5902), .QN(n8341) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n14151), .CK(n5901), .QN(n8276) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n14153), .CK(n5901), .QN(n8340) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n14151), .CK(n5899), .QN(n8278) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n14153), .CK(n5899), .QN(n8342) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n14151), .CK(n5898), .QN(n8266) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n14153), .CK(n5898), .QN(n8330) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n14151), .CK(n5897), .QN(n8291) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n14153), .CK(n5897), .QN(n8355) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n14151), .CK(n5896), .QN(n8279) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n14153), .CK(n5896), .QN(n8343) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n14151), .CK(n5895), .QN(n8275) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n14153), .CK(n5895), .QN(n8339) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n14151), .CK(n5894), .QN(n8290) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n14153), .CK(n5894), .QN(n8354) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n14151), .CK(n5893), .QN(n8280) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n14153), .CK(n5893), .QN(n8344) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n14151), .CK(n5892), .QN(n8286) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n14153), .CK(n5892), .QN(n8350) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n14151), .CK(n5891), .QN(n8267) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n14153), .CK(n5891), .QN(n8331) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n14151), .CK(n5890), .QN(n8265) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n14153), .CK(n5890), .QN(n8329) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n14151), .CK(n5888), .QN(n8272) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n14153), .CK(n5888), .QN(n8336) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n14151), .CK(n5887), .QN(n8293) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n14153), .CK(n5887), .QN(n8357) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n14151), .CK(n5886), .QN(n8274) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n14153), .CK(n5886), .QN(n8338) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n14151), .CK(n5885), .QN(n8285) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n14153), .CK(n5885), .QN(n8349) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n14151), .CK(n5884), .QN(n8269) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n14153), .CK(n5884), .QN(n8333) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n14151), .CK(n5883), .QN(n8270) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n14153), .CK(n5883), .QN(n8334) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n14151), .CK(n5882), .QN(n8295) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n14153), .CK(n5882), .QN(n8359) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n14151), .CK(n5881), .QN(n8273) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n14153), .CK(n5881), .QN(n8337) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n14151), .CK(n5880), .QN(n8271) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n14153), .CK(n5880), .QN(n8335) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n14151), .CK(n5879), .QN(n8283) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n14153), .CK(n5879), .QN(n8347) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n14151), .CK(n5909), .QN(n8281) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n14153), .CK(n5909), .QN(n8345) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n14151), .CK(n5908), .QN(n8288) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n14153), .CK(n5908), .QN(n8352) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n14151), .CK(n5907), .QN(n8292) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n14153), .CK(n5907), .QN(n8356) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n14151), .CK(n5906), .QN(n8268) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n14153), .CK(n5906), .QN(n8332) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n14151), .CK(n5905), .QN(n8294) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n14153), .CK(n5905), .QN(n8358) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n14151), .CK(n5904), .QN(n8289) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n14153), .CK(n5904), .QN(n8353) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n14151), .CK(n5903), .QN(n8287) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n14153), .CK(n5903), .QN(n8351) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n14151), .CK(n5900), .QN(n8282) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n14153), .CK(n5900), .QN(n8346) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n14151), .CK(n5889), .QN(n8284) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n14153), .CK(n5889), .QN(n8348) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n14151), .CK(n5878), .QN(n8296) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n14153), .CK(n5878), .QN(n8360) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n14150), .CK(n5902), .QN(n8245) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n14152), .CK(n5902), .QN(n8309) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n14150), .CK(n5901), .QN(n8244) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n14152), .CK(n5901), .QN(n8308) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n14150), .CK(n5899), .QN(n8246) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n14152), .CK(n5899), .QN(n8310) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n14150), .CK(n5898), .QN(n8234) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n14152), .CK(n5898), .QN(n8298) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n14150), .CK(n5897), .QN(n8259) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n14152), .CK(n5897), .QN(n8323) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n14150), .CK(n5896), .QN(n8247) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n14152), .CK(n5896), .QN(n8311) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n14150), .CK(n5895), .QN(n8243) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n14152), .CK(n5895), .QN(n8307) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n14150), .CK(n5894), .QN(n8258) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n14152), .CK(n5894), .QN(n8322) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n14150), .CK(n5893), .QN(n8248) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n14152), .CK(n5893), .QN(n8312) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n14150), .CK(n5892), .QN(n8254) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n14152), .CK(n5892), .QN(n8318) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n14150), .CK(n5891), .QN(n8235) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n14152), .CK(n5891), .QN(n8299) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n14150), .CK(n5890), .QN(n8233) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n14152), .CK(n5890), .QN(n8297) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n14150), .CK(n5888), .QN(n8240) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n14152), .CK(n5888), .QN(n8304) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n14150), .CK(n5887), .QN(n8261) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n14152), .CK(n5887), .QN(n8325) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n14150), .CK(n5886), .QN(n8242) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n14152), .CK(n5886), .QN(n8306) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n14150), .CK(n5885), .QN(n8253) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n14152), .CK(n5885), .QN(n8317) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n14150), .CK(n5884), .QN(n8237) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n14152), .CK(n5884), .QN(n8301) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n14150), .CK(n5883), .QN(n8238) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n14152), .CK(n5883), .QN(n8302) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n14150), .CK(n5882), .QN(n8263) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n14152), .CK(n5882), .QN(n8327) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n14150), .CK(n5881), .QN(n8241) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n14152), .CK(n5881), .QN(n8305) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n14150), .CK(n5880), .QN(n8239) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n14152), .CK(n5880), .QN(n8303) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n14150), .CK(n5879), .QN(n8251) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n14152), .CK(n5879), .QN(n8315) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n14150), .CK(n5909), .QN(n8249) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n14152), .CK(n5909), .QN(n8313) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n14150), .CK(n5908), .QN(n8256) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n14152), .CK(n5908), .QN(n8320) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n14150), .CK(n5907), .QN(n8260) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n14152), .CK(n5907), .QN(n8324) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n14150), .CK(n5906), .QN(n8236) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n14152), .CK(n5906), .QN(n8300) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n14150), .CK(n5905), .QN(n8262) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n14152), .CK(n5905), .QN(n8326) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n14150), .CK(n5904), .QN(n8257) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n14152), .CK(n5904), .QN(n8321) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n14150), .CK(n5903), .QN(n8255) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n14152), .CK(n5903), .QN(n8319) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n14150), .CK(n5900), .QN(n8250) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n14152), .CK(n5900), .QN(n8314) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n14150), .CK(n5889), .QN(n8252) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n14152), .CK(n5889), .QN(n8316) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n14150), .CK(n5878), .QN(n8264) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n14152), .CK(n5878), .QN(n8328) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n14137), .CK(n5902), .QN(n7829) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n14137), .CK(n5901), .QN(n7828) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n14137), .CK(n5899), .QN(n7830) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n14137), .CK(n5898), .QN(n7818) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n14137), .CK(n5897), .QN(n7843) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n14137), .CK(n5896), .QN(n7831) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n14137), .CK(n5895), .QN(n7827) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n14137), .CK(n5894), .QN(n7842) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n14137), .CK(n5893), .QN(n7832) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n14137), .CK(n5892), .QN(n7838) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n14137), .CK(n5891), .QN(n7819) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n14137), .CK(n5890), .QN(n7817) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n14137), .CK(n5888), .QN(n7824) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n14137), .CK(n5887), .QN(n7845) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n14137), .CK(n5886), .QN(n7826) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n14137), .CK(n5885), .QN(n7837) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n14137), .CK(n5884), .QN(n7821) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n14137), .CK(n5883), .QN(n7822) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n14137), .CK(n5882), .QN(n7847) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n14137), .CK(n5881), .QN(n7825) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n14137), .CK(n5880), .QN(n7823) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n14137), .CK(n5879), .QN(n7835) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n14137), .CK(n5909), .QN(n7833) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n14137), .CK(n5908), .QN(n7840) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n14137), .CK(n5907), .QN(n7844) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n14137), .CK(n5906), .QN(n7820) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n14137), .CK(n5905), .QN(n7846) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n14137), .CK(n5904), .QN(n7841) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n14137), .CK(n5903), .QN(n7839) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n14137), .CK(n5900), .QN(n7834) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n14137), .CK(n5889), .QN(n7836) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n14137), .CK(n5878), .QN(n7848) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n14134), .CK(n5902), .QN(n7733) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n14134), .CK(n5901), .QN(n7732) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n14134), .CK(n5899), .QN(n7734) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n14134), .CK(n5898), .QN(n7722) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n14134), .CK(n5897), .QN(n7747) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n14134), .CK(n5896), .QN(n7735) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n14134), .CK(n5895), .QN(n7731) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n14134), .CK(n5894), .QN(n7746) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n14134), .CK(n5893), .QN(n7736) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n14134), .CK(n5892), .QN(n7742) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n14134), .CK(n5891), .QN(n7723) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n14134), .CK(n5890), .QN(n7721) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n14134), .CK(n5888), .QN(n7728) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n14134), .CK(n5887), .QN(n7749) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n14134), .CK(n5886), .QN(n7730) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n14134), .CK(n5885), .QN(n7741) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n14134), .CK(n5884), .QN(n7725) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n14134), .CK(n5883), .QN(n7726) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n14134), .CK(n5882), .QN(n7751) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n14134), .CK(n5881), .QN(n7729) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n14134), .CK(n5880), .QN(n7727) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n14134), .CK(n5879), .QN(n7739) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n14134), .CK(n5909), .QN(n7737) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n14134), .CK(n5908), .QN(n7744) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n14134), .CK(n5907), .QN(n7748) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n14134), .CK(n5906), .QN(n7724) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n14134), .CK(n5905), .QN(n7750) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n14134), .CK(n5904), .QN(n7745) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n14134), .CK(n5903), .QN(n7743) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n14134), .CK(n5900), .QN(n7738) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n14134), .CK(n5889), .QN(n7740) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n14134), .CK(n5878), .QN(n7752) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n14136), .CK(n5902), .QN(n7797) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n14136), .CK(n5901), .QN(n7796) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n14136), .CK(n5899), .QN(n7798) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n14136), .CK(n5898), .QN(n7786) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n14136), .CK(n5897), .QN(n7811) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n14136), .CK(n5896), .QN(n7799) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n14136), .CK(n5895), .QN(n7795) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n14136), .CK(n5894), .QN(n7810) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n14136), .CK(n5893), .QN(n7800) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n14136), .CK(n5892), .QN(n7806) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n14136), .CK(n5891), .QN(n7787) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n14136), .CK(n5890), .QN(n7785) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n14136), .CK(n5888), .QN(n7792) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n14136), .CK(n5887), .QN(n7813) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n14136), .CK(n5886), .QN(n7794) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n14136), .CK(n5885), .QN(n7805) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n14136), .CK(n5884), .QN(n7789) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n14136), .CK(n5883), .QN(n7790) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n14136), .CK(n5882), .QN(n7815) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n14136), .CK(n5881), .QN(n7793) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n14136), .CK(n5880), .QN(n7791) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n14136), .CK(n5879), .QN(n7803) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n14136), .CK(n5909), .QN(n7801) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n14136), .CK(n5908), .QN(n7808) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n14136), .CK(n5907), .QN(n7812) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n14136), .CK(n5906), .QN(n7788) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n14136), .CK(n5905), .QN(n7814) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n14136), .CK(n5904), .QN(n7809) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n14136), .CK(n5903), .QN(n7807) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n14136), .CK(n5900), .QN(n7802) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n14136), .CK(n5889), .QN(n7804) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n14136), .CK(n5878), .QN(n7816) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n32730), .CK(n5902), .QN(n7701) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n32730), .CK(n5901), .QN(n7700) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n14133), .CK(n5899), .QN(n7702) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n32730), .CK(n5898), .QN(n7690) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n32730), .CK(n5897), .QN(n7715) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n32730), .CK(n5896), .QN(n7703) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n32730), .CK(n5895), .QN(n7699) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n32730), .CK(n5894), .QN(n7714) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n14133), .CK(n5893), .QN(n7704) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n32730), .CK(n5892), .QN(n7710) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n32730), .CK(n5891), .QN(n7691) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n14133), .CK(n5890), .QN(n7689) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n32730), .CK(n5888), .QN(n7696) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n14133), .CK(n5887), .QN(n7717) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n14133), .CK(n5886), .QN(n7698) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n14133), .CK(n5885), .QN(n7709) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n14133), .CK(n5884), .QN(n7693) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n14133), .CK(n5883), .QN(n7694) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n32730), .CK(n5882), .QN(n7719) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n14133), .CK(n5881), .QN(n7697) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n14133), .CK(n5880), .QN(n7695) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n32730), .CK(n5879), .QN(n7707) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n32730), .CK(n5909), .QN(n7705) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n14133), .CK(n5908), .QN(n7712) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n14133), .CK(n5907), .QN(n7716) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n14133), .CK(n5906), .QN(n7692) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n14133), .CK(n5905), .QN(n7718) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n14133), .CK(n5904), .QN(n7713) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n14133), .CK(n5903), .QN(n7711) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n14133), .CK(n5900), .QN(n7706) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n14133), .CK(n5889), .QN(n7708) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n32730), .CK(n5878), .QN(n7720) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n14135), .CK(n5902), .QN(n7765) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n14135), .CK(n5901), .QN(n7764) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n14135), .CK(n5899), .QN(n7766) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n14135), .CK(n5898), .QN(n7754) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n14135), .CK(n5897), .QN(n7779) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n14135), .CK(n5896), .QN(n7767) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n14135), .CK(n5895), .QN(n7763) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n14135), .CK(n5894), .QN(n7778) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n14135), .CK(n5893), .QN(n7768) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n14135), .CK(n5892), .QN(n7774) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n14135), .CK(n5891), .QN(n7755) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n14135), .CK(n5890), .QN(n7753) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n14135), .CK(n5888), .QN(n7760) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n14135), .CK(n5887), .QN(n7781) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n14135), .CK(n5886), .QN(n7762) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n14135), .CK(n5885), .QN(n7773) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n14135), .CK(n5884), .QN(n7757) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n14135), .CK(n5883), .QN(n7758) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n14135), .CK(n5882), .QN(n7783) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n14135), .CK(n5881), .QN(n7761) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n14135), .CK(n5880), .QN(n7759) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n14135), .CK(n5879), .QN(n7771) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n14135), .CK(n5909), .QN(n7769) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n14135), .CK(n5908), .QN(n7776) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n14135), .CK(n5907), .QN(n7780) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n14135), .CK(n5906), .QN(n7756) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n14135), .CK(n5905), .QN(n7782) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n14135), .CK(n5904), .QN(n7777) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n14135), .CK(n5903), .QN(n7775) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n14135), .CK(n5900), .QN(n7770) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n14135), .CK(n5889), .QN(n7772) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n14135), .CK(n5878), .QN(n7784) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n14132), .CK(n5902), .QN(n7669) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n14132), .CK(n5901), .QN(n7668) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n14132), .CK(n5899), .QN(n7670) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n14132), .CK(n5898), .QN(n7658) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n14132), .CK(n5897), .QN(n7683) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n14132), .CK(n5896), .QN(n7671) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n14132), .CK(n5895), .QN(n7667) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n14132), .CK(n5894), .QN(n7682) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n14132), .CK(n5893), .QN(n7672) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n14132), .CK(n5892), .QN(n7678) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n14132), .CK(n5891), .QN(n7659) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n14132), .CK(n5890), .QN(n7657) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n14132), .CK(n5888), .QN(n7664) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n14132), .CK(n5887), .QN(n7685) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n14132), .CK(n5886), .QN(n7666) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n14132), .CK(n5885), .QN(n7677) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n14132), .CK(n5884), .QN(n7661) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n14132), .CK(n5883), .QN(n7662) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n14132), .CK(n5882), .QN(n7687) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n14132), .CK(n5881), .QN(n7665) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n14132), .CK(n5880), .QN(n7663) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n14132), .CK(n5879), .QN(n7675) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n14132), .CK(n5909), .QN(n7673) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n14132), .CK(n5908), .QN(n7680) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n14132), .CK(n5907), .QN(n7684) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n14132), .CK(n5906), .QN(n7660) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n14132), .CK(n5905), .QN(n7686) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n14132), .CK(n5904), .QN(n7681) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n14132), .CK(n5903), .QN(n7679) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n14132), .CK(n5900), .QN(n7674) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n14132), .CK(n5889), .QN(n7676) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n14132), .CK(n5878), .QN(n7688) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n14131), .CK(n5902), .QN(n7637) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n14131), .CK(n5901), .QN(n7636) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n14131), .CK(n5899), .QN(n7638) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n14131), .CK(n5898), .QN(n7626) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n14131), .CK(n5897), .QN(n7651) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n14131), .CK(n5896), .QN(n7639) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n14131), .CK(n5895), .QN(n7635) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n14131), .CK(n5894), .QN(n7650) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n14131), .CK(n5893), .QN(n7640) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n14131), .CK(n5892), .QN(n7646) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n14131), .CK(n5891), .QN(n7627) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n14131), .CK(n5890), .QN(n7625) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n14131), .CK(n5888), .QN(n7632) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n14131), .CK(n5887), .QN(n7653) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n14131), .CK(n5886), .QN(n7634) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n14131), .CK(n5885), .QN(n7645) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n14131), .CK(n5884), .QN(n7629) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n14131), .CK(n5883), .QN(n7630) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n14131), .CK(n5882), .QN(n7655) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n14131), .CK(n5881), .QN(n7633) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n14131), .CK(n5880), .QN(n7631) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n14131), .CK(n5879), .QN(n7643) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n14131), .CK(n5909), .QN(n7641) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n14131), .CK(n5908), .QN(n7648) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n14131), .CK(n5907), .QN(n7652) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n14131), .CK(n5906), .QN(n7628) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n14131), .CK(n5905), .QN(n7654) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n14131), .CK(n5904), .QN(n7649) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n14131), .CK(n5903), .QN(n7647) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n14131), .CK(n5900), .QN(n7642) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n14131), .CK(n5889), .QN(n7644) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n14131), .CK(n5878), .QN(n7656) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n14130), .CK(n5902), .QN(n7605) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n14130), .CK(n5901), .QN(n7604) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n14130), .CK(n5899), .QN(n7606) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n14130), .CK(n5898), .QN(n7594) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n14130), .CK(n5897), .QN(n7619) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n14130), .CK(n5896), .QN(n7607) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n14130), .CK(n5895), .QN(n7603) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n14130), .CK(n5894), .QN(n7618) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n14130), .CK(n5893), .QN(n7608) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n14130), .CK(n5892), .QN(n7614) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n14130), .CK(n5891), .QN(n7595) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n14130), .CK(n5890), .QN(n7593) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n14130), .CK(n5888), .QN(n7600) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n14130), .CK(n5887), .QN(n7621) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n14130), .CK(n5886), .QN(n7602) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n14130), .CK(n5885), .QN(n7613) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n14130), .CK(n5884), .QN(n7597) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n14130), .CK(n5883), .QN(n7598) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n14130), .CK(n5882), .QN(n7623) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n14130), .CK(n5881), .QN(n7601) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n14130), .CK(n5880), .QN(n7599) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n14130), .CK(n5879), .QN(n7611) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n14130), .CK(n5909), .QN(n7609) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n14130), .CK(n5908), .QN(n7616) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n14130), .CK(n5907), .QN(n7620) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n14130), .CK(n5906), .QN(n7596) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n14130), .CK(n5905), .QN(n7622) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n14130), .CK(n5904), .QN(n7617) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n14130), .CK(n5903), .QN(n7615) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n14130), .CK(n5900), .QN(n7610) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n14130), .CK(n5889), .QN(n7612) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n14130), .CK(n5878), .QN(n7624) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n20327), .CK(n5902), .QN(n7573) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n20327), .CK(n5901), .QN(n7572) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n20327), .CK(n5899), .QN(n7574) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n20327), .CK(n5898), .QN(n7562) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n20327), .CK(n5897), .QN(n7587) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n20327), .CK(n5896), .QN(n7575) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n20327), .CK(n5895), .QN(n7571) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n20327), .CK(n5894), .QN(n7586) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n20327), .CK(n5893), .QN(n7576) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n20327), .CK(n5892), .QN(n7582) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n20327), .CK(n5891), .QN(n7563) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n20327), .CK(n5890), .QN(n7561) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n20327), .CK(n5888), .QN(n7568) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n20327), .CK(n5887), .QN(n7589) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n20327), .CK(n5886), .QN(n7570) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n20327), .CK(n5885), .QN(n7581) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n20327), .CK(n5884), .QN(n7565) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n20327), .CK(n5883), .QN(n7566) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n20327), .CK(n5882), .QN(n7591) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n20327), .CK(n5881), .QN(n7569) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n20327), .CK(n5880), .QN(n7567) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n20327), .CK(n5879), .QN(n7579) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n20327), .CK(n5909), .QN(n7577) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n20327), .CK(n5908), .QN(n7584) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n20327), .CK(n5907), .QN(n7588) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n20327), .CK(n5906), .QN(n7564) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n20327), .CK(n5905), .QN(n7590) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n20327), .CK(n5904), .QN(n7585) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n20327), .CK(n5903), .QN(n7583) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n20327), .CK(n5900), .QN(n7578) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n20327), .CK(n5889), .QN(n7580) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n20327), .CK(n5878), .QN(n7592) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n32723), .CK(n5902), .QN(n7541) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n32723), .CK(n5901), .QN(n7540) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n32723), .CK(n5899), .QN(n7542) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n32723), .CK(n5898), .QN(n7530) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n32723), .CK(n5897), .QN(n7555) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n32723), .CK(n5896), .QN(n7543) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n32723), .CK(n5895), .QN(n7539) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n32723), .CK(n5894), .QN(n7554) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n32723), .CK(n5893), .QN(n7544) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n32723), .CK(n5892), .QN(n7550) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n32723), .CK(n5891), .QN(n7531) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n32723), .CK(n5890), .QN(n7529) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n32723), .CK(n5888), .QN(n7536) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n32723), .CK(n5887), .QN(n7557) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n32723), .CK(n5886), .QN(n7538) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n32723), .CK(n5885), .QN(n7549) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n32723), .CK(n5884), .QN(n7533) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n32723), .CK(n5883), .QN(n7534) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n32723), .CK(n5882), .QN(n7559) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n32723), .CK(n5881), .QN(n7537) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n32723), .CK(n5880), .QN(n7535) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n32723), .CK(n5879), .QN(n7547) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n32723), .CK(n5909), .QN(n7545) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n32723), .CK(n5908), .QN(n7552) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n32723), .CK(n5907), .QN(n7556) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n32723), .CK(n5906), .QN(n7532) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n32723), .CK(n5905), .QN(n7558) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n32723), .CK(n5904), .QN(n7553) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n32723), .CK(n5903), .QN(n7551) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n32723), .CK(n5900), .QN(n7546) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n32723), .CK(n5889), .QN(n7548) );
  DFF_X1 \OUT1_reg[30]  ( .D(n5778), .CK(n5809), .Q(OUT1[30]) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n32725), .CK(n5904), .Q(n7425) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n32725), .CK(n5880), .Q(n7407) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n32725), .CK(n5884), .Q(n7405) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n32724), .CK(n5909), .Q(n7417) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n32725), .CK(n5879), .Q(n7419) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n32724), .CK(n5883), .Q(n7406) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n32724), .CK(n5885), .Q(n7421) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n32725), .CK(n5891), .Q(n7403) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n32725), .CK(n5893), .Q(n7416) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n32725), .CK(n5902), .Q(n7413) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n32725), .CK(n5895), .Q(n7411) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n32724), .CK(n5901), .Q(n7412) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n5913), .CK(n5894), .Q(n7426) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n32724), .CK(n5898), .Q(n7402) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n32725), .CK(n5908), .Q(n7424) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n32725), .CK(n5906), .Q(n7404) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n32724), .CK(n5896), .Q(n7415) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n32724), .CK(n5897), .Q(n7427) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n32724), .CK(n5881), .Q(n7409) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n32724), .CK(n5903), .Q(n7423) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n32724), .CK(n5889), .Q(n7420) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n32724), .CK(n5890), .Q(n7401) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n32724), .CK(n5886), .Q(n7410) );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n32724), .CK(n5878), .Q(n7432) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n32724), .CK(n5888), .Q(n7408) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n32724), .CK(n5892), .Q(n7422) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n32724), .CK(n5882), .Q(n7431) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n32724), .CK(n5907), .Q(n7428) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n32725), .CK(n5887), .Q(n7429) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n32724), .CK(n5905), .Q(n7430) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n32724), .CK(n5899), .Q(n7414) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n5913), .CK(n5900), .Q(n7418) );
  BUF_X2 U3844 ( .A(n5913), .Z(n32724) );
  NAND2_X2 U3845 ( .A1(RST), .A2(DATAIN[5]), .ZN(n14150) );
  NAND2_X2 U3846 ( .A1(RST), .A2(DATAIN[0]), .ZN(n14155) );
  NAND2_X2 U3847 ( .A1(RST), .A2(DATAIN[7]), .ZN(n14148) );
  INV_X4 U3848 ( .A(n34216), .ZN(n5910) );
  INV_X4 U3849 ( .A(n34214), .ZN(n5912) );
  INV_X4 U3850 ( .A(n34215), .ZN(n5911) );
  BUF_X2 U3851 ( .A(n5913), .Z(n32725) );
  BUF_X2 U3852 ( .A(n34210), .Z(n32665) );
  NAND2_X2 U3853 ( .A1(RST), .A2(DATAIN[1]), .ZN(n14154) );
  NAND2_X2 U3854 ( .A1(RST), .A2(DATAIN[3]), .ZN(n14152) );
  NAND2_X2 U3855 ( .A1(RST), .A2(DATAIN[2]), .ZN(n14153) );
  AND2_X1 U3856 ( .A1(RST), .A2(DATAIN[27]), .ZN(n32683) );
  BUF_X1 U3857 ( .A(n14133), .Z(n32730) );
  NAND2_X2 U3858 ( .A1(RST), .A2(DATAIN[18]), .ZN(n14137) );
  BUF_X1 U3859 ( .A(n14138), .Z(n32729) );
  NAND2_X2 U3860 ( .A1(RST), .A2(DATAIN[21]), .ZN(n14134) );
  NAND2_X2 U3861 ( .A1(RST), .A2(DATAIN[20]), .ZN(n14135) );
  NAND2_X2 U3862 ( .A1(RST), .A2(DATAIN[15]), .ZN(n14140) );
  NAND2_X2 U3863 ( .A1(RST), .A2(DATAIN[19]), .ZN(n14136) );
  NAND2_X2 U3864 ( .A1(RST), .A2(DATAIN[14]), .ZN(n14141) );
  NAND2_X2 U3865 ( .A1(RST), .A2(DATAIN[13]), .ZN(n14142) );
  NAND2_X2 U3866 ( .A1(RST), .A2(DATAIN[12]), .ZN(n14143) );
  NAND2_X2 U3867 ( .A1(RST), .A2(DATAIN[10]), .ZN(n14145) );
  NAND2_X2 U3868 ( .A1(RST), .A2(DATAIN[11]), .ZN(n14144) );
  OR2_X1 U3869 ( .A1(n33498), .A2(n33499), .ZN(n34173) );
  BUF_X2 U3870 ( .A(n34186), .Z(n32666) );
  OR2_X1 U3871 ( .A1(n33498), .A2(n33504), .ZN(n34181) );
  OR2_X1 U3872 ( .A1(n33493), .A2(n33500), .ZN(n34175) );
  OR2_X1 U3873 ( .A1(n33502), .A2(n33506), .ZN(n34163) );
  OR2_X1 U3874 ( .A1(n33493), .A2(n33504), .ZN(n34164) );
  BUF_X2 U3875 ( .A(n34162), .Z(n32667) );
  OR2_X1 U3876 ( .A1(n33498), .A2(n33505), .ZN(n34159) );
  OR2_X1 U3877 ( .A1(n33506), .A2(n33486), .ZN(n34160) );
  OR2_X1 U3878 ( .A1(n33500), .A2(n33506), .ZN(n34157) );
  OR2_X1 U3879 ( .A1(n33493), .A2(n33486), .ZN(n34174) );
  OR2_X1 U3880 ( .A1(n33505), .A2(n33501), .ZN(n34172) );
  OR2_X1 U3881 ( .A1(n33506), .A2(n33503), .ZN(n34197) );
  OR2_X1 U3882 ( .A1(n33500), .A2(n33501), .ZN(n34195) );
  OR2_X1 U3883 ( .A1(n33506), .A2(n33499), .ZN(n34187) );
  OR2_X1 U3884 ( .A1(n33501), .A2(n33499), .ZN(n34196) );
  OR2_X1 U3885 ( .A1(n33493), .A2(n33503), .ZN(n34188) );
  NAND2_X2 U3886 ( .A1(n32791), .A2(n5811), .ZN(n33475) );
  NAND2_X2 U3887 ( .A1(RST), .A2(n32790), .ZN(n33476) );
  NAND2_X2 U3888 ( .A1(RST), .A2(DATAIN[4]), .ZN(n14151) );
  NAND2_X2 U3889 ( .A1(RST), .A2(DATAIN[6]), .ZN(n14149) );
  INV_X2 U3890 ( .A(n34197), .ZN(n32668) );
  INV_X2 U3891 ( .A(n34195), .ZN(n32669) );
  INV_X2 U3892 ( .A(n34187), .ZN(n32670) );
  NOR2_X4 U3893 ( .A1(n33493), .A2(n33492), .ZN(n34185) );
  NOR2_X4 U3894 ( .A1(n33501), .A2(n33492), .ZN(n34183) );
  INV_X2 U3895 ( .A(n34181), .ZN(n32671) );
  INV_X2 U3896 ( .A(n34175), .ZN(n32672) );
  INV_X2 U3897 ( .A(n34173), .ZN(n32673) );
  INV_X2 U3898 ( .A(n34163), .ZN(n32674) );
  NOR2_X4 U3899 ( .A1(n33498), .A2(n33492), .ZN(n34161) );
  INV_X2 U3900 ( .A(n34159), .ZN(n32675) );
  INV_X2 U3901 ( .A(n34157), .ZN(n32676) );
  INV_X2 U3902 ( .A(n34164), .ZN(n32677) );
  INV_X2 U3903 ( .A(n34160), .ZN(n32678) );
  INV_X2 U3904 ( .A(n34174), .ZN(n32679) );
  INV_X2 U3905 ( .A(n34172), .ZN(n32680) );
  NOR2_X4 U3906 ( .A1(n33506), .A2(n33492), .ZN(n34184) );
  NOR2_X4 U3907 ( .A1(n33501), .A2(n33503), .ZN(n34182) );
  INV_X2 U3908 ( .A(n34196), .ZN(n32681) );
  INV_X2 U3909 ( .A(n34188), .ZN(n32682) );
  NOR2_X4 U3910 ( .A1(n33493), .A2(n33499), .ZN(n34170) );
  NOR2_X4 U3911 ( .A1(n33502), .A2(n33501), .ZN(n34198) );
  NOR2_X4 U3912 ( .A1(n33506), .A2(n33504), .ZN(n34200) );
  NOR2_X4 U3913 ( .A1(n33498), .A2(n33503), .ZN(n34194) );
  NAND2_X2 U3914 ( .A1(RST), .A2(DATAIN[23]), .ZN(n14132) );
  BUF_X1 U3915 ( .A(n14139), .Z(n32728) );
  BUF_X1 U3916 ( .A(n14146), .Z(n32727) );
  BUF_X1 U3917 ( .A(n14147), .Z(n32726) );
  BUF_X1 U3918 ( .A(n34199), .Z(n32721) );
  BUF_X1 U3919 ( .A(n34169), .Z(n32717) );
  BUF_X1 U3920 ( .A(n34158), .Z(n32716) );
  BUF_X1 U3921 ( .A(n34176), .Z(n32719) );
  BUF_X1 U3922 ( .A(n34193), .Z(n32720) );
  BUF_X1 U3923 ( .A(n34171), .Z(n32718) );
  INV_X1 U3924 ( .A(ADD_WR[0]), .ZN(n33520) );
  INV_X1 U3925 ( .A(ADD_WR[1]), .ZN(n33521) );
  INV_X1 U3926 ( .A(ADD_WR[2]), .ZN(n33519) );
  INV_X1 U3927 ( .A(ADD_WR[3]), .ZN(n33516) );
  BUF_X1 U3928 ( .A(n33465), .Z(n32714) );
  BUF_X1 U3929 ( .A(n33466), .Z(n32715) );
  BUF_X1 U3930 ( .A(n33464), .Z(n32713) );
  BUF_X1 U3931 ( .A(n33462), .Z(n32711) );
  BUF_X1 U3932 ( .A(n33460), .Z(n32709) );
  BUF_X1 U3933 ( .A(n33453), .Z(n32706) );
  BUF_X1 U3934 ( .A(n33454), .Z(n32707) );
  BUF_X1 U3935 ( .A(n33451), .Z(n32704) );
  BUF_X1 U3936 ( .A(n33452), .Z(n32705) );
  BUF_X1 U3937 ( .A(n33449), .Z(n32702) );
  BUF_X1 U3938 ( .A(n33450), .Z(n32703) );
  BUF_X1 U3939 ( .A(n33447), .Z(n32700) );
  BUF_X1 U3940 ( .A(n33448), .Z(n32701) );
  BUF_X1 U3941 ( .A(n33441), .Z(n32698) );
  BUF_X1 U3942 ( .A(n33442), .Z(n32699) );
  BUF_X1 U3943 ( .A(n33439), .Z(n32696) );
  BUF_X1 U3944 ( .A(n33440), .Z(n32697) );
  BUF_X1 U3945 ( .A(n33437), .Z(n32694) );
  BUF_X1 U3946 ( .A(n33438), .Z(n32695) );
  BUF_X1 U3947 ( .A(n33435), .Z(n32692) );
  BUF_X1 U3948 ( .A(n33436), .Z(n32693) );
  BUF_X1 U3949 ( .A(n33430), .Z(n32691) );
  BUF_X1 U3950 ( .A(n33428), .Z(n32689) );
  BUF_X1 U3951 ( .A(n33425), .Z(n32686) );
  BUF_X1 U3952 ( .A(n33426), .Z(n32687) );
  BUF_X1 U3953 ( .A(n33424), .Z(n32685) );
  NAND2_X1 U3954 ( .A1(RST), .A2(DATAIN[22]), .ZN(n14133) );
  INV_X1 U3955 ( .A(ADD_WR[4]), .ZN(n33517) );
  BUF_X1 U3956 ( .A(n33463), .Z(n32712) );
  BUF_X1 U3957 ( .A(n33461), .Z(n32710) );
  BUF_X1 U3958 ( .A(n33459), .Z(n32708) );
  BUF_X1 U3959 ( .A(n33429), .Z(n32690) );
  BUF_X1 U3960 ( .A(n33427), .Z(n32688) );
  BUF_X1 U3961 ( .A(n33423), .Z(n32684) );
  NAND2_X1 U3962 ( .A1(RST), .A2(DATAIN[16]), .ZN(n14139) );
  NAND2_X1 U3963 ( .A1(RST), .A2(DATAIN[8]), .ZN(n14147) );
  NAND2_X1 U3964 ( .A1(RST), .A2(DATAIN[17]), .ZN(n14138) );
  NAND2_X1 U3965 ( .A1(RST), .A2(DATAIN[9]), .ZN(n14146) );
  BUF_X2 U3966 ( .A(n34209), .Z(n32722) );
  NAND2_X2 U3967 ( .A1(RST), .A2(DATAIN[24]), .ZN(n14131) );
  NAND2_X2 U3968 ( .A1(RST), .A2(DATAIN[25]), .ZN(n14130) );
  NAND2_X2 U3969 ( .A1(RST), .A2(DATAIN[26]), .ZN(n20327) );
  INV_X2 U3970 ( .A(n32683), .ZN(n32723) );
  NAND4_X1 U3971 ( .A1(EN), .A2(RST), .A3(RD2), .A4(n34209), .ZN(n34210) );
  NOR2_X1 U3972 ( .A1(n33506), .A2(n33505), .ZN(n34199) );
  NOR2_X1 U3973 ( .A1(n33502), .A2(n33498), .ZN(n34176) );
  NOR2_X1 U3974 ( .A1(n33493), .A2(n33505), .ZN(n34171) );
  NOR2_X1 U3975 ( .A1(n33493), .A2(n33502), .ZN(n34158) );
  NAND2_X1 U3976 ( .A1(WR), .A2(EN), .ZN(n32731) );
  NOR2_X1 U3977 ( .A1(n33516), .A2(n32731), .ZN(n32733) );
  NAND2_X1 U3978 ( .A1(ADD_WR[4]), .A2(n32733), .ZN(n32745) );
  NAND3_X1 U3979 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(ADD_WR[1]), .ZN(n32740)
         );
  OAI21_X1 U3980 ( .B1(n32745), .B2(n32740), .A(RST), .ZN(n1045) );
  NAND3_X1 U3981 ( .A1(ADD_WR[2]), .A2(ADD_WR[1]), .A3(n33520), .ZN(n32738) );
  OAI21_X1 U3982 ( .B1(n32745), .B2(n32738), .A(RST), .ZN(n1046) );
  NAND3_X1 U3983 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(n33519), .ZN(n32737) );
  OAI21_X1 U3984 ( .B1(n32745), .B2(n32737), .A(RST), .ZN(n1047) );
  NAND3_X1 U3985 ( .A1(ADD_WR[1]), .A2(n33520), .A3(n33519), .ZN(n32736) );
  OAI21_X1 U3986 ( .B1(n32745), .B2(n32736), .A(RST), .ZN(n1048) );
  NOR2_X1 U3987 ( .A1(ADD_WR[3]), .A2(n32731), .ZN(n32735) );
  NAND2_X1 U3988 ( .A1(ADD_WR[4]), .A2(n32735), .ZN(n32732) );
  OAI21_X1 U3989 ( .B1(n32740), .B2(n32732), .A(RST), .ZN(n1049) );
  OAI21_X1 U3990 ( .B1(n32738), .B2(n32732), .A(RST), .ZN(n1050) );
  NAND3_X1 U3991 ( .A1(ADD_WR[2]), .A2(ADD_WR[0]), .A3(n33521), .ZN(n32744) );
  OAI21_X1 U3992 ( .B1(n32732), .B2(n32744), .A(RST), .ZN(n1051) );
  NAND3_X1 U3993 ( .A1(ADD_WR[2]), .A2(n33520), .A3(n33521), .ZN(n32743) );
  OAI21_X1 U3994 ( .B1(n32732), .B2(n32743), .A(RST), .ZN(n1052) );
  OAI21_X1 U3995 ( .B1(n32737), .B2(n32732), .A(RST), .ZN(n1053) );
  OAI21_X1 U3996 ( .B1(n32736), .B2(n32732), .A(RST), .ZN(n1054) );
  NAND3_X1 U3997 ( .A1(ADD_WR[0]), .A2(n33519), .A3(n33521), .ZN(n32742) );
  OAI21_X1 U3998 ( .B1(n32732), .B2(n32742), .A(RST), .ZN(n1055) );
  NAND3_X1 U3999 ( .A1(n33520), .A2(n33519), .A3(n33521), .ZN(n32741) );
  OAI21_X1 U4000 ( .B1(n32732), .B2(n32741), .A(RST), .ZN(n1056) );
  NAND2_X1 U4001 ( .A1(n32733), .A2(n33517), .ZN(n32734) );
  OAI21_X1 U4002 ( .B1(n32740), .B2(n32734), .A(RST), .ZN(n1057) );
  OAI21_X1 U4003 ( .B1(n32738), .B2(n32734), .A(RST), .ZN(n1058) );
  OAI21_X1 U4004 ( .B1(n32744), .B2(n32734), .A(RST), .ZN(n1059) );
  OAI21_X1 U4005 ( .B1(n32743), .B2(n32734), .A(RST), .ZN(n1060) );
  OAI21_X1 U4006 ( .B1(n32737), .B2(n32734), .A(RST), .ZN(n1061) );
  OAI21_X1 U4007 ( .B1(n32736), .B2(n32734), .A(RST), .ZN(n1062) );
  OAI21_X1 U4008 ( .B1(n32742), .B2(n32734), .A(RST), .ZN(n1063) );
  OAI21_X1 U4009 ( .B1(n32741), .B2(n32734), .A(RST), .ZN(n1064) );
  NAND2_X1 U4010 ( .A1(n32735), .A2(n33517), .ZN(n32739) );
  OAI21_X1 U4011 ( .B1(n32744), .B2(n32739), .A(RST), .ZN(n1065) );
  OAI21_X1 U4012 ( .B1(n32743), .B2(n32739), .A(RST), .ZN(n1066) );
  OAI21_X1 U4013 ( .B1(n32742), .B2(n32739), .A(RST), .ZN(n1067) );
  OAI21_X1 U4014 ( .B1(n32741), .B2(n32739), .A(RST), .ZN(n1068) );
  OAI21_X1 U4015 ( .B1(n32736), .B2(n32739), .A(RST), .ZN(n1069) );
  OAI21_X1 U4016 ( .B1(n32737), .B2(n32739), .A(RST), .ZN(n1070) );
  OAI21_X1 U4017 ( .B1(n32738), .B2(n32739), .A(RST), .ZN(n1071) );
  OAI21_X1 U4018 ( .B1(n32740), .B2(n32739), .A(RST), .ZN(n1072) );
  OAI21_X1 U4019 ( .B1(n32745), .B2(n32741), .A(RST), .ZN(n1073) );
  OAI21_X1 U4020 ( .B1(n32745), .B2(n32742), .A(RST), .ZN(n1074) );
  OAI21_X1 U4021 ( .B1(n32745), .B2(n32743), .A(RST), .ZN(n1075) );
  OAI21_X1 U4022 ( .B1(n32745), .B2(n32744), .A(RST), .ZN(n1076) );
  NAND2_X1 U4023 ( .A1(EN), .A2(RD1), .ZN(n32746) );
  NAND2_X1 U4024 ( .A1(RST), .A2(n32746), .ZN(n5811) );
  NOR2_X1 U4025 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .ZN(n32747) );
  NAND2_X1 U4026 ( .A1(ADD_RD1[3]), .A2(n32747), .ZN(n32755) );
  INV_X1 U4027 ( .A(ADD_RD1[2]), .ZN(n32748) );
  INV_X1 U4028 ( .A(ADD_RD1[1]), .ZN(n32786) );
  NAND2_X1 U4029 ( .A1(n32748), .A2(n32786), .ZN(n32771) );
  NOR2_X1 U4030 ( .A1(n32755), .A2(n32771), .ZN(n33424) );
  NAND2_X1 U4031 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[1]), .ZN(n32763) );
  INV_X1 U4032 ( .A(ADD_RD1[3]), .ZN(n32749) );
  NAND3_X1 U4033 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[0]), .A3(n32749), .ZN(n32768)
         );
  NOR2_X1 U4034 ( .A1(n32763), .A2(n32768), .ZN(n33423) );
  AOI22_X1 U4035 ( .A1(n7424), .A2(n32685), .B1(n7416), .B2(n32684), .ZN(
        n32754) );
  NAND2_X1 U4036 ( .A1(ADD_RD1[2]), .A2(n32786), .ZN(n32770) );
  INV_X1 U4037 ( .A(ADD_RD1[4]), .ZN(n32762) );
  NAND3_X1 U4038 ( .A1(ADD_RD1[0]), .A2(n32762), .A3(n32749), .ZN(n32775) );
  NOR2_X1 U4039 ( .A1(n32770), .A2(n32775), .ZN(n33426) );
  NOR2_X1 U4040 ( .A1(n32771), .A2(n32775), .ZN(n33425) );
  AOI22_X1 U4041 ( .A1(n7430), .A2(n32687), .B1(n7420), .B2(n32686), .ZN(
        n32753) );
  INV_X1 U4042 ( .A(ADD_RD1[0]), .ZN(n32750) );
  NAND3_X1 U4043 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .A3(n32750), .ZN(n32760)
         );
  NOR2_X1 U4044 ( .A1(n32771), .A2(n32760), .ZN(n33428) );
  NAND2_X1 U4045 ( .A1(n32747), .A2(n32749), .ZN(n32769) );
  NOR2_X1 U4046 ( .A1(n32770), .A2(n32769), .ZN(n33427) );
  AOI22_X1 U4047 ( .A1(n7426), .A2(n32689), .B1(n7425), .B2(n32688), .ZN(
        n32752) );
  NAND2_X1 U4048 ( .A1(ADD_RD1[1]), .A2(n32748), .ZN(n32774) );
  NOR2_X1 U4049 ( .A1(n32755), .A2(n32774), .ZN(n33430) );
  NAND3_X1 U4050 ( .A1(ADD_RD1[4]), .A2(n32750), .A3(n32749), .ZN(n32773) );
  NOR2_X1 U4051 ( .A1(n32763), .A2(n32773), .ZN(n33429) );
  AOI22_X1 U4052 ( .A1(n7419), .A2(n32691), .B1(n7422), .B2(n32690), .ZN(
        n32751) );
  NAND4_X1 U4053 ( .A1(n32754), .A2(n32753), .A3(n32752), .A4(n32751), .ZN(
        n32783) );
  NOR2_X1 U4054 ( .A1(n32763), .A2(n32769), .ZN(n33436) );
  NOR2_X1 U4055 ( .A1(n32771), .A2(n32768), .ZN(n33435) );
  AOI22_X1 U4056 ( .A1(n7404), .A2(n32693), .B1(n7410), .B2(n32692), .ZN(
        n32759) );
  NOR2_X1 U4057 ( .A1(n32763), .A2(n32760), .ZN(n33438) );
  NOR2_X1 U4058 ( .A1(n32768), .A2(n32774), .ZN(n33437) );
  AOI22_X1 U4059 ( .A1(n7412), .A2(n32695), .B1(n7408), .B2(n32694), .ZN(
        n32758) );
  NOR2_X1 U4060 ( .A1(n32770), .A2(n32760), .ZN(n33440) );
  NOR2_X1 U4061 ( .A1(n32755), .A2(n32770), .ZN(n33439) );
  AOI22_X1 U4062 ( .A1(n7402), .A2(n32697), .B1(n7409), .B2(n32696), .ZN(
        n32757) );
  NAND3_X1 U4063 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(ADD_RD1[3]), .ZN(
        n32761) );
  NOR2_X1 U4064 ( .A1(n32770), .A2(n32761), .ZN(n33442) );
  NOR2_X1 U4065 ( .A1(n32755), .A2(n32763), .ZN(n33441) );
  AOI22_X1 U4066 ( .A1(n7414), .A2(n32699), .B1(n7406), .B2(n32698), .ZN(
        n32756) );
  NAND4_X1 U4067 ( .A1(n32759), .A2(n32758), .A3(n32757), .A4(n32756), .ZN(
        n32782) );
  NOR2_X1 U4068 ( .A1(n32771), .A2(n32761), .ZN(n33448) );
  NOR2_X1 U4069 ( .A1(n32763), .A2(n32775), .ZN(n33447) );
  AOI22_X1 U4070 ( .A1(n7411), .A2(n32701), .B1(n7428), .B2(n32700), .ZN(
        n32767) );
  NOR2_X1 U4071 ( .A1(n32769), .A2(n32774), .ZN(n33450) );
  NOR2_X1 U4072 ( .A1(n32760), .A2(n32774), .ZN(n33449) );
  AOI22_X1 U4073 ( .A1(n7418), .A2(n32703), .B1(n7415), .B2(n32702), .ZN(
        n32766) );
  NOR2_X1 U4074 ( .A1(n32770), .A2(n32773), .ZN(n33452) );
  NOR2_X1 U4075 ( .A1(n32774), .A2(n32761), .ZN(n33451) );
  AOI22_X1 U4076 ( .A1(n7401), .A2(n32705), .B1(n7427), .B2(n32704), .ZN(
        n32765) );
  NOR2_X1 U4077 ( .A1(n32763), .A2(n32761), .ZN(n33454) );
  NAND3_X1 U4078 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n32762), .ZN(n32772)
         );
  NOR2_X1 U4079 ( .A1(n32763), .A2(n32772), .ZN(n33453) );
  AOI22_X1 U4080 ( .A1(n7413), .A2(n32707), .B1(n7405), .B2(n32706), .ZN(
        n32764) );
  NAND4_X1 U4081 ( .A1(n32767), .A2(n32766), .A3(n32765), .A4(n32764), .ZN(
        n32781) );
  NOR2_X1 U4082 ( .A1(n32768), .A2(n32770), .ZN(n33460) );
  NOR2_X1 U4083 ( .A1(n32771), .A2(n32769), .ZN(n33459) );
  AOI22_X1 U4084 ( .A1(n7403), .A2(n32709), .B1(n7432), .B2(n32708), .ZN(
        n32779) );
  NOR2_X1 U4085 ( .A1(n32770), .A2(n32772), .ZN(n33462) );
  NOR2_X1 U4086 ( .A1(n32771), .A2(n32772), .ZN(n33461) );
  AOI22_X1 U4087 ( .A1(n7431), .A2(n32711), .B1(n7417), .B2(n32710), .ZN(
        n32778) );
  NOR2_X1 U4088 ( .A1(n32771), .A2(n32773), .ZN(n33464) );
  NOR2_X1 U4089 ( .A1(n32774), .A2(n32772), .ZN(n33463) );
  AOI22_X1 U4090 ( .A1(n7421), .A2(n32713), .B1(n7407), .B2(n32712), .ZN(
        n32777) );
  NOR2_X1 U4091 ( .A1(n32774), .A2(n32773), .ZN(n33466) );
  NOR2_X1 U4092 ( .A1(n32775), .A2(n32774), .ZN(n33465) );
  AOI22_X1 U4093 ( .A1(n7429), .A2(n32715), .B1(n7423), .B2(n32714), .ZN(
        n32776) );
  NAND4_X1 U4094 ( .A1(n32779), .A2(n32778), .A3(n32777), .A4(n32776), .ZN(
        n32780) );
  NOR4_X1 U4095 ( .A1(n32783), .A2(n32782), .A3(n32781), .A4(n32780), .ZN(
        n32792) );
  OAI22_X1 U4096 ( .A1(n33517), .A2(ADD_RD1[4]), .B1(n33516), .B2(ADD_RD1[3]), 
        .ZN(n32784) );
  AOI221_X1 U4097 ( .B1(n33517), .B2(ADD_RD1[4]), .C1(ADD_RD1[3]), .C2(n33516), 
        .A(n32784), .ZN(n32789) );
  OAI22_X1 U4098 ( .A1(n33520), .A2(ADD_RD1[0]), .B1(n33519), .B2(ADD_RD1[2]), 
        .ZN(n32785) );
  AOI221_X1 U4099 ( .B1(n33520), .B2(ADD_RD1[0]), .C1(ADD_RD1[2]), .C2(n33519), 
        .A(n32785), .ZN(n32788) );
  AOI22_X1 U4100 ( .A1(ADD_WR[1]), .A2(n32786), .B1(ADD_RD1[1]), .B2(n33521), 
        .ZN(n32787) );
  NAND4_X1 U4101 ( .A1(WR), .A2(n32789), .A3(n32788), .A4(n32787), .ZN(n32790)
         );
  NAND2_X1 U4102 ( .A1(RST), .A2(DATAIN[31]), .ZN(n34213) );
  INV_X1 U4103 ( .A(n32790), .ZN(n32791) );
  OAI22_X1 U4104 ( .A1(n32792), .A2(n33476), .B1(n34213), .B2(n33475), .ZN(
        n5777) );
  AOI22_X1 U4105 ( .A1(n32685), .A2(n7456), .B1(n32684), .B2(n7448), .ZN(
        n32796) );
  AOI22_X1 U4106 ( .A1(n32687), .A2(n7462), .B1(n32686), .B2(n7452), .ZN(
        n32795) );
  AOI22_X1 U4107 ( .A1(n32689), .A2(n7458), .B1(n32688), .B2(n7457), .ZN(
        n32794) );
  AOI22_X1 U4108 ( .A1(n32691), .A2(n7451), .B1(n32690), .B2(n7454), .ZN(
        n32793) );
  NAND4_X1 U4109 ( .A1(n32796), .A2(n32795), .A3(n32794), .A4(n32793), .ZN(
        n32812) );
  AOI22_X1 U4110 ( .A1(n32693), .A2(n7436), .B1(n32692), .B2(n7442), .ZN(
        n32800) );
  AOI22_X1 U4111 ( .A1(n32695), .A2(n7444), .B1(n32694), .B2(n7440), .ZN(
        n32799) );
  AOI22_X1 U4112 ( .A1(n32697), .A2(n7434), .B1(n32696), .B2(n7441), .ZN(
        n32798) );
  AOI22_X1 U4113 ( .A1(n32699), .A2(n7446), .B1(n32698), .B2(n7438), .ZN(
        n32797) );
  NAND4_X1 U4114 ( .A1(n32800), .A2(n32799), .A3(n32798), .A4(n32797), .ZN(
        n32811) );
  AOI22_X1 U4115 ( .A1(n32701), .A2(n7443), .B1(n32700), .B2(n7460), .ZN(
        n32804) );
  AOI22_X1 U4116 ( .A1(n32703), .A2(n7450), .B1(n32702), .B2(n7447), .ZN(
        n32803) );
  AOI22_X1 U4117 ( .A1(n32705), .A2(n7433), .B1(n32704), .B2(n7459), .ZN(
        n32802) );
  AOI22_X1 U4118 ( .A1(n32707), .A2(n7445), .B1(n32706), .B2(n7437), .ZN(
        n32801) );
  NAND4_X1 U4119 ( .A1(n32804), .A2(n32803), .A3(n32802), .A4(n32801), .ZN(
        n32810) );
  AOI22_X1 U4120 ( .A1(n32709), .A2(n7435), .B1(n32708), .B2(n7464), .ZN(
        n32808) );
  AOI22_X1 U4121 ( .A1(n32711), .A2(n7463), .B1(n32710), .B2(n7449), .ZN(
        n32807) );
  AOI22_X1 U4122 ( .A1(n32713), .A2(n7453), .B1(n32712), .B2(n7439), .ZN(
        n32806) );
  AOI22_X1 U4123 ( .A1(n32715), .A2(n7461), .B1(n32714), .B2(n7455), .ZN(
        n32805) );
  NAND4_X1 U4124 ( .A1(n32808), .A2(n32807), .A3(n32806), .A4(n32805), .ZN(
        n32809) );
  NOR4_X1 U4125 ( .A1(n32812), .A2(n32811), .A3(n32810), .A4(n32809), .ZN(
        n32813) );
  NAND2_X1 U4126 ( .A1(RST), .A2(DATAIN[30]), .ZN(n34214) );
  OAI22_X1 U4127 ( .A1(n32813), .A2(n33476), .B1(n33475), .B2(n34214), .ZN(
        n5778) );
  AOI22_X1 U4128 ( .A1(n32685), .A2(n7488), .B1(n32684), .B2(n7480), .ZN(
        n32817) );
  AOI22_X1 U4129 ( .A1(n32687), .A2(n7494), .B1(n32686), .B2(n7484), .ZN(
        n32816) );
  AOI22_X1 U4130 ( .A1(n32689), .A2(n7490), .B1(n32688), .B2(n7489), .ZN(
        n32815) );
  AOI22_X1 U4131 ( .A1(n32691), .A2(n7483), .B1(n32690), .B2(n7486), .ZN(
        n32814) );
  NAND4_X1 U4132 ( .A1(n32817), .A2(n32816), .A3(n32815), .A4(n32814), .ZN(
        n32833) );
  AOI22_X1 U4133 ( .A1(n32693), .A2(n7468), .B1(n32692), .B2(n7474), .ZN(
        n32821) );
  AOI22_X1 U4134 ( .A1(n32695), .A2(n7476), .B1(n32694), .B2(n7472), .ZN(
        n32820) );
  AOI22_X1 U4135 ( .A1(n32697), .A2(n7466), .B1(n32696), .B2(n7473), .ZN(
        n32819) );
  AOI22_X1 U4136 ( .A1(n32699), .A2(n7478), .B1(n32698), .B2(n7470), .ZN(
        n32818) );
  NAND4_X1 U4137 ( .A1(n32821), .A2(n32820), .A3(n32819), .A4(n32818), .ZN(
        n32832) );
  AOI22_X1 U4138 ( .A1(n32701), .A2(n7475), .B1(n32700), .B2(n7492), .ZN(
        n32825) );
  AOI22_X1 U4139 ( .A1(n32703), .A2(n7482), .B1(n32702), .B2(n7479), .ZN(
        n32824) );
  AOI22_X1 U4140 ( .A1(n32705), .A2(n7465), .B1(n32704), .B2(n7491), .ZN(
        n32823) );
  AOI22_X1 U4141 ( .A1(n32707), .A2(n7477), .B1(n32706), .B2(n7469), .ZN(
        n32822) );
  NAND4_X1 U4142 ( .A1(n32825), .A2(n32824), .A3(n32823), .A4(n32822), .ZN(
        n32831) );
  AOI22_X1 U4143 ( .A1(n32709), .A2(n7467), .B1(n32708), .B2(n7496), .ZN(
        n32829) );
  AOI22_X1 U4144 ( .A1(n32711), .A2(n7495), .B1(n32710), .B2(n7481), .ZN(
        n32828) );
  AOI22_X1 U4145 ( .A1(n32713), .A2(n7485), .B1(n32712), .B2(n7471), .ZN(
        n32827) );
  AOI22_X1 U4146 ( .A1(n32715), .A2(n7493), .B1(n32714), .B2(n7487), .ZN(
        n32826) );
  NAND4_X1 U4147 ( .A1(n32829), .A2(n32828), .A3(n32827), .A4(n32826), .ZN(
        n32830) );
  NOR4_X1 U4148 ( .A1(n32833), .A2(n32832), .A3(n32831), .A4(n32830), .ZN(
        n32834) );
  NAND2_X1 U4149 ( .A1(RST), .A2(DATAIN[29]), .ZN(n34215) );
  OAI22_X1 U4150 ( .A1(n32834), .A2(n33476), .B1(n33475), .B2(n34215), .ZN(
        n5779) );
  AOI22_X1 U4151 ( .A1(n32685), .A2(n7520), .B1(n32684), .B2(n7512), .ZN(
        n32838) );
  AOI22_X1 U4152 ( .A1(n32687), .A2(n7526), .B1(n32686), .B2(n7516), .ZN(
        n32837) );
  AOI22_X1 U4153 ( .A1(n32689), .A2(n7522), .B1(n32688), .B2(n7521), .ZN(
        n32836) );
  AOI22_X1 U4154 ( .A1(n32691), .A2(n7515), .B1(n32690), .B2(n7518), .ZN(
        n32835) );
  NAND4_X1 U4155 ( .A1(n32838), .A2(n32837), .A3(n32836), .A4(n32835), .ZN(
        n32854) );
  AOI22_X1 U4156 ( .A1(n32693), .A2(n7500), .B1(n32692), .B2(n7506), .ZN(
        n32842) );
  AOI22_X1 U4157 ( .A1(n32695), .A2(n7508), .B1(n32694), .B2(n7504), .ZN(
        n32841) );
  AOI22_X1 U4158 ( .A1(n32697), .A2(n7498), .B1(n32696), .B2(n7505), .ZN(
        n32840) );
  AOI22_X1 U4159 ( .A1(n32699), .A2(n7510), .B1(n32698), .B2(n7502), .ZN(
        n32839) );
  NAND4_X1 U4160 ( .A1(n32842), .A2(n32841), .A3(n32840), .A4(n32839), .ZN(
        n32853) );
  AOI22_X1 U4161 ( .A1(n32701), .A2(n7507), .B1(n32700), .B2(n7524), .ZN(
        n32846) );
  AOI22_X1 U4162 ( .A1(n32703), .A2(n7514), .B1(n32702), .B2(n7511), .ZN(
        n32845) );
  AOI22_X1 U4163 ( .A1(n32705), .A2(n7497), .B1(n32704), .B2(n7523), .ZN(
        n32844) );
  AOI22_X1 U4164 ( .A1(n32707), .A2(n7509), .B1(n32706), .B2(n7501), .ZN(
        n32843) );
  NAND4_X1 U4165 ( .A1(n32846), .A2(n32845), .A3(n32844), .A4(n32843), .ZN(
        n32852) );
  AOI22_X1 U4166 ( .A1(n32709), .A2(n7499), .B1(n32708), .B2(n7528), .ZN(
        n32850) );
  AOI22_X1 U4167 ( .A1(n32711), .A2(n7527), .B1(n32710), .B2(n7513), .ZN(
        n32849) );
  AOI22_X1 U4168 ( .A1(n32713), .A2(n7517), .B1(n32712), .B2(n7503), .ZN(
        n32848) );
  AOI22_X1 U4169 ( .A1(n32715), .A2(n7525), .B1(n32714), .B2(n7519), .ZN(
        n32847) );
  NAND4_X1 U4170 ( .A1(n32850), .A2(n32849), .A3(n32848), .A4(n32847), .ZN(
        n32851) );
  NOR4_X1 U4171 ( .A1(n32854), .A2(n32853), .A3(n32852), .A4(n32851), .ZN(
        n32855) );
  NAND2_X1 U4172 ( .A1(RST), .A2(DATAIN[28]), .ZN(n34216) );
  OAI22_X1 U4173 ( .A1(n32855), .A2(n33476), .B1(n33475), .B2(n34216), .ZN(
        n5780) );
  AOI22_X1 U4174 ( .A1(n32685), .A2(n7552), .B1(n32684), .B2(n7544), .ZN(
        n32859) );
  AOI22_X1 U4175 ( .A1(n32687), .A2(n7558), .B1(n32686), .B2(n7548), .ZN(
        n32858) );
  AOI22_X1 U4176 ( .A1(n32689), .A2(n7554), .B1(n32688), .B2(n7553), .ZN(
        n32857) );
  AOI22_X1 U4177 ( .A1(n32691), .A2(n7547), .B1(n32690), .B2(n7550), .ZN(
        n32856) );
  NAND4_X1 U4178 ( .A1(n32859), .A2(n32858), .A3(n32857), .A4(n32856), .ZN(
        n32875) );
  AOI22_X1 U4179 ( .A1(n32693), .A2(n7532), .B1(n32692), .B2(n7538), .ZN(
        n32863) );
  AOI22_X1 U4180 ( .A1(n32695), .A2(n7540), .B1(n32694), .B2(n7536), .ZN(
        n32862) );
  AOI22_X1 U4181 ( .A1(n32697), .A2(n7530), .B1(n32696), .B2(n7537), .ZN(
        n32861) );
  AOI22_X1 U4182 ( .A1(n32699), .A2(n7542), .B1(n32698), .B2(n7534), .ZN(
        n32860) );
  NAND4_X1 U4183 ( .A1(n32863), .A2(n32862), .A3(n32861), .A4(n32860), .ZN(
        n32874) );
  AOI22_X1 U4184 ( .A1(n32701), .A2(n7539), .B1(n32700), .B2(n7556), .ZN(
        n32867) );
  AOI22_X1 U4185 ( .A1(n32703), .A2(n7546), .B1(n32702), .B2(n7543), .ZN(
        n32866) );
  AOI22_X1 U4186 ( .A1(n32705), .A2(n7529), .B1(n32704), .B2(n7555), .ZN(
        n32865) );
  AOI22_X1 U4187 ( .A1(n32707), .A2(n7541), .B1(n32706), .B2(n7533), .ZN(
        n32864) );
  NAND4_X1 U4188 ( .A1(n32867), .A2(n32866), .A3(n32865), .A4(n32864), .ZN(
        n32873) );
  AOI22_X1 U4189 ( .A1(n32709), .A2(n7531), .B1(n32708), .B2(n7560), .ZN(
        n32871) );
  AOI22_X1 U4190 ( .A1(n32711), .A2(n7559), .B1(n32710), .B2(n7545), .ZN(
        n32870) );
  AOI22_X1 U4191 ( .A1(n32713), .A2(n7549), .B1(n32712), .B2(n7535), .ZN(
        n32869) );
  AOI22_X1 U4192 ( .A1(n32715), .A2(n7557), .B1(n32714), .B2(n7551), .ZN(
        n32868) );
  NAND4_X1 U4193 ( .A1(n32871), .A2(n32870), .A3(n32869), .A4(n32868), .ZN(
        n32872) );
  NOR4_X1 U4194 ( .A1(n32875), .A2(n32874), .A3(n32873), .A4(n32872), .ZN(
        n32876) );
  OAI22_X1 U4195 ( .A1(n32876), .A2(n33476), .B1(n33475), .B2(n32723), .ZN(
        n5781) );
  AOI22_X1 U4196 ( .A1(n32685), .A2(n7584), .B1(n32684), .B2(n7576), .ZN(
        n32880) );
  AOI22_X1 U4197 ( .A1(n32687), .A2(n7590), .B1(n32686), .B2(n7580), .ZN(
        n32879) );
  AOI22_X1 U4198 ( .A1(n32689), .A2(n7586), .B1(n32688), .B2(n7585), .ZN(
        n32878) );
  AOI22_X1 U4199 ( .A1(n32691), .A2(n7579), .B1(n32690), .B2(n7582), .ZN(
        n32877) );
  NAND4_X1 U4200 ( .A1(n32880), .A2(n32879), .A3(n32878), .A4(n32877), .ZN(
        n32896) );
  AOI22_X1 U4201 ( .A1(n32693), .A2(n7564), .B1(n32692), .B2(n7570), .ZN(
        n32884) );
  AOI22_X1 U4202 ( .A1(n32695), .A2(n7572), .B1(n32694), .B2(n7568), .ZN(
        n32883) );
  AOI22_X1 U4203 ( .A1(n32697), .A2(n7562), .B1(n32696), .B2(n7569), .ZN(
        n32882) );
  AOI22_X1 U4204 ( .A1(n32699), .A2(n7574), .B1(n32698), .B2(n7566), .ZN(
        n32881) );
  NAND4_X1 U4205 ( .A1(n32884), .A2(n32883), .A3(n32882), .A4(n32881), .ZN(
        n32895) );
  AOI22_X1 U4206 ( .A1(n32701), .A2(n7571), .B1(n32700), .B2(n7588), .ZN(
        n32888) );
  AOI22_X1 U4207 ( .A1(n32703), .A2(n7578), .B1(n32702), .B2(n7575), .ZN(
        n32887) );
  AOI22_X1 U4208 ( .A1(n32705), .A2(n7561), .B1(n32704), .B2(n7587), .ZN(
        n32886) );
  AOI22_X1 U4209 ( .A1(n32707), .A2(n7573), .B1(n32706), .B2(n7565), .ZN(
        n32885) );
  NAND4_X1 U4210 ( .A1(n32888), .A2(n32887), .A3(n32886), .A4(n32885), .ZN(
        n32894) );
  AOI22_X1 U4211 ( .A1(n32709), .A2(n7563), .B1(n32708), .B2(n7592), .ZN(
        n32892) );
  AOI22_X1 U4212 ( .A1(n32711), .A2(n7591), .B1(n32710), .B2(n7577), .ZN(
        n32891) );
  AOI22_X1 U4213 ( .A1(n32713), .A2(n7581), .B1(n32712), .B2(n7567), .ZN(
        n32890) );
  AOI22_X1 U4214 ( .A1(n32715), .A2(n7589), .B1(n32714), .B2(n7583), .ZN(
        n32889) );
  NAND4_X1 U4215 ( .A1(n32892), .A2(n32891), .A3(n32890), .A4(n32889), .ZN(
        n32893) );
  NOR4_X1 U4216 ( .A1(n32896), .A2(n32895), .A3(n32894), .A4(n32893), .ZN(
        n32897) );
  OAI22_X1 U4217 ( .A1(n32897), .A2(n33476), .B1(n33475), .B2(n20327), .ZN(
        n5782) );
  AOI22_X1 U4218 ( .A1(n32685), .A2(n7616), .B1(n32684), .B2(n7608), .ZN(
        n32901) );
  AOI22_X1 U4219 ( .A1(n32687), .A2(n7622), .B1(n32686), .B2(n7612), .ZN(
        n32900) );
  AOI22_X1 U4220 ( .A1(n32689), .A2(n7618), .B1(n32688), .B2(n7617), .ZN(
        n32899) );
  AOI22_X1 U4221 ( .A1(n32691), .A2(n7611), .B1(n32690), .B2(n7614), .ZN(
        n32898) );
  NAND4_X1 U4222 ( .A1(n32901), .A2(n32900), .A3(n32899), .A4(n32898), .ZN(
        n32917) );
  AOI22_X1 U4223 ( .A1(n32693), .A2(n7596), .B1(n32692), .B2(n7602), .ZN(
        n32905) );
  AOI22_X1 U4224 ( .A1(n32695), .A2(n7604), .B1(n32694), .B2(n7600), .ZN(
        n32904) );
  AOI22_X1 U4225 ( .A1(n32697), .A2(n7594), .B1(n32696), .B2(n7601), .ZN(
        n32903) );
  AOI22_X1 U4226 ( .A1(n32699), .A2(n7606), .B1(n32698), .B2(n7598), .ZN(
        n32902) );
  NAND4_X1 U4227 ( .A1(n32905), .A2(n32904), .A3(n32903), .A4(n32902), .ZN(
        n32916) );
  AOI22_X1 U4228 ( .A1(n32701), .A2(n7603), .B1(n32700), .B2(n7620), .ZN(
        n32909) );
  AOI22_X1 U4229 ( .A1(n32703), .A2(n7610), .B1(n32702), .B2(n7607), .ZN(
        n32908) );
  AOI22_X1 U4230 ( .A1(n32705), .A2(n7593), .B1(n32704), .B2(n7619), .ZN(
        n32907) );
  AOI22_X1 U4231 ( .A1(n32707), .A2(n7605), .B1(n32706), .B2(n7597), .ZN(
        n32906) );
  NAND4_X1 U4232 ( .A1(n32909), .A2(n32908), .A3(n32907), .A4(n32906), .ZN(
        n32915) );
  AOI22_X1 U4233 ( .A1(n32709), .A2(n7595), .B1(n32708), .B2(n7624), .ZN(
        n32913) );
  AOI22_X1 U4234 ( .A1(n32711), .A2(n7623), .B1(n32710), .B2(n7609), .ZN(
        n32912) );
  AOI22_X1 U4235 ( .A1(n32713), .A2(n7613), .B1(n32712), .B2(n7599), .ZN(
        n32911) );
  AOI22_X1 U4236 ( .A1(n32715), .A2(n7621), .B1(n32714), .B2(n7615), .ZN(
        n32910) );
  NAND4_X1 U4237 ( .A1(n32913), .A2(n32912), .A3(n32911), .A4(n32910), .ZN(
        n32914) );
  NOR4_X1 U4238 ( .A1(n32917), .A2(n32916), .A3(n32915), .A4(n32914), .ZN(
        n32918) );
  OAI22_X1 U4239 ( .A1(n32918), .A2(n33476), .B1(n33475), .B2(n14130), .ZN(
        n5783) );
  AOI22_X1 U4240 ( .A1(n32685), .A2(n7648), .B1(n32684), .B2(n7640), .ZN(
        n32922) );
  AOI22_X1 U4241 ( .A1(n32687), .A2(n7654), .B1(n32686), .B2(n7644), .ZN(
        n32921) );
  AOI22_X1 U4242 ( .A1(n32689), .A2(n7650), .B1(n32688), .B2(n7649), .ZN(
        n32920) );
  AOI22_X1 U4243 ( .A1(n32691), .A2(n7643), .B1(n32690), .B2(n7646), .ZN(
        n32919) );
  NAND4_X1 U4244 ( .A1(n32922), .A2(n32921), .A3(n32920), .A4(n32919), .ZN(
        n32938) );
  AOI22_X1 U4245 ( .A1(n32693), .A2(n7628), .B1(n32692), .B2(n7634), .ZN(
        n32926) );
  AOI22_X1 U4246 ( .A1(n32695), .A2(n7636), .B1(n32694), .B2(n7632), .ZN(
        n32925) );
  AOI22_X1 U4247 ( .A1(n32697), .A2(n7626), .B1(n32696), .B2(n7633), .ZN(
        n32924) );
  AOI22_X1 U4248 ( .A1(n32699), .A2(n7638), .B1(n32698), .B2(n7630), .ZN(
        n32923) );
  NAND4_X1 U4249 ( .A1(n32926), .A2(n32925), .A3(n32924), .A4(n32923), .ZN(
        n32937) );
  AOI22_X1 U4250 ( .A1(n32701), .A2(n7635), .B1(n32700), .B2(n7652), .ZN(
        n32930) );
  AOI22_X1 U4251 ( .A1(n32703), .A2(n7642), .B1(n32702), .B2(n7639), .ZN(
        n32929) );
  AOI22_X1 U4252 ( .A1(n32705), .A2(n7625), .B1(n32704), .B2(n7651), .ZN(
        n32928) );
  AOI22_X1 U4253 ( .A1(n32707), .A2(n7637), .B1(n32706), .B2(n7629), .ZN(
        n32927) );
  NAND4_X1 U4254 ( .A1(n32930), .A2(n32929), .A3(n32928), .A4(n32927), .ZN(
        n32936) );
  AOI22_X1 U4255 ( .A1(n32709), .A2(n7627), .B1(n32708), .B2(n7656), .ZN(
        n32934) );
  AOI22_X1 U4256 ( .A1(n32711), .A2(n7655), .B1(n32710), .B2(n7641), .ZN(
        n32933) );
  AOI22_X1 U4257 ( .A1(n32713), .A2(n7645), .B1(n32712), .B2(n7631), .ZN(
        n32932) );
  AOI22_X1 U4258 ( .A1(n32715), .A2(n7653), .B1(n32714), .B2(n7647), .ZN(
        n32931) );
  NAND4_X1 U4259 ( .A1(n32934), .A2(n32933), .A3(n32932), .A4(n32931), .ZN(
        n32935) );
  NOR4_X1 U4260 ( .A1(n32938), .A2(n32937), .A3(n32936), .A4(n32935), .ZN(
        n32939) );
  OAI22_X1 U4261 ( .A1(n32939), .A2(n33476), .B1(n33475), .B2(n14131), .ZN(
        n5784) );
  AOI22_X1 U4262 ( .A1(n32685), .A2(n7680), .B1(n32684), .B2(n7672), .ZN(
        n32943) );
  AOI22_X1 U4263 ( .A1(n32687), .A2(n7686), .B1(n32686), .B2(n7676), .ZN(
        n32942) );
  AOI22_X1 U4264 ( .A1(n32689), .A2(n7682), .B1(n32688), .B2(n7681), .ZN(
        n32941) );
  AOI22_X1 U4265 ( .A1(n32691), .A2(n7675), .B1(n32690), .B2(n7678), .ZN(
        n32940) );
  NAND4_X1 U4266 ( .A1(n32943), .A2(n32942), .A3(n32941), .A4(n32940), .ZN(
        n32959) );
  AOI22_X1 U4267 ( .A1(n32693), .A2(n7660), .B1(n32692), .B2(n7666), .ZN(
        n32947) );
  AOI22_X1 U4268 ( .A1(n32695), .A2(n7668), .B1(n32694), .B2(n7664), .ZN(
        n32946) );
  AOI22_X1 U4269 ( .A1(n32697), .A2(n7658), .B1(n32696), .B2(n7665), .ZN(
        n32945) );
  AOI22_X1 U4270 ( .A1(n32699), .A2(n7670), .B1(n32698), .B2(n7662), .ZN(
        n32944) );
  NAND4_X1 U4271 ( .A1(n32947), .A2(n32946), .A3(n32945), .A4(n32944), .ZN(
        n32958) );
  AOI22_X1 U4272 ( .A1(n32701), .A2(n7667), .B1(n32700), .B2(n7684), .ZN(
        n32951) );
  AOI22_X1 U4273 ( .A1(n32703), .A2(n7674), .B1(n32702), .B2(n7671), .ZN(
        n32950) );
  AOI22_X1 U4274 ( .A1(n32705), .A2(n7657), .B1(n32704), .B2(n7683), .ZN(
        n32949) );
  AOI22_X1 U4275 ( .A1(n32707), .A2(n7669), .B1(n32706), .B2(n7661), .ZN(
        n32948) );
  NAND4_X1 U4276 ( .A1(n32951), .A2(n32950), .A3(n32949), .A4(n32948), .ZN(
        n32957) );
  AOI22_X1 U4277 ( .A1(n32709), .A2(n7659), .B1(n32708), .B2(n7688), .ZN(
        n32955) );
  AOI22_X1 U4278 ( .A1(n32711), .A2(n7687), .B1(n32710), .B2(n7673), .ZN(
        n32954) );
  AOI22_X1 U4279 ( .A1(n32713), .A2(n7677), .B1(n32712), .B2(n7663), .ZN(
        n32953) );
  AOI22_X1 U4280 ( .A1(n32715), .A2(n7685), .B1(n32714), .B2(n7679), .ZN(
        n32952) );
  NAND4_X1 U4281 ( .A1(n32955), .A2(n32954), .A3(n32953), .A4(n32952), .ZN(
        n32956) );
  NOR4_X1 U4282 ( .A1(n32959), .A2(n32958), .A3(n32957), .A4(n32956), .ZN(
        n32960) );
  OAI22_X1 U4283 ( .A1(n32960), .A2(n33476), .B1(n33475), .B2(n14132), .ZN(
        n5785) );
  AOI22_X1 U4284 ( .A1(n32685), .A2(n7712), .B1(n32684), .B2(n7704), .ZN(
        n32964) );
  AOI22_X1 U4285 ( .A1(n32687), .A2(n7718), .B1(n32686), .B2(n7708), .ZN(
        n32963) );
  AOI22_X1 U4286 ( .A1(n32689), .A2(n7714), .B1(n32688), .B2(n7713), .ZN(
        n32962) );
  AOI22_X1 U4287 ( .A1(n32691), .A2(n7707), .B1(n32690), .B2(n7710), .ZN(
        n32961) );
  NAND4_X1 U4288 ( .A1(n32964), .A2(n32963), .A3(n32962), .A4(n32961), .ZN(
        n32980) );
  AOI22_X1 U4289 ( .A1(n32693), .A2(n7692), .B1(n32692), .B2(n7698), .ZN(
        n32968) );
  AOI22_X1 U4290 ( .A1(n32695), .A2(n7700), .B1(n32694), .B2(n7696), .ZN(
        n32967) );
  AOI22_X1 U4291 ( .A1(n32697), .A2(n7690), .B1(n32696), .B2(n7697), .ZN(
        n32966) );
  AOI22_X1 U4292 ( .A1(n32699), .A2(n7702), .B1(n32698), .B2(n7694), .ZN(
        n32965) );
  NAND4_X1 U4293 ( .A1(n32968), .A2(n32967), .A3(n32966), .A4(n32965), .ZN(
        n32979) );
  AOI22_X1 U4294 ( .A1(n32701), .A2(n7699), .B1(n32700), .B2(n7716), .ZN(
        n32972) );
  AOI22_X1 U4295 ( .A1(n32703), .A2(n7706), .B1(n32702), .B2(n7703), .ZN(
        n32971) );
  AOI22_X1 U4296 ( .A1(n32705), .A2(n7689), .B1(n32704), .B2(n7715), .ZN(
        n32970) );
  AOI22_X1 U4297 ( .A1(n32707), .A2(n7701), .B1(n32706), .B2(n7693), .ZN(
        n32969) );
  NAND4_X1 U4298 ( .A1(n32972), .A2(n32971), .A3(n32970), .A4(n32969), .ZN(
        n32978) );
  AOI22_X1 U4299 ( .A1(n32709), .A2(n7691), .B1(n32708), .B2(n7720), .ZN(
        n32976) );
  AOI22_X1 U4300 ( .A1(n32711), .A2(n7719), .B1(n32710), .B2(n7705), .ZN(
        n32975) );
  AOI22_X1 U4301 ( .A1(n32713), .A2(n7709), .B1(n32712), .B2(n7695), .ZN(
        n32974) );
  AOI22_X1 U4302 ( .A1(n32715), .A2(n7717), .B1(n32714), .B2(n7711), .ZN(
        n32973) );
  NAND4_X1 U4303 ( .A1(n32976), .A2(n32975), .A3(n32974), .A4(n32973), .ZN(
        n32977) );
  NOR4_X1 U4304 ( .A1(n32980), .A2(n32979), .A3(n32978), .A4(n32977), .ZN(
        n32981) );
  OAI22_X1 U4305 ( .A1(n32981), .A2(n33476), .B1(n33475), .B2(n32730), .ZN(
        n5786) );
  AOI22_X1 U4306 ( .A1(n32685), .A2(n7744), .B1(n32684), .B2(n7736), .ZN(
        n32985) );
  AOI22_X1 U4307 ( .A1(n32687), .A2(n7750), .B1(n32686), .B2(n7740), .ZN(
        n32984) );
  AOI22_X1 U4308 ( .A1(n32689), .A2(n7746), .B1(n32688), .B2(n7745), .ZN(
        n32983) );
  AOI22_X1 U4309 ( .A1(n32691), .A2(n7739), .B1(n32690), .B2(n7742), .ZN(
        n32982) );
  NAND4_X1 U4310 ( .A1(n32985), .A2(n32984), .A3(n32983), .A4(n32982), .ZN(
        n33001) );
  AOI22_X1 U4311 ( .A1(n32693), .A2(n7724), .B1(n32692), .B2(n7730), .ZN(
        n32989) );
  AOI22_X1 U4312 ( .A1(n32695), .A2(n7732), .B1(n32694), .B2(n7728), .ZN(
        n32988) );
  AOI22_X1 U4313 ( .A1(n32697), .A2(n7722), .B1(n32696), .B2(n7729), .ZN(
        n32987) );
  AOI22_X1 U4314 ( .A1(n32699), .A2(n7734), .B1(n32698), .B2(n7726), .ZN(
        n32986) );
  NAND4_X1 U4315 ( .A1(n32989), .A2(n32988), .A3(n32987), .A4(n32986), .ZN(
        n33000) );
  AOI22_X1 U4316 ( .A1(n32701), .A2(n7731), .B1(n32700), .B2(n7748), .ZN(
        n32993) );
  AOI22_X1 U4317 ( .A1(n32703), .A2(n7738), .B1(n32702), .B2(n7735), .ZN(
        n32992) );
  AOI22_X1 U4318 ( .A1(n32705), .A2(n7721), .B1(n32704), .B2(n7747), .ZN(
        n32991) );
  AOI22_X1 U4319 ( .A1(n32707), .A2(n7733), .B1(n32706), .B2(n7725), .ZN(
        n32990) );
  NAND4_X1 U4320 ( .A1(n32993), .A2(n32992), .A3(n32991), .A4(n32990), .ZN(
        n32999) );
  AOI22_X1 U4321 ( .A1(n32709), .A2(n7723), .B1(n32708), .B2(n7752), .ZN(
        n32997) );
  AOI22_X1 U4322 ( .A1(n32711), .A2(n7751), .B1(n32710), .B2(n7737), .ZN(
        n32996) );
  AOI22_X1 U4323 ( .A1(n32713), .A2(n7741), .B1(n32712), .B2(n7727), .ZN(
        n32995) );
  AOI22_X1 U4324 ( .A1(n32715), .A2(n7749), .B1(n32714), .B2(n7743), .ZN(
        n32994) );
  NAND4_X1 U4325 ( .A1(n32997), .A2(n32996), .A3(n32995), .A4(n32994), .ZN(
        n32998) );
  NOR4_X1 U4326 ( .A1(n33001), .A2(n33000), .A3(n32999), .A4(n32998), .ZN(
        n33002) );
  OAI22_X1 U4327 ( .A1(n33002), .A2(n33476), .B1(n33475), .B2(n14134), .ZN(
        n5787) );
  AOI22_X1 U4328 ( .A1(n32685), .A2(n7776), .B1(n32684), .B2(n7768), .ZN(
        n33006) );
  AOI22_X1 U4329 ( .A1(n32687), .A2(n7782), .B1(n32686), .B2(n7772), .ZN(
        n33005) );
  AOI22_X1 U4330 ( .A1(n32689), .A2(n7778), .B1(n32688), .B2(n7777), .ZN(
        n33004) );
  AOI22_X1 U4331 ( .A1(n32691), .A2(n7771), .B1(n32690), .B2(n7774), .ZN(
        n33003) );
  NAND4_X1 U4332 ( .A1(n33006), .A2(n33005), .A3(n33004), .A4(n33003), .ZN(
        n33022) );
  AOI22_X1 U4333 ( .A1(n32693), .A2(n7756), .B1(n32692), .B2(n7762), .ZN(
        n33010) );
  AOI22_X1 U4334 ( .A1(n32695), .A2(n7764), .B1(n32694), .B2(n7760), .ZN(
        n33009) );
  AOI22_X1 U4335 ( .A1(n32697), .A2(n7754), .B1(n32696), .B2(n7761), .ZN(
        n33008) );
  AOI22_X1 U4336 ( .A1(n32699), .A2(n7766), .B1(n32698), .B2(n7758), .ZN(
        n33007) );
  NAND4_X1 U4337 ( .A1(n33010), .A2(n33009), .A3(n33008), .A4(n33007), .ZN(
        n33021) );
  AOI22_X1 U4338 ( .A1(n32701), .A2(n7763), .B1(n32700), .B2(n7780), .ZN(
        n33014) );
  AOI22_X1 U4339 ( .A1(n32703), .A2(n7770), .B1(n32702), .B2(n7767), .ZN(
        n33013) );
  AOI22_X1 U4340 ( .A1(n32705), .A2(n7753), .B1(n32704), .B2(n7779), .ZN(
        n33012) );
  AOI22_X1 U4341 ( .A1(n32707), .A2(n7765), .B1(n32706), .B2(n7757), .ZN(
        n33011) );
  NAND4_X1 U4342 ( .A1(n33014), .A2(n33013), .A3(n33012), .A4(n33011), .ZN(
        n33020) );
  AOI22_X1 U4343 ( .A1(n32709), .A2(n7755), .B1(n32708), .B2(n7784), .ZN(
        n33018) );
  AOI22_X1 U4344 ( .A1(n32711), .A2(n7783), .B1(n32710), .B2(n7769), .ZN(
        n33017) );
  AOI22_X1 U4345 ( .A1(n32713), .A2(n7773), .B1(n32712), .B2(n7759), .ZN(
        n33016) );
  AOI22_X1 U4346 ( .A1(n32715), .A2(n7781), .B1(n32714), .B2(n7775), .ZN(
        n33015) );
  NAND4_X1 U4347 ( .A1(n33018), .A2(n33017), .A3(n33016), .A4(n33015), .ZN(
        n33019) );
  NOR4_X1 U4348 ( .A1(n33022), .A2(n33021), .A3(n33020), .A4(n33019), .ZN(
        n33023) );
  OAI22_X1 U4349 ( .A1(n33023), .A2(n33476), .B1(n33475), .B2(n14135), .ZN(
        n5788) );
  AOI22_X1 U4350 ( .A1(n32685), .A2(n7808), .B1(n32684), .B2(n7800), .ZN(
        n33027) );
  AOI22_X1 U4351 ( .A1(n32687), .A2(n7814), .B1(n32686), .B2(n7804), .ZN(
        n33026) );
  AOI22_X1 U4352 ( .A1(n32689), .A2(n7810), .B1(n32688), .B2(n7809), .ZN(
        n33025) );
  AOI22_X1 U4353 ( .A1(n32691), .A2(n7803), .B1(n32690), .B2(n7806), .ZN(
        n33024) );
  NAND4_X1 U4354 ( .A1(n33027), .A2(n33026), .A3(n33025), .A4(n33024), .ZN(
        n33043) );
  AOI22_X1 U4355 ( .A1(n32693), .A2(n7788), .B1(n32692), .B2(n7794), .ZN(
        n33031) );
  AOI22_X1 U4356 ( .A1(n32695), .A2(n7796), .B1(n32694), .B2(n7792), .ZN(
        n33030) );
  AOI22_X1 U4357 ( .A1(n32697), .A2(n7786), .B1(n32696), .B2(n7793), .ZN(
        n33029) );
  AOI22_X1 U4358 ( .A1(n32699), .A2(n7798), .B1(n32698), .B2(n7790), .ZN(
        n33028) );
  NAND4_X1 U4359 ( .A1(n33031), .A2(n33030), .A3(n33029), .A4(n33028), .ZN(
        n33042) );
  AOI22_X1 U4360 ( .A1(n32701), .A2(n7795), .B1(n32700), .B2(n7812), .ZN(
        n33035) );
  AOI22_X1 U4361 ( .A1(n32703), .A2(n7802), .B1(n32702), .B2(n7799), .ZN(
        n33034) );
  AOI22_X1 U4362 ( .A1(n32705), .A2(n7785), .B1(n32704), .B2(n7811), .ZN(
        n33033) );
  AOI22_X1 U4363 ( .A1(n32707), .A2(n7797), .B1(n32706), .B2(n7789), .ZN(
        n33032) );
  NAND4_X1 U4364 ( .A1(n33035), .A2(n33034), .A3(n33033), .A4(n33032), .ZN(
        n33041) );
  AOI22_X1 U4365 ( .A1(n32709), .A2(n7787), .B1(n32708), .B2(n7816), .ZN(
        n33039) );
  AOI22_X1 U4366 ( .A1(n32711), .A2(n7815), .B1(n32710), .B2(n7801), .ZN(
        n33038) );
  AOI22_X1 U4367 ( .A1(n32713), .A2(n7805), .B1(n32712), .B2(n7791), .ZN(
        n33037) );
  AOI22_X1 U4368 ( .A1(n32715), .A2(n7813), .B1(n32714), .B2(n7807), .ZN(
        n33036) );
  NAND4_X1 U4369 ( .A1(n33039), .A2(n33038), .A3(n33037), .A4(n33036), .ZN(
        n33040) );
  NOR4_X1 U4370 ( .A1(n33043), .A2(n33042), .A3(n33041), .A4(n33040), .ZN(
        n33044) );
  OAI22_X1 U4371 ( .A1(n33044), .A2(n33476), .B1(n33475), .B2(n14136), .ZN(
        n5789) );
  AOI22_X1 U4372 ( .A1(n33424), .A2(n7840), .B1(n32684), .B2(n7832), .ZN(
        n33048) );
  AOI22_X1 U4373 ( .A1(n32687), .A2(n7846), .B1(n32686), .B2(n7836), .ZN(
        n33047) );
  AOI22_X1 U4374 ( .A1(n33428), .A2(n7842), .B1(n32688), .B2(n7841), .ZN(
        n33046) );
  AOI22_X1 U4375 ( .A1(n33430), .A2(n7835), .B1(n32690), .B2(n7838), .ZN(
        n33045) );
  NAND4_X1 U4376 ( .A1(n33048), .A2(n33047), .A3(n33046), .A4(n33045), .ZN(
        n33064) );
  AOI22_X1 U4377 ( .A1(n32693), .A2(n7820), .B1(n32692), .B2(n7826), .ZN(
        n33052) );
  AOI22_X1 U4378 ( .A1(n32695), .A2(n7828), .B1(n32694), .B2(n7824), .ZN(
        n33051) );
  AOI22_X1 U4379 ( .A1(n33440), .A2(n7818), .B1(n32696), .B2(n7825), .ZN(
        n33050) );
  AOI22_X1 U4380 ( .A1(n33442), .A2(n7830), .B1(n32698), .B2(n7822), .ZN(
        n33049) );
  NAND4_X1 U4381 ( .A1(n33052), .A2(n33051), .A3(n33050), .A4(n33049), .ZN(
        n33063) );
  AOI22_X1 U4382 ( .A1(n32701), .A2(n7827), .B1(n32700), .B2(n7844), .ZN(
        n33056) );
  AOI22_X1 U4383 ( .A1(n32703), .A2(n7834), .B1(n32702), .B2(n7831), .ZN(
        n33055) );
  AOI22_X1 U4384 ( .A1(n32705), .A2(n7817), .B1(n32704), .B2(n7843), .ZN(
        n33054) );
  AOI22_X1 U4385 ( .A1(n32707), .A2(n7829), .B1(n32706), .B2(n7821), .ZN(
        n33053) );
  NAND4_X1 U4386 ( .A1(n33056), .A2(n33055), .A3(n33054), .A4(n33053), .ZN(
        n33062) );
  AOI22_X1 U4387 ( .A1(n32709), .A2(n7819), .B1(n32708), .B2(n7848), .ZN(
        n33060) );
  AOI22_X1 U4388 ( .A1(n32711), .A2(n7847), .B1(n32710), .B2(n7833), .ZN(
        n33059) );
  AOI22_X1 U4389 ( .A1(n32713), .A2(n7837), .B1(n32712), .B2(n7823), .ZN(
        n33058) );
  AOI22_X1 U4390 ( .A1(n32715), .A2(n7845), .B1(n32714), .B2(n7839), .ZN(
        n33057) );
  NAND4_X1 U4391 ( .A1(n33060), .A2(n33059), .A3(n33058), .A4(n33057), .ZN(
        n33061) );
  NOR4_X1 U4392 ( .A1(n33064), .A2(n33063), .A3(n33062), .A4(n33061), .ZN(
        n33065) );
  OAI22_X1 U4393 ( .A1(n33065), .A2(n33476), .B1(n33475), .B2(n14137), .ZN(
        n5790) );
  AOI22_X1 U4394 ( .A1(n33424), .A2(n7872), .B1(n32684), .B2(n7864), .ZN(
        n33069) );
  AOI22_X1 U4395 ( .A1(n33426), .A2(n7878), .B1(n32686), .B2(n7868), .ZN(
        n33068) );
  AOI22_X1 U4396 ( .A1(n33428), .A2(n7874), .B1(n32688), .B2(n7873), .ZN(
        n33067) );
  AOI22_X1 U4397 ( .A1(n33430), .A2(n7867), .B1(n32690), .B2(n7870), .ZN(
        n33066) );
  NAND4_X1 U4398 ( .A1(n33069), .A2(n33068), .A3(n33067), .A4(n33066), .ZN(
        n33085) );
  AOI22_X1 U4399 ( .A1(n32693), .A2(n7852), .B1(n32692), .B2(n7858), .ZN(
        n33073) );
  AOI22_X1 U4400 ( .A1(n32695), .A2(n7860), .B1(n32694), .B2(n7856), .ZN(
        n33072) );
  AOI22_X1 U4401 ( .A1(n33440), .A2(n7850), .B1(n32696), .B2(n7857), .ZN(
        n33071) );
  AOI22_X1 U4402 ( .A1(n33442), .A2(n7862), .B1(n32698), .B2(n7854), .ZN(
        n33070) );
  NAND4_X1 U4403 ( .A1(n33073), .A2(n33072), .A3(n33071), .A4(n33070), .ZN(
        n33084) );
  AOI22_X1 U4404 ( .A1(n32701), .A2(n7859), .B1(n32700), .B2(n7876), .ZN(
        n33077) );
  AOI22_X1 U4405 ( .A1(n33450), .A2(n7866), .B1(n32702), .B2(n7863), .ZN(
        n33076) );
  AOI22_X1 U4406 ( .A1(n33452), .A2(n7849), .B1(n32704), .B2(n7875), .ZN(
        n33075) );
  AOI22_X1 U4407 ( .A1(n33454), .A2(n7861), .B1(n32706), .B2(n7853), .ZN(
        n33074) );
  NAND4_X1 U4408 ( .A1(n33077), .A2(n33076), .A3(n33075), .A4(n33074), .ZN(
        n33083) );
  AOI22_X1 U4409 ( .A1(n32709), .A2(n7851), .B1(n32708), .B2(n7880), .ZN(
        n33081) );
  AOI22_X1 U4410 ( .A1(n33462), .A2(n7879), .B1(n32710), .B2(n7865), .ZN(
        n33080) );
  AOI22_X1 U4411 ( .A1(n33464), .A2(n7869), .B1(n32712), .B2(n7855), .ZN(
        n33079) );
  AOI22_X1 U4412 ( .A1(n32715), .A2(n7877), .B1(n32714), .B2(n7871), .ZN(
        n33078) );
  NAND4_X1 U4413 ( .A1(n33081), .A2(n33080), .A3(n33079), .A4(n33078), .ZN(
        n33082) );
  NOR4_X1 U4414 ( .A1(n33085), .A2(n33084), .A3(n33083), .A4(n33082), .ZN(
        n33086) );
  OAI22_X1 U4415 ( .A1(n33086), .A2(n33476), .B1(n33475), .B2(n32729), .ZN(
        n5791) );
  AOI22_X1 U4416 ( .A1(n33424), .A2(n7904), .B1(n32684), .B2(n7896), .ZN(
        n33090) );
  AOI22_X1 U4417 ( .A1(n33426), .A2(n7910), .B1(n32686), .B2(n7900), .ZN(
        n33089) );
  AOI22_X1 U4418 ( .A1(n33428), .A2(n7906), .B1(n32688), .B2(n7905), .ZN(
        n33088) );
  AOI22_X1 U4419 ( .A1(n33430), .A2(n7899), .B1(n32690), .B2(n7902), .ZN(
        n33087) );
  NAND4_X1 U4420 ( .A1(n33090), .A2(n33089), .A3(n33088), .A4(n33087), .ZN(
        n33106) );
  AOI22_X1 U4421 ( .A1(n33436), .A2(n7884), .B1(n32692), .B2(n7890), .ZN(
        n33094) );
  AOI22_X1 U4422 ( .A1(n33438), .A2(n7892), .B1(n32694), .B2(n7888), .ZN(
        n33093) );
  AOI22_X1 U4423 ( .A1(n33440), .A2(n7882), .B1(n32696), .B2(n7889), .ZN(
        n33092) );
  AOI22_X1 U4424 ( .A1(n33442), .A2(n7894), .B1(n32698), .B2(n7886), .ZN(
        n33091) );
  NAND4_X1 U4425 ( .A1(n33094), .A2(n33093), .A3(n33092), .A4(n33091), .ZN(
        n33105) );
  AOI22_X1 U4426 ( .A1(n33448), .A2(n7891), .B1(n32700), .B2(n7908), .ZN(
        n33098) );
  AOI22_X1 U4427 ( .A1(n33450), .A2(n7898), .B1(n32702), .B2(n7895), .ZN(
        n33097) );
  AOI22_X1 U4428 ( .A1(n33452), .A2(n7881), .B1(n32704), .B2(n7907), .ZN(
        n33096) );
  AOI22_X1 U4429 ( .A1(n33454), .A2(n7893), .B1(n32706), .B2(n7885), .ZN(
        n33095) );
  NAND4_X1 U4430 ( .A1(n33098), .A2(n33097), .A3(n33096), .A4(n33095), .ZN(
        n33104) );
  AOI22_X1 U4431 ( .A1(n33460), .A2(n7883), .B1(n32708), .B2(n7912), .ZN(
        n33102) );
  AOI22_X1 U4432 ( .A1(n33462), .A2(n7911), .B1(n32710), .B2(n7897), .ZN(
        n33101) );
  AOI22_X1 U4433 ( .A1(n33464), .A2(n7901), .B1(n32712), .B2(n7887), .ZN(
        n33100) );
  AOI22_X1 U4434 ( .A1(n33466), .A2(n7909), .B1(n32714), .B2(n7903), .ZN(
        n33099) );
  NAND4_X1 U4435 ( .A1(n33102), .A2(n33101), .A3(n33100), .A4(n33099), .ZN(
        n33103) );
  NOR4_X1 U4436 ( .A1(n33106), .A2(n33105), .A3(n33104), .A4(n33103), .ZN(
        n33107) );
  OAI22_X1 U4437 ( .A1(n33107), .A2(n33476), .B1(n33475), .B2(n32728), .ZN(
        n5792) );
  AOI22_X1 U4438 ( .A1(n33424), .A2(n7936), .B1(n32684), .B2(n7928), .ZN(
        n33111) );
  AOI22_X1 U4439 ( .A1(n33426), .A2(n7942), .B1(n32686), .B2(n7932), .ZN(
        n33110) );
  AOI22_X1 U4440 ( .A1(n33428), .A2(n7938), .B1(n32688), .B2(n7937), .ZN(
        n33109) );
  AOI22_X1 U4441 ( .A1(n33430), .A2(n7931), .B1(n32690), .B2(n7934), .ZN(
        n33108) );
  NAND4_X1 U4442 ( .A1(n33111), .A2(n33110), .A3(n33109), .A4(n33108), .ZN(
        n33127) );
  AOI22_X1 U4443 ( .A1(n33436), .A2(n7916), .B1(n32692), .B2(n7922), .ZN(
        n33115) );
  AOI22_X1 U4444 ( .A1(n33438), .A2(n7924), .B1(n32694), .B2(n7920), .ZN(
        n33114) );
  AOI22_X1 U4445 ( .A1(n33440), .A2(n7914), .B1(n32696), .B2(n7921), .ZN(
        n33113) );
  AOI22_X1 U4446 ( .A1(n33442), .A2(n7926), .B1(n32698), .B2(n7918), .ZN(
        n33112) );
  NAND4_X1 U4447 ( .A1(n33115), .A2(n33114), .A3(n33113), .A4(n33112), .ZN(
        n33126) );
  AOI22_X1 U4448 ( .A1(n33448), .A2(n7923), .B1(n32700), .B2(n7940), .ZN(
        n33119) );
  AOI22_X1 U4449 ( .A1(n33450), .A2(n7930), .B1(n32702), .B2(n7927), .ZN(
        n33118) );
  AOI22_X1 U4450 ( .A1(n33452), .A2(n7913), .B1(n32704), .B2(n7939), .ZN(
        n33117) );
  AOI22_X1 U4451 ( .A1(n33454), .A2(n7925), .B1(n32706), .B2(n7917), .ZN(
        n33116) );
  NAND4_X1 U4452 ( .A1(n33119), .A2(n33118), .A3(n33117), .A4(n33116), .ZN(
        n33125) );
  AOI22_X1 U4453 ( .A1(n33460), .A2(n7915), .B1(n32708), .B2(n7944), .ZN(
        n33123) );
  AOI22_X1 U4454 ( .A1(n33462), .A2(n7943), .B1(n32710), .B2(n7929), .ZN(
        n33122) );
  AOI22_X1 U4455 ( .A1(n33464), .A2(n7933), .B1(n32712), .B2(n7919), .ZN(
        n33121) );
  AOI22_X1 U4456 ( .A1(n33466), .A2(n7941), .B1(n32714), .B2(n7935), .ZN(
        n33120) );
  NAND4_X1 U4457 ( .A1(n33123), .A2(n33122), .A3(n33121), .A4(n33120), .ZN(
        n33124) );
  NOR4_X1 U4458 ( .A1(n33127), .A2(n33126), .A3(n33125), .A4(n33124), .ZN(
        n33128) );
  OAI22_X1 U4459 ( .A1(n33128), .A2(n33476), .B1(n33475), .B2(n14140), .ZN(
        n5793) );
  AOI22_X1 U4460 ( .A1(n32685), .A2(n7968), .B1(n32684), .B2(n7960), .ZN(
        n33132) );
  AOI22_X1 U4461 ( .A1(n33426), .A2(n7974), .B1(n32686), .B2(n7964), .ZN(
        n33131) );
  AOI22_X1 U4462 ( .A1(n32689), .A2(n7970), .B1(n32688), .B2(n7969), .ZN(
        n33130) );
  AOI22_X1 U4463 ( .A1(n32691), .A2(n7963), .B1(n32690), .B2(n7966), .ZN(
        n33129) );
  NAND4_X1 U4464 ( .A1(n33132), .A2(n33131), .A3(n33130), .A4(n33129), .ZN(
        n33148) );
  AOI22_X1 U4465 ( .A1(n33436), .A2(n7948), .B1(n32692), .B2(n7954), .ZN(
        n33136) );
  AOI22_X1 U4466 ( .A1(n33438), .A2(n7956), .B1(n32694), .B2(n7952), .ZN(
        n33135) );
  AOI22_X1 U4467 ( .A1(n32697), .A2(n7946), .B1(n32696), .B2(n7953), .ZN(
        n33134) );
  AOI22_X1 U4468 ( .A1(n32699), .A2(n7958), .B1(n32698), .B2(n7950), .ZN(
        n33133) );
  NAND4_X1 U4469 ( .A1(n33136), .A2(n33135), .A3(n33134), .A4(n33133), .ZN(
        n33147) );
  AOI22_X1 U4470 ( .A1(n33448), .A2(n7955), .B1(n32700), .B2(n7972), .ZN(
        n33140) );
  AOI22_X1 U4471 ( .A1(n33450), .A2(n7962), .B1(n32702), .B2(n7959), .ZN(
        n33139) );
  AOI22_X1 U4472 ( .A1(n33452), .A2(n7945), .B1(n32704), .B2(n7971), .ZN(
        n33138) );
  AOI22_X1 U4473 ( .A1(n33454), .A2(n7957), .B1(n32706), .B2(n7949), .ZN(
        n33137) );
  NAND4_X1 U4474 ( .A1(n33140), .A2(n33139), .A3(n33138), .A4(n33137), .ZN(
        n33146) );
  AOI22_X1 U4475 ( .A1(n33460), .A2(n7947), .B1(n32708), .B2(n7976), .ZN(
        n33144) );
  AOI22_X1 U4476 ( .A1(n33462), .A2(n7975), .B1(n32710), .B2(n7961), .ZN(
        n33143) );
  AOI22_X1 U4477 ( .A1(n33464), .A2(n7965), .B1(n32712), .B2(n7951), .ZN(
        n33142) );
  AOI22_X1 U4478 ( .A1(n33466), .A2(n7973), .B1(n32714), .B2(n7967), .ZN(
        n33141) );
  NAND4_X1 U4479 ( .A1(n33144), .A2(n33143), .A3(n33142), .A4(n33141), .ZN(
        n33145) );
  NOR4_X1 U4480 ( .A1(n33148), .A2(n33147), .A3(n33146), .A4(n33145), .ZN(
        n33149) );
  OAI22_X1 U4481 ( .A1(n33149), .A2(n33476), .B1(n33475), .B2(n14141), .ZN(
        n5794) );
  AOI22_X1 U4482 ( .A1(n33424), .A2(n8000), .B1(n32684), .B2(n7992), .ZN(
        n33153) );
  AOI22_X1 U4483 ( .A1(n33426), .A2(n8006), .B1(n32686), .B2(n7996), .ZN(
        n33152) );
  AOI22_X1 U4484 ( .A1(n33428), .A2(n8002), .B1(n32688), .B2(n8001), .ZN(
        n33151) );
  AOI22_X1 U4485 ( .A1(n33430), .A2(n7995), .B1(n32690), .B2(n7998), .ZN(
        n33150) );
  NAND4_X1 U4486 ( .A1(n33153), .A2(n33152), .A3(n33151), .A4(n33150), .ZN(
        n33169) );
  AOI22_X1 U4487 ( .A1(n33436), .A2(n7980), .B1(n32692), .B2(n7986), .ZN(
        n33157) );
  AOI22_X1 U4488 ( .A1(n33438), .A2(n7988), .B1(n32694), .B2(n7984), .ZN(
        n33156) );
  AOI22_X1 U4489 ( .A1(n33440), .A2(n7978), .B1(n32696), .B2(n7985), .ZN(
        n33155) );
  AOI22_X1 U4490 ( .A1(n33442), .A2(n7990), .B1(n32698), .B2(n7982), .ZN(
        n33154) );
  NAND4_X1 U4491 ( .A1(n33157), .A2(n33156), .A3(n33155), .A4(n33154), .ZN(
        n33168) );
  AOI22_X1 U4492 ( .A1(n33448), .A2(n7987), .B1(n32700), .B2(n8004), .ZN(
        n33161) );
  AOI22_X1 U4493 ( .A1(n32703), .A2(n7994), .B1(n32702), .B2(n7991), .ZN(
        n33160) );
  AOI22_X1 U4494 ( .A1(n33452), .A2(n7977), .B1(n32704), .B2(n8003), .ZN(
        n33159) );
  AOI22_X1 U4495 ( .A1(n32707), .A2(n7989), .B1(n32706), .B2(n7981), .ZN(
        n33158) );
  NAND4_X1 U4496 ( .A1(n33161), .A2(n33160), .A3(n33159), .A4(n33158), .ZN(
        n33167) );
  AOI22_X1 U4497 ( .A1(n33460), .A2(n7979), .B1(n32708), .B2(n8008), .ZN(
        n33165) );
  AOI22_X1 U4498 ( .A1(n32711), .A2(n8007), .B1(n32710), .B2(n7993), .ZN(
        n33164) );
  AOI22_X1 U4499 ( .A1(n33464), .A2(n7997), .B1(n32712), .B2(n7983), .ZN(
        n33163) );
  AOI22_X1 U4500 ( .A1(n33466), .A2(n8005), .B1(n32714), .B2(n7999), .ZN(
        n33162) );
  NAND4_X1 U4501 ( .A1(n33165), .A2(n33164), .A3(n33163), .A4(n33162), .ZN(
        n33166) );
  NOR4_X1 U4502 ( .A1(n33169), .A2(n33168), .A3(n33167), .A4(n33166), .ZN(
        n33170) );
  OAI22_X1 U4503 ( .A1(n33170), .A2(n33476), .B1(n33475), .B2(n14142), .ZN(
        n5795) );
  AOI22_X1 U4504 ( .A1(n32685), .A2(n8032), .B1(n33423), .B2(n8024), .ZN(
        n33174) );
  AOI22_X1 U4505 ( .A1(n32687), .A2(n8038), .B1(n33425), .B2(n8028), .ZN(
        n33173) );
  AOI22_X1 U4506 ( .A1(n32689), .A2(n8034), .B1(n33427), .B2(n8033), .ZN(
        n33172) );
  AOI22_X1 U4507 ( .A1(n32691), .A2(n8027), .B1(n33429), .B2(n8030), .ZN(
        n33171) );
  NAND4_X1 U4508 ( .A1(n33174), .A2(n33173), .A3(n33172), .A4(n33171), .ZN(
        n33190) );
  AOI22_X1 U4509 ( .A1(n32693), .A2(n8012), .B1(n33435), .B2(n8018), .ZN(
        n33178) );
  AOI22_X1 U4510 ( .A1(n32695), .A2(n8020), .B1(n33437), .B2(n8016), .ZN(
        n33177) );
  AOI22_X1 U4511 ( .A1(n32697), .A2(n8010), .B1(n33439), .B2(n8017), .ZN(
        n33176) );
  AOI22_X1 U4512 ( .A1(n32699), .A2(n8022), .B1(n33441), .B2(n8014), .ZN(
        n33175) );
  NAND4_X1 U4513 ( .A1(n33178), .A2(n33177), .A3(n33176), .A4(n33175), .ZN(
        n33189) );
  AOI22_X1 U4514 ( .A1(n33448), .A2(n8019), .B1(n32700), .B2(n8036), .ZN(
        n33182) );
  AOI22_X1 U4515 ( .A1(n32703), .A2(n8026), .B1(n33449), .B2(n8023), .ZN(
        n33181) );
  AOI22_X1 U4516 ( .A1(n32705), .A2(n8009), .B1(n33451), .B2(n8035), .ZN(
        n33180) );
  AOI22_X1 U4517 ( .A1(n33454), .A2(n8021), .B1(n32706), .B2(n8013), .ZN(
        n33179) );
  NAND4_X1 U4518 ( .A1(n33182), .A2(n33181), .A3(n33180), .A4(n33179), .ZN(
        n33188) );
  AOI22_X1 U4519 ( .A1(n32709), .A2(n8011), .B1(n32708), .B2(n8040), .ZN(
        n33186) );
  AOI22_X1 U4520 ( .A1(n32711), .A2(n8039), .B1(n33461), .B2(n8025), .ZN(
        n33185) );
  AOI22_X1 U4521 ( .A1(n32713), .A2(n8029), .B1(n33463), .B2(n8015), .ZN(
        n33184) );
  AOI22_X1 U4522 ( .A1(n33466), .A2(n8037), .B1(n32714), .B2(n8031), .ZN(
        n33183) );
  NAND4_X1 U4523 ( .A1(n33186), .A2(n33185), .A3(n33184), .A4(n33183), .ZN(
        n33187) );
  NOR4_X1 U4524 ( .A1(n33190), .A2(n33189), .A3(n33188), .A4(n33187), .ZN(
        n33191) );
  OAI22_X1 U4525 ( .A1(n33191), .A2(n33476), .B1(n33475), .B2(n14143), .ZN(
        n5796) );
  AOI22_X1 U4526 ( .A1(n32685), .A2(n8064), .B1(n33423), .B2(n8056), .ZN(
        n33195) );
  AOI22_X1 U4527 ( .A1(n32687), .A2(n8070), .B1(n33425), .B2(n8060), .ZN(
        n33194) );
  AOI22_X1 U4528 ( .A1(n32689), .A2(n8066), .B1(n33427), .B2(n8065), .ZN(
        n33193) );
  AOI22_X1 U4529 ( .A1(n32691), .A2(n8059), .B1(n33429), .B2(n8062), .ZN(
        n33192) );
  NAND4_X1 U4530 ( .A1(n33195), .A2(n33194), .A3(n33193), .A4(n33192), .ZN(
        n33211) );
  AOI22_X1 U4531 ( .A1(n32693), .A2(n8044), .B1(n33435), .B2(n8050), .ZN(
        n33199) );
  AOI22_X1 U4532 ( .A1(n32695), .A2(n8052), .B1(n33437), .B2(n8048), .ZN(
        n33198) );
  AOI22_X1 U4533 ( .A1(n32697), .A2(n8042), .B1(n33439), .B2(n8049), .ZN(
        n33197) );
  AOI22_X1 U4534 ( .A1(n32699), .A2(n8054), .B1(n33441), .B2(n8046), .ZN(
        n33196) );
  NAND4_X1 U4535 ( .A1(n33199), .A2(n33198), .A3(n33197), .A4(n33196), .ZN(
        n33210) );
  AOI22_X1 U4536 ( .A1(n32701), .A2(n8051), .B1(n33447), .B2(n8068), .ZN(
        n33203) );
  AOI22_X1 U4537 ( .A1(n32703), .A2(n8058), .B1(n33449), .B2(n8055), .ZN(
        n33202) );
  AOI22_X1 U4538 ( .A1(n32705), .A2(n8041), .B1(n33451), .B2(n8067), .ZN(
        n33201) );
  AOI22_X1 U4539 ( .A1(n32707), .A2(n8053), .B1(n33453), .B2(n8045), .ZN(
        n33200) );
  NAND4_X1 U4540 ( .A1(n33203), .A2(n33202), .A3(n33201), .A4(n33200), .ZN(
        n33209) );
  AOI22_X1 U4541 ( .A1(n32709), .A2(n8043), .B1(n33459), .B2(n8072), .ZN(
        n33207) );
  AOI22_X1 U4542 ( .A1(n32711), .A2(n8071), .B1(n33461), .B2(n8057), .ZN(
        n33206) );
  AOI22_X1 U4543 ( .A1(n32713), .A2(n8061), .B1(n33463), .B2(n8047), .ZN(
        n33205) );
  AOI22_X1 U4544 ( .A1(n32715), .A2(n8069), .B1(n33465), .B2(n8063), .ZN(
        n33204) );
  NAND4_X1 U4545 ( .A1(n33207), .A2(n33206), .A3(n33205), .A4(n33204), .ZN(
        n33208) );
  NOR4_X1 U4546 ( .A1(n33211), .A2(n33210), .A3(n33209), .A4(n33208), .ZN(
        n33212) );
  OAI22_X1 U4547 ( .A1(n33212), .A2(n33476), .B1(n33475), .B2(n14144), .ZN(
        n5797) );
  AOI22_X1 U4548 ( .A1(n32685), .A2(n8096), .B1(n33423), .B2(n8088), .ZN(
        n33216) );
  AOI22_X1 U4549 ( .A1(n32687), .A2(n8102), .B1(n33425), .B2(n8092), .ZN(
        n33215) );
  AOI22_X1 U4550 ( .A1(n32689), .A2(n8098), .B1(n33427), .B2(n8097), .ZN(
        n33214) );
  AOI22_X1 U4551 ( .A1(n32691), .A2(n8091), .B1(n33429), .B2(n8094), .ZN(
        n33213) );
  NAND4_X1 U4552 ( .A1(n33216), .A2(n33215), .A3(n33214), .A4(n33213), .ZN(
        n33232) );
  AOI22_X1 U4553 ( .A1(n32693), .A2(n8076), .B1(n33435), .B2(n8082), .ZN(
        n33220) );
  AOI22_X1 U4554 ( .A1(n32695), .A2(n8084), .B1(n33437), .B2(n8080), .ZN(
        n33219) );
  AOI22_X1 U4555 ( .A1(n32697), .A2(n8074), .B1(n33439), .B2(n8081), .ZN(
        n33218) );
  AOI22_X1 U4556 ( .A1(n32699), .A2(n8086), .B1(n33441), .B2(n8078), .ZN(
        n33217) );
  NAND4_X1 U4557 ( .A1(n33220), .A2(n33219), .A3(n33218), .A4(n33217), .ZN(
        n33231) );
  AOI22_X1 U4558 ( .A1(n32701), .A2(n8083), .B1(n33447), .B2(n8100), .ZN(
        n33224) );
  AOI22_X1 U4559 ( .A1(n32703), .A2(n8090), .B1(n33449), .B2(n8087), .ZN(
        n33223) );
  AOI22_X1 U4560 ( .A1(n32705), .A2(n8073), .B1(n33451), .B2(n8099), .ZN(
        n33222) );
  AOI22_X1 U4561 ( .A1(n32707), .A2(n8085), .B1(n33453), .B2(n8077), .ZN(
        n33221) );
  NAND4_X1 U4562 ( .A1(n33224), .A2(n33223), .A3(n33222), .A4(n33221), .ZN(
        n33230) );
  AOI22_X1 U4563 ( .A1(n32709), .A2(n8075), .B1(n33459), .B2(n8104), .ZN(
        n33228) );
  AOI22_X1 U4564 ( .A1(n32711), .A2(n8103), .B1(n33461), .B2(n8089), .ZN(
        n33227) );
  AOI22_X1 U4565 ( .A1(n32713), .A2(n8093), .B1(n33463), .B2(n8079), .ZN(
        n33226) );
  AOI22_X1 U4566 ( .A1(n32715), .A2(n8101), .B1(n33465), .B2(n8095), .ZN(
        n33225) );
  NAND4_X1 U4567 ( .A1(n33228), .A2(n33227), .A3(n33226), .A4(n33225), .ZN(
        n33229) );
  NOR4_X1 U4568 ( .A1(n33232), .A2(n33231), .A3(n33230), .A4(n33229), .ZN(
        n33233) );
  OAI22_X1 U4569 ( .A1(n33233), .A2(n33476), .B1(n33475), .B2(n14145), .ZN(
        n5798) );
  AOI22_X1 U4570 ( .A1(n32685), .A2(n8128), .B1(n33423), .B2(n8120), .ZN(
        n33237) );
  AOI22_X1 U4571 ( .A1(n32687), .A2(n8134), .B1(n33425), .B2(n8124), .ZN(
        n33236) );
  AOI22_X1 U4572 ( .A1(n32689), .A2(n8130), .B1(n33427), .B2(n8129), .ZN(
        n33235) );
  AOI22_X1 U4573 ( .A1(n32691), .A2(n8123), .B1(n33429), .B2(n8126), .ZN(
        n33234) );
  NAND4_X1 U4574 ( .A1(n33237), .A2(n33236), .A3(n33235), .A4(n33234), .ZN(
        n33253) );
  AOI22_X1 U4575 ( .A1(n32693), .A2(n8108), .B1(n33435), .B2(n8114), .ZN(
        n33241) );
  AOI22_X1 U4576 ( .A1(n32695), .A2(n8116), .B1(n33437), .B2(n8112), .ZN(
        n33240) );
  AOI22_X1 U4577 ( .A1(n32697), .A2(n8106), .B1(n33439), .B2(n8113), .ZN(
        n33239) );
  AOI22_X1 U4578 ( .A1(n32699), .A2(n8118), .B1(n33441), .B2(n8110), .ZN(
        n33238) );
  NAND4_X1 U4579 ( .A1(n33241), .A2(n33240), .A3(n33239), .A4(n33238), .ZN(
        n33252) );
  AOI22_X1 U4580 ( .A1(n32701), .A2(n8115), .B1(n33447), .B2(n8132), .ZN(
        n33245) );
  AOI22_X1 U4581 ( .A1(n32703), .A2(n8122), .B1(n33449), .B2(n8119), .ZN(
        n33244) );
  AOI22_X1 U4582 ( .A1(n32705), .A2(n8105), .B1(n33451), .B2(n8131), .ZN(
        n33243) );
  AOI22_X1 U4583 ( .A1(n32707), .A2(n8117), .B1(n33453), .B2(n8109), .ZN(
        n33242) );
  NAND4_X1 U4584 ( .A1(n33245), .A2(n33244), .A3(n33243), .A4(n33242), .ZN(
        n33251) );
  AOI22_X1 U4585 ( .A1(n32709), .A2(n8107), .B1(n33459), .B2(n8136), .ZN(
        n33249) );
  AOI22_X1 U4586 ( .A1(n32711), .A2(n8135), .B1(n33461), .B2(n8121), .ZN(
        n33248) );
  AOI22_X1 U4587 ( .A1(n32713), .A2(n8125), .B1(n33463), .B2(n8111), .ZN(
        n33247) );
  AOI22_X1 U4588 ( .A1(n32715), .A2(n8133), .B1(n33465), .B2(n8127), .ZN(
        n33246) );
  NAND4_X1 U4589 ( .A1(n33249), .A2(n33248), .A3(n33247), .A4(n33246), .ZN(
        n33250) );
  NOR4_X1 U4590 ( .A1(n33253), .A2(n33252), .A3(n33251), .A4(n33250), .ZN(
        n33254) );
  OAI22_X1 U4591 ( .A1(n33254), .A2(n33476), .B1(n33475), .B2(n32727), .ZN(
        n5799) );
  AOI22_X1 U4592 ( .A1(n32685), .A2(n8160), .B1(n33423), .B2(n8152), .ZN(
        n33258) );
  AOI22_X1 U4593 ( .A1(n32687), .A2(n8166), .B1(n33425), .B2(n8156), .ZN(
        n33257) );
  AOI22_X1 U4594 ( .A1(n32689), .A2(n8162), .B1(n33427), .B2(n8161), .ZN(
        n33256) );
  AOI22_X1 U4595 ( .A1(n32691), .A2(n8155), .B1(n33429), .B2(n8158), .ZN(
        n33255) );
  NAND4_X1 U4596 ( .A1(n33258), .A2(n33257), .A3(n33256), .A4(n33255), .ZN(
        n33274) );
  AOI22_X1 U4597 ( .A1(n33436), .A2(n8140), .B1(n32692), .B2(n8146), .ZN(
        n33262) );
  AOI22_X1 U4598 ( .A1(n33438), .A2(n8148), .B1(n32694), .B2(n8144), .ZN(
        n33261) );
  AOI22_X1 U4599 ( .A1(n32697), .A2(n8138), .B1(n33439), .B2(n8145), .ZN(
        n33260) );
  AOI22_X1 U4600 ( .A1(n32699), .A2(n8150), .B1(n33441), .B2(n8142), .ZN(
        n33259) );
  NAND4_X1 U4601 ( .A1(n33262), .A2(n33261), .A3(n33260), .A4(n33259), .ZN(
        n33273) );
  AOI22_X1 U4602 ( .A1(n32701), .A2(n8147), .B1(n33447), .B2(n8164), .ZN(
        n33266) );
  AOI22_X1 U4603 ( .A1(n32703), .A2(n8154), .B1(n33449), .B2(n8151), .ZN(
        n33265) );
  AOI22_X1 U4604 ( .A1(n32705), .A2(n8137), .B1(n33451), .B2(n8163), .ZN(
        n33264) );
  AOI22_X1 U4605 ( .A1(n32707), .A2(n8149), .B1(n33453), .B2(n8141), .ZN(
        n33263) );
  NAND4_X1 U4606 ( .A1(n33266), .A2(n33265), .A3(n33264), .A4(n33263), .ZN(
        n33272) );
  AOI22_X1 U4607 ( .A1(n32709), .A2(n8139), .B1(n33459), .B2(n8168), .ZN(
        n33270) );
  AOI22_X1 U4608 ( .A1(n32711), .A2(n8167), .B1(n33461), .B2(n8153), .ZN(
        n33269) );
  AOI22_X1 U4609 ( .A1(n32713), .A2(n8157), .B1(n33463), .B2(n8143), .ZN(
        n33268) );
  AOI22_X1 U4610 ( .A1(n32715), .A2(n8165), .B1(n33465), .B2(n8159), .ZN(
        n33267) );
  NAND4_X1 U4611 ( .A1(n33270), .A2(n33269), .A3(n33268), .A4(n33267), .ZN(
        n33271) );
  NOR4_X1 U4612 ( .A1(n33274), .A2(n33273), .A3(n33272), .A4(n33271), .ZN(
        n33275) );
  OAI22_X1 U4613 ( .A1(n33275), .A2(n33476), .B1(n33475), .B2(n32726), .ZN(
        n5800) );
  AOI22_X1 U4614 ( .A1(n33424), .A2(n8192), .B1(n33423), .B2(n8184), .ZN(
        n33279) );
  AOI22_X1 U4615 ( .A1(n33426), .A2(n8198), .B1(n33425), .B2(n8188), .ZN(
        n33278) );
  AOI22_X1 U4616 ( .A1(n33428), .A2(n8194), .B1(n33427), .B2(n8193), .ZN(
        n33277) );
  AOI22_X1 U4617 ( .A1(n33430), .A2(n8187), .B1(n33429), .B2(n8190), .ZN(
        n33276) );
  NAND4_X1 U4618 ( .A1(n33279), .A2(n33278), .A3(n33277), .A4(n33276), .ZN(
        n33295) );
  AOI22_X1 U4619 ( .A1(n33436), .A2(n8172), .B1(n33435), .B2(n8178), .ZN(
        n33283) );
  AOI22_X1 U4620 ( .A1(n33438), .A2(n8180), .B1(n33437), .B2(n8176), .ZN(
        n33282) );
  AOI22_X1 U4621 ( .A1(n33440), .A2(n8170), .B1(n33439), .B2(n8177), .ZN(
        n33281) );
  AOI22_X1 U4622 ( .A1(n33442), .A2(n8182), .B1(n33441), .B2(n8174), .ZN(
        n33280) );
  NAND4_X1 U4623 ( .A1(n33283), .A2(n33282), .A3(n33281), .A4(n33280), .ZN(
        n33294) );
  AOI22_X1 U4624 ( .A1(n33448), .A2(n8179), .B1(n33447), .B2(n8196), .ZN(
        n33287) );
  AOI22_X1 U4625 ( .A1(n33450), .A2(n8186), .B1(n33449), .B2(n8183), .ZN(
        n33286) );
  AOI22_X1 U4626 ( .A1(n33452), .A2(n8169), .B1(n33451), .B2(n8195), .ZN(
        n33285) );
  AOI22_X1 U4627 ( .A1(n33454), .A2(n8181), .B1(n33453), .B2(n8173), .ZN(
        n33284) );
  NAND4_X1 U4628 ( .A1(n33287), .A2(n33286), .A3(n33285), .A4(n33284), .ZN(
        n33293) );
  AOI22_X1 U4629 ( .A1(n33460), .A2(n8171), .B1(n33459), .B2(n8200), .ZN(
        n33291) );
  AOI22_X1 U4630 ( .A1(n33462), .A2(n8199), .B1(n33461), .B2(n8185), .ZN(
        n33290) );
  AOI22_X1 U4631 ( .A1(n33464), .A2(n8189), .B1(n33463), .B2(n8175), .ZN(
        n33289) );
  AOI22_X1 U4632 ( .A1(n33466), .A2(n8197), .B1(n33465), .B2(n8191), .ZN(
        n33288) );
  NAND4_X1 U4633 ( .A1(n33291), .A2(n33290), .A3(n33289), .A4(n33288), .ZN(
        n33292) );
  NOR4_X1 U4634 ( .A1(n33295), .A2(n33294), .A3(n33293), .A4(n33292), .ZN(
        n33296) );
  OAI22_X1 U4635 ( .A1(n33296), .A2(n33476), .B1(n33475), .B2(n14148), .ZN(
        n5801) );
  AOI22_X1 U4636 ( .A1(n33424), .A2(n8224), .B1(n33423), .B2(n8216), .ZN(
        n33300) );
  AOI22_X1 U4637 ( .A1(n33426), .A2(n8230), .B1(n33425), .B2(n8220), .ZN(
        n33299) );
  AOI22_X1 U4638 ( .A1(n33428), .A2(n8226), .B1(n33427), .B2(n8225), .ZN(
        n33298) );
  AOI22_X1 U4639 ( .A1(n33430), .A2(n8219), .B1(n33429), .B2(n8222), .ZN(
        n33297) );
  NAND4_X1 U4640 ( .A1(n33300), .A2(n33299), .A3(n33298), .A4(n33297), .ZN(
        n33316) );
  AOI22_X1 U4641 ( .A1(n33436), .A2(n8204), .B1(n33435), .B2(n8210), .ZN(
        n33304) );
  AOI22_X1 U4642 ( .A1(n33438), .A2(n8212), .B1(n33437), .B2(n8208), .ZN(
        n33303) );
  AOI22_X1 U4643 ( .A1(n33440), .A2(n8202), .B1(n33439), .B2(n8209), .ZN(
        n33302) );
  AOI22_X1 U4644 ( .A1(n33442), .A2(n8214), .B1(n33441), .B2(n8206), .ZN(
        n33301) );
  NAND4_X1 U4645 ( .A1(n33304), .A2(n33303), .A3(n33302), .A4(n33301), .ZN(
        n33315) );
  AOI22_X1 U4646 ( .A1(n33448), .A2(n8211), .B1(n33447), .B2(n8228), .ZN(
        n33308) );
  AOI22_X1 U4647 ( .A1(n33450), .A2(n8218), .B1(n33449), .B2(n8215), .ZN(
        n33307) );
  AOI22_X1 U4648 ( .A1(n33452), .A2(n8201), .B1(n33451), .B2(n8227), .ZN(
        n33306) );
  AOI22_X1 U4649 ( .A1(n33454), .A2(n8213), .B1(n33453), .B2(n8205), .ZN(
        n33305) );
  NAND4_X1 U4650 ( .A1(n33308), .A2(n33307), .A3(n33306), .A4(n33305), .ZN(
        n33314) );
  AOI22_X1 U4651 ( .A1(n33460), .A2(n8203), .B1(n33459), .B2(n8232), .ZN(
        n33312) );
  AOI22_X1 U4652 ( .A1(n33462), .A2(n8231), .B1(n33461), .B2(n8217), .ZN(
        n33311) );
  AOI22_X1 U4653 ( .A1(n33464), .A2(n8221), .B1(n33463), .B2(n8207), .ZN(
        n33310) );
  AOI22_X1 U4654 ( .A1(n33466), .A2(n8229), .B1(n33465), .B2(n8223), .ZN(
        n33309) );
  NAND4_X1 U4655 ( .A1(n33312), .A2(n33311), .A3(n33310), .A4(n33309), .ZN(
        n33313) );
  NOR4_X1 U4656 ( .A1(n33316), .A2(n33315), .A3(n33314), .A4(n33313), .ZN(
        n33317) );
  OAI22_X1 U4657 ( .A1(n33317), .A2(n33476), .B1(n33475), .B2(n14149), .ZN(
        n5802) );
  AOI22_X1 U4658 ( .A1(n32685), .A2(n8256), .B1(n33423), .B2(n8248), .ZN(
        n33321) );
  AOI22_X1 U4659 ( .A1(n33426), .A2(n8262), .B1(n33425), .B2(n8252), .ZN(
        n33320) );
  AOI22_X1 U4660 ( .A1(n33428), .A2(n8258), .B1(n33427), .B2(n8257), .ZN(
        n33319) );
  AOI22_X1 U4661 ( .A1(n33430), .A2(n8251), .B1(n33429), .B2(n8254), .ZN(
        n33318) );
  NAND4_X1 U4662 ( .A1(n33321), .A2(n33320), .A3(n33319), .A4(n33318), .ZN(
        n33337) );
  AOI22_X1 U4663 ( .A1(n33436), .A2(n8236), .B1(n33435), .B2(n8242), .ZN(
        n33325) );
  AOI22_X1 U4664 ( .A1(n33438), .A2(n8244), .B1(n33437), .B2(n8240), .ZN(
        n33324) );
  AOI22_X1 U4665 ( .A1(n32697), .A2(n8234), .B1(n32696), .B2(n8241), .ZN(
        n33323) );
  AOI22_X1 U4666 ( .A1(n33442), .A2(n8246), .B1(n33441), .B2(n8238), .ZN(
        n33322) );
  NAND4_X1 U4667 ( .A1(n33325), .A2(n33324), .A3(n33323), .A4(n33322), .ZN(
        n33336) );
  AOI22_X1 U4668 ( .A1(n32701), .A2(n8243), .B1(n33447), .B2(n8260), .ZN(
        n33329) );
  AOI22_X1 U4669 ( .A1(n32703), .A2(n8250), .B1(n32702), .B2(n8247), .ZN(
        n33328) );
  AOI22_X1 U4670 ( .A1(n32705), .A2(n8233), .B1(n32704), .B2(n8259), .ZN(
        n33327) );
  AOI22_X1 U4671 ( .A1(n33454), .A2(n8245), .B1(n33453), .B2(n8237), .ZN(
        n33326) );
  NAND4_X1 U4672 ( .A1(n33329), .A2(n33328), .A3(n33327), .A4(n33326), .ZN(
        n33335) );
  AOI22_X1 U4673 ( .A1(n33460), .A2(n8235), .B1(n33459), .B2(n8264), .ZN(
        n33333) );
  AOI22_X1 U4674 ( .A1(n32711), .A2(n8263), .B1(n32710), .B2(n8249), .ZN(
        n33332) );
  AOI22_X1 U4675 ( .A1(n32713), .A2(n8253), .B1(n32712), .B2(n8239), .ZN(
        n33331) );
  AOI22_X1 U4676 ( .A1(n33466), .A2(n8261), .B1(n33465), .B2(n8255), .ZN(
        n33330) );
  NAND4_X1 U4677 ( .A1(n33333), .A2(n33332), .A3(n33331), .A4(n33330), .ZN(
        n33334) );
  NOR4_X1 U4678 ( .A1(n33337), .A2(n33336), .A3(n33335), .A4(n33334), .ZN(
        n33338) );
  OAI22_X1 U4679 ( .A1(n33338), .A2(n33476), .B1(n33475), .B2(n14150), .ZN(
        n5803) );
  AOI22_X1 U4680 ( .A1(n32685), .A2(n8288), .B1(n33423), .B2(n8280), .ZN(
        n33342) );
  AOI22_X1 U4681 ( .A1(n33426), .A2(n8294), .B1(n33425), .B2(n8284), .ZN(
        n33341) );
  AOI22_X1 U4682 ( .A1(n32689), .A2(n8290), .B1(n33427), .B2(n8289), .ZN(
        n33340) );
  AOI22_X1 U4683 ( .A1(n32691), .A2(n8283), .B1(n33429), .B2(n8286), .ZN(
        n33339) );
  NAND4_X1 U4684 ( .A1(n33342), .A2(n33341), .A3(n33340), .A4(n33339), .ZN(
        n33358) );
  AOI22_X1 U4685 ( .A1(n33436), .A2(n8268), .B1(n33435), .B2(n8274), .ZN(
        n33346) );
  AOI22_X1 U4686 ( .A1(n33438), .A2(n8276), .B1(n33437), .B2(n8272), .ZN(
        n33345) );
  AOI22_X1 U4687 ( .A1(n33440), .A2(n8266), .B1(n33439), .B2(n8273), .ZN(
        n33344) );
  AOI22_X1 U4688 ( .A1(n32699), .A2(n8278), .B1(n33441), .B2(n8270), .ZN(
        n33343) );
  NAND4_X1 U4689 ( .A1(n33346), .A2(n33345), .A3(n33344), .A4(n33343), .ZN(
        n33357) );
  AOI22_X1 U4690 ( .A1(n33448), .A2(n8275), .B1(n33447), .B2(n8292), .ZN(
        n33350) );
  AOI22_X1 U4691 ( .A1(n32703), .A2(n8282), .B1(n33449), .B2(n8279), .ZN(
        n33349) );
  AOI22_X1 U4692 ( .A1(n33452), .A2(n8265), .B1(n33451), .B2(n8291), .ZN(
        n33348) );
  AOI22_X1 U4693 ( .A1(n32707), .A2(n8277), .B1(n33453), .B2(n8269), .ZN(
        n33347) );
  NAND4_X1 U4694 ( .A1(n33350), .A2(n33349), .A3(n33348), .A4(n33347), .ZN(
        n33356) );
  AOI22_X1 U4695 ( .A1(n33460), .A2(n8267), .B1(n33459), .B2(n8296), .ZN(
        n33354) );
  AOI22_X1 U4696 ( .A1(n33462), .A2(n8295), .B1(n33461), .B2(n8281), .ZN(
        n33353) );
  AOI22_X1 U4697 ( .A1(n33464), .A2(n8285), .B1(n33463), .B2(n8271), .ZN(
        n33352) );
  AOI22_X1 U4698 ( .A1(n32715), .A2(n8293), .B1(n33465), .B2(n8287), .ZN(
        n33351) );
  NAND4_X1 U4699 ( .A1(n33354), .A2(n33353), .A3(n33352), .A4(n33351), .ZN(
        n33355) );
  NOR4_X1 U4700 ( .A1(n33358), .A2(n33357), .A3(n33356), .A4(n33355), .ZN(
        n33359) );
  OAI22_X1 U4701 ( .A1(n33359), .A2(n33476), .B1(n33475), .B2(n14151), .ZN(
        n5804) );
  AOI22_X1 U4702 ( .A1(n33424), .A2(n8320), .B1(n32684), .B2(n8312), .ZN(
        n33363) );
  AOI22_X1 U4703 ( .A1(n32687), .A2(n8326), .B1(n32686), .B2(n8316), .ZN(
        n33362) );
  AOI22_X1 U4704 ( .A1(n32689), .A2(n8322), .B1(n32688), .B2(n8321), .ZN(
        n33361) );
  AOI22_X1 U4705 ( .A1(n32691), .A2(n8315), .B1(n32690), .B2(n8318), .ZN(
        n33360) );
  NAND4_X1 U4706 ( .A1(n33363), .A2(n33362), .A3(n33361), .A4(n33360), .ZN(
        n33379) );
  AOI22_X1 U4707 ( .A1(n33436), .A2(n8300), .B1(n32692), .B2(n8306), .ZN(
        n33367) );
  AOI22_X1 U4708 ( .A1(n33438), .A2(n8308), .B1(n32694), .B2(n8304), .ZN(
        n33366) );
  AOI22_X1 U4709 ( .A1(n33440), .A2(n8298), .B1(n32696), .B2(n8305), .ZN(
        n33365) );
  AOI22_X1 U4710 ( .A1(n33442), .A2(n8310), .B1(n32698), .B2(n8302), .ZN(
        n33364) );
  NAND4_X1 U4711 ( .A1(n33367), .A2(n33366), .A3(n33365), .A4(n33364), .ZN(
        n33378) );
  AOI22_X1 U4712 ( .A1(n33448), .A2(n8307), .B1(n32700), .B2(n8324), .ZN(
        n33371) );
  AOI22_X1 U4713 ( .A1(n33450), .A2(n8314), .B1(n32702), .B2(n8311), .ZN(
        n33370) );
  AOI22_X1 U4714 ( .A1(n32705), .A2(n8297), .B1(n32704), .B2(n8323), .ZN(
        n33369) );
  AOI22_X1 U4715 ( .A1(n33454), .A2(n8309), .B1(n32706), .B2(n8301), .ZN(
        n33368) );
  NAND4_X1 U4716 ( .A1(n33371), .A2(n33370), .A3(n33369), .A4(n33368), .ZN(
        n33377) );
  AOI22_X1 U4717 ( .A1(n32709), .A2(n8299), .B1(n32708), .B2(n8328), .ZN(
        n33375) );
  AOI22_X1 U4718 ( .A1(n33462), .A2(n8327), .B1(n32710), .B2(n8313), .ZN(
        n33374) );
  AOI22_X1 U4719 ( .A1(n33464), .A2(n8317), .B1(n32712), .B2(n8303), .ZN(
        n33373) );
  AOI22_X1 U4720 ( .A1(n33466), .A2(n8325), .B1(n32714), .B2(n8319), .ZN(
        n33372) );
  NAND4_X1 U4721 ( .A1(n33375), .A2(n33374), .A3(n33373), .A4(n33372), .ZN(
        n33376) );
  NOR4_X1 U4722 ( .A1(n33379), .A2(n33378), .A3(n33377), .A4(n33376), .ZN(
        n33380) );
  OAI22_X1 U4723 ( .A1(n33380), .A2(n33476), .B1(n33475), .B2(n14152), .ZN(
        n5805) );
  AOI22_X1 U4724 ( .A1(n33424), .A2(n8352), .B1(n32684), .B2(n8344), .ZN(
        n33384) );
  AOI22_X1 U4725 ( .A1(n33426), .A2(n8358), .B1(n32686), .B2(n8348), .ZN(
        n33383) );
  AOI22_X1 U4726 ( .A1(n33428), .A2(n8354), .B1(n32688), .B2(n8353), .ZN(
        n33382) );
  AOI22_X1 U4727 ( .A1(n33430), .A2(n8347), .B1(n32690), .B2(n8350), .ZN(
        n33381) );
  NAND4_X1 U4728 ( .A1(n33384), .A2(n33383), .A3(n33382), .A4(n33381), .ZN(
        n33400) );
  AOI22_X1 U4729 ( .A1(n32693), .A2(n8332), .B1(n33435), .B2(n8338), .ZN(
        n33388) );
  AOI22_X1 U4730 ( .A1(n32695), .A2(n8340), .B1(n33437), .B2(n8336), .ZN(
        n33387) );
  AOI22_X1 U4731 ( .A1(n32697), .A2(n8330), .B1(n33439), .B2(n8337), .ZN(
        n33386) );
  AOI22_X1 U4732 ( .A1(n32699), .A2(n8342), .B1(n32698), .B2(n8334), .ZN(
        n33385) );
  NAND4_X1 U4733 ( .A1(n33388), .A2(n33387), .A3(n33386), .A4(n33385), .ZN(
        n33399) );
  AOI22_X1 U4734 ( .A1(n32701), .A2(n8339), .B1(n33447), .B2(n8356), .ZN(
        n33392) );
  AOI22_X1 U4735 ( .A1(n33450), .A2(n8346), .B1(n33449), .B2(n8343), .ZN(
        n33391) );
  AOI22_X1 U4736 ( .A1(n33452), .A2(n8329), .B1(n33451), .B2(n8355), .ZN(
        n33390) );
  AOI22_X1 U4737 ( .A1(n33454), .A2(n8341), .B1(n33453), .B2(n8333), .ZN(
        n33389) );
  NAND4_X1 U4738 ( .A1(n33392), .A2(n33391), .A3(n33390), .A4(n33389), .ZN(
        n33398) );
  AOI22_X1 U4739 ( .A1(n32709), .A2(n8331), .B1(n33459), .B2(n8360), .ZN(
        n33396) );
  AOI22_X1 U4740 ( .A1(n33462), .A2(n8359), .B1(n33461), .B2(n8345), .ZN(
        n33395) );
  AOI22_X1 U4741 ( .A1(n32713), .A2(n8349), .B1(n33463), .B2(n8335), .ZN(
        n33394) );
  AOI22_X1 U4742 ( .A1(n33466), .A2(n8357), .B1(n33465), .B2(n8351), .ZN(
        n33393) );
  NAND4_X1 U4743 ( .A1(n33396), .A2(n33395), .A3(n33394), .A4(n33393), .ZN(
        n33397) );
  NOR4_X1 U4744 ( .A1(n33400), .A2(n33399), .A3(n33398), .A4(n33397), .ZN(
        n33401) );
  OAI22_X1 U4745 ( .A1(n33401), .A2(n33476), .B1(n33475), .B2(n14153), .ZN(
        n5806) );
  AOI22_X1 U4746 ( .A1(n32685), .A2(n8384), .B1(n33423), .B2(n8376), .ZN(
        n33405) );
  AOI22_X1 U4747 ( .A1(n32687), .A2(n8390), .B1(n33425), .B2(n8380), .ZN(
        n33404) );
  AOI22_X1 U4748 ( .A1(n33428), .A2(n8386), .B1(n33427), .B2(n8385), .ZN(
        n33403) );
  AOI22_X1 U4749 ( .A1(n33430), .A2(n8379), .B1(n33429), .B2(n8382), .ZN(
        n33402) );
  NAND4_X1 U4750 ( .A1(n33405), .A2(n33404), .A3(n33403), .A4(n33402), .ZN(
        n33421) );
  AOI22_X1 U4751 ( .A1(n32693), .A2(n8364), .B1(n33435), .B2(n8370), .ZN(
        n33409) );
  AOI22_X1 U4752 ( .A1(n32695), .A2(n8372), .B1(n33437), .B2(n8368), .ZN(
        n33408) );
  AOI22_X1 U4753 ( .A1(n33440), .A2(n8362), .B1(n33439), .B2(n8369), .ZN(
        n33407) );
  AOI22_X1 U4754 ( .A1(n33442), .A2(n8374), .B1(n33441), .B2(n8366), .ZN(
        n33406) );
  NAND4_X1 U4755 ( .A1(n33409), .A2(n33408), .A3(n33407), .A4(n33406), .ZN(
        n33420) );
  AOI22_X1 U4756 ( .A1(n33448), .A2(n8371), .B1(n33447), .B2(n8388), .ZN(
        n33413) );
  AOI22_X1 U4757 ( .A1(n33450), .A2(n8378), .B1(n33449), .B2(n8375), .ZN(
        n33412) );
  AOI22_X1 U4758 ( .A1(n32705), .A2(n8361), .B1(n33451), .B2(n8387), .ZN(
        n33411) );
  AOI22_X1 U4759 ( .A1(n32707), .A2(n8373), .B1(n33453), .B2(n8365), .ZN(
        n33410) );
  NAND4_X1 U4760 ( .A1(n33413), .A2(n33412), .A3(n33411), .A4(n33410), .ZN(
        n33419) );
  AOI22_X1 U4761 ( .A1(n33460), .A2(n8363), .B1(n33459), .B2(n8392), .ZN(
        n33417) );
  AOI22_X1 U4762 ( .A1(n33462), .A2(n8391), .B1(n33461), .B2(n8377), .ZN(
        n33416) );
  AOI22_X1 U4763 ( .A1(n33464), .A2(n8381), .B1(n33463), .B2(n8367), .ZN(
        n33415) );
  AOI22_X1 U4764 ( .A1(n32715), .A2(n8389), .B1(n33465), .B2(n8383), .ZN(
        n33414) );
  NAND4_X1 U4765 ( .A1(n33417), .A2(n33416), .A3(n33415), .A4(n33414), .ZN(
        n33418) );
  NOR4_X1 U4766 ( .A1(n33421), .A2(n33420), .A3(n33419), .A4(n33418), .ZN(
        n33422) );
  OAI22_X1 U4767 ( .A1(n33422), .A2(n33476), .B1(n33475), .B2(n14154), .ZN(
        n5807) );
  AOI22_X1 U4768 ( .A1(n33424), .A2(n8416), .B1(n32684), .B2(n8408), .ZN(
        n33434) );
  AOI22_X1 U4769 ( .A1(n32687), .A2(n8422), .B1(n32686), .B2(n8412), .ZN(
        n33433) );
  AOI22_X1 U4770 ( .A1(n32689), .A2(n8418), .B1(n32688), .B2(n8417), .ZN(
        n33432) );
  AOI22_X1 U4771 ( .A1(n32691), .A2(n8411), .B1(n32690), .B2(n8414), .ZN(
        n33431) );
  NAND4_X1 U4772 ( .A1(n33434), .A2(n33433), .A3(n33432), .A4(n33431), .ZN(
        n33474) );
  AOI22_X1 U4773 ( .A1(n32693), .A2(n8396), .B1(n32692), .B2(n8402), .ZN(
        n33446) );
  AOI22_X1 U4774 ( .A1(n32695), .A2(n8404), .B1(n32694), .B2(n8400), .ZN(
        n33445) );
  AOI22_X1 U4775 ( .A1(n32697), .A2(n8394), .B1(n32696), .B2(n8401), .ZN(
        n33444) );
  AOI22_X1 U4776 ( .A1(n32699), .A2(n8406), .B1(n32698), .B2(n8398), .ZN(
        n33443) );
  NAND4_X1 U4777 ( .A1(n33446), .A2(n33445), .A3(n33444), .A4(n33443), .ZN(
        n33473) );
  AOI22_X1 U4778 ( .A1(n32701), .A2(n8403), .B1(n32700), .B2(n8420), .ZN(
        n33458) );
  AOI22_X1 U4779 ( .A1(n33450), .A2(n8410), .B1(n32702), .B2(n8407), .ZN(
        n33457) );
  AOI22_X1 U4780 ( .A1(n33452), .A2(n8393), .B1(n32704), .B2(n8419), .ZN(
        n33456) );
  AOI22_X1 U4781 ( .A1(n32707), .A2(n8405), .B1(n32706), .B2(n8397), .ZN(
        n33455) );
  NAND4_X1 U4782 ( .A1(n33458), .A2(n33457), .A3(n33456), .A4(n33455), .ZN(
        n33472) );
  AOI22_X1 U4783 ( .A1(n33460), .A2(n8395), .B1(n32708), .B2(n8424), .ZN(
        n33470) );
  AOI22_X1 U4784 ( .A1(n32711), .A2(n8423), .B1(n32710), .B2(n8409), .ZN(
        n33469) );
  AOI22_X1 U4785 ( .A1(n32713), .A2(n8413), .B1(n32712), .B2(n8399), .ZN(
        n33468) );
  AOI22_X1 U4786 ( .A1(n32715), .A2(n8421), .B1(n32714), .B2(n8415), .ZN(
        n33467) );
  NAND4_X1 U4787 ( .A1(n33470), .A2(n33469), .A3(n33468), .A4(n33467), .ZN(
        n33471) );
  NOR4_X1 U4788 ( .A1(n33474), .A2(n33473), .A3(n33472), .A4(n33471), .ZN(
        n33477) );
  OAI22_X1 U4789 ( .A1(n33477), .A2(n33476), .B1(n33475), .B2(n14155), .ZN(
        n5808) );
  INV_X1 U4790 ( .A(ADD_RD2[2]), .ZN(n33478) );
  INV_X1 U4791 ( .A(ADD_RD2[1]), .ZN(n33522) );
  NAND2_X1 U4792 ( .A1(n33478), .A2(n33522), .ZN(n33493) );
  NOR2_X1 U4793 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .ZN(n33479) );
  INV_X1 U4794 ( .A(ADD_RD2[4]), .ZN(n33484) );
  NAND2_X1 U4795 ( .A1(n33479), .A2(n33484), .ZN(n33502) );
  NAND3_X1 U4796 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n33484), .ZN(n33500)
         );
  NAND2_X1 U4797 ( .A1(ADD_RD2[2]), .A2(n33522), .ZN(n33506) );
  AOI22_X1 U4798 ( .A1(n7432), .A2(n34158), .B1(n7431), .B2(n32676), .ZN(
        n33483) );
  INV_X1 U4799 ( .A(ADD_RD2[3]), .ZN(n33491) );
  NAND3_X1 U4800 ( .A1(ADD_RD2[0]), .A2(n33484), .A3(n33491), .ZN(n33486) );
  NAND2_X1 U4801 ( .A1(ADD_RD2[1]), .A2(n33478), .ZN(n33498) );
  NAND2_X1 U4802 ( .A1(ADD_RD2[4]), .A2(n33479), .ZN(n33505) );
  AOI22_X1 U4803 ( .A1(n7430), .A2(n32678), .B1(n7429), .B2(n32675), .ZN(
        n33482) );
  NAND2_X1 U4804 ( .A1(ADD_RD2[2]), .A2(ADD_RD2[1]), .ZN(n33501) );
  NOR2_X1 U4805 ( .A1(n33486), .A2(n33501), .ZN(n34162) );
  NAND3_X1 U4806 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(ADD_RD2[3]), .ZN(
        n33492) );
  AOI22_X1 U4807 ( .A1(n7428), .A2(n32667), .B1(n7427), .B2(n34161), .ZN(
        n33481) );
  INV_X1 U4808 ( .A(ADD_RD2[0]), .ZN(n33485) );
  NAND3_X1 U4809 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .A3(n33485), .ZN(n33504)
         );
  AOI22_X1 U4810 ( .A1(n7426), .A2(n32677), .B1(n7425), .B2(n32674), .ZN(
        n33480) );
  NAND4_X1 U4811 ( .A1(n33483), .A2(n33482), .A3(n33481), .A4(n33480), .ZN(
        n33514) );
  NAND3_X1 U4812 ( .A1(ADD_RD2[3]), .A2(n33485), .A3(n33484), .ZN(n33499) );
  NOR2_X1 U4813 ( .A1(n33486), .A2(n33498), .ZN(n34169) );
  AOI22_X1 U4814 ( .A1(n7424), .A2(n34170), .B1(n7423), .B2(n32717), .ZN(
        n33490) );
  AOI22_X1 U4815 ( .A1(n7422), .A2(n32680), .B1(n7421), .B2(n32718), .ZN(
        n33489) );
  AOI22_X1 U4816 ( .A1(n7420), .A2(n32679), .B1(n7419), .B2(n32673), .ZN(
        n33488) );
  AOI22_X1 U4817 ( .A1(n7418), .A2(n32719), .B1(n7417), .B2(n32672), .ZN(
        n33487) );
  NAND4_X1 U4818 ( .A1(n33490), .A2(n33489), .A3(n33488), .A4(n33487), .ZN(
        n33513) );
  NAND3_X1 U4819 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[0]), .A3(n33491), .ZN(n33503)
         );
  AOI22_X1 U4820 ( .A1(n7416), .A2(n34182), .B1(n7415), .B2(n32671), .ZN(
        n33497) );
  AOI22_X1 U4821 ( .A1(n7414), .A2(n34184), .B1(n7413), .B2(n34183), .ZN(
        n33496) );
  NOR2_X1 U4822 ( .A1(n33501), .A2(n33504), .ZN(n34186) );
  AOI22_X1 U4823 ( .A1(n7412), .A2(n32666), .B1(n7411), .B2(n34185), .ZN(
        n33495) );
  AOI22_X1 U4824 ( .A1(n7410), .A2(n32682), .B1(n7409), .B2(n32670), .ZN(
        n33494) );
  NAND4_X1 U4825 ( .A1(n33497), .A2(n33496), .A3(n33495), .A4(n33494), .ZN(
        n33512) );
  NOR2_X1 U4826 ( .A1(n33500), .A2(n33498), .ZN(n34193) );
  AOI22_X1 U4827 ( .A1(n7408), .A2(n34194), .B1(n7407), .B2(n32720), .ZN(
        n33510) );
  AOI22_X1 U4828 ( .A1(n7406), .A2(n32681), .B1(n7405), .B2(n32669), .ZN(
        n33509) );
  AOI22_X1 U4829 ( .A1(n7404), .A2(n34198), .B1(n7403), .B2(n32668), .ZN(
        n33508) );
  AOI22_X1 U4830 ( .A1(n7402), .A2(n34200), .B1(n7401), .B2(n32721), .ZN(
        n33507) );
  NAND4_X1 U4831 ( .A1(n33510), .A2(n33509), .A3(n33508), .A4(n33507), .ZN(
        n33511) );
  NOR4_X1 U4832 ( .A1(n33514), .A2(n33513), .A3(n33512), .A4(n33511), .ZN(
        n33526) );
  OAI22_X1 U4833 ( .A1(n33517), .A2(ADD_RD2[4]), .B1(n33516), .B2(ADD_RD2[3]), 
        .ZN(n33515) );
  AOI221_X1 U4834 ( .B1(n33517), .B2(ADD_RD2[4]), .C1(ADD_RD2[3]), .C2(n33516), 
        .A(n33515), .ZN(n33525) );
  OAI22_X1 U4835 ( .A1(n33520), .A2(ADD_RD2[0]), .B1(n33519), .B2(ADD_RD2[2]), 
        .ZN(n33518) );
  AOI221_X1 U4836 ( .B1(n33520), .B2(ADD_RD2[0]), .C1(ADD_RD2[2]), .C2(n33519), 
        .A(n33518), .ZN(n33524) );
  AOI22_X1 U4837 ( .A1(ADD_WR[1]), .A2(n33522), .B1(ADD_RD2[1]), .B2(n33521), 
        .ZN(n33523) );
  NAND4_X1 U4838 ( .A1(WR), .A2(n33525), .A3(n33524), .A4(n33523), .ZN(n34209)
         );
  OAI22_X1 U4839 ( .A1(n33526), .A2(n32665), .B1(n34213), .B2(n32722), .ZN(
        n5812) );
  AOI22_X1 U4840 ( .A1(n7464), .A2(n34158), .B1(n7463), .B2(n32676), .ZN(
        n33530) );
  AOI22_X1 U4841 ( .A1(n7462), .A2(n32678), .B1(n7461), .B2(n32675), .ZN(
        n33529) );
  AOI22_X1 U4842 ( .A1(n7460), .A2(n32667), .B1(n7459), .B2(n34161), .ZN(
        n33528) );
  AOI22_X1 U4843 ( .A1(n7458), .A2(n32677), .B1(n7457), .B2(n32674), .ZN(
        n33527) );
  NAND4_X1 U4844 ( .A1(n33530), .A2(n33529), .A3(n33528), .A4(n33527), .ZN(
        n33546) );
  AOI22_X1 U4845 ( .A1(n7456), .A2(n34170), .B1(n7455), .B2(n32717), .ZN(
        n33534) );
  AOI22_X1 U4846 ( .A1(n7454), .A2(n32680), .B1(n7453), .B2(n32718), .ZN(
        n33533) );
  AOI22_X1 U4847 ( .A1(n7452), .A2(n32679), .B1(n7451), .B2(n32673), .ZN(
        n33532) );
  AOI22_X1 U4848 ( .A1(n7450), .A2(n32719), .B1(n7449), .B2(n32672), .ZN(
        n33531) );
  NAND4_X1 U4849 ( .A1(n33534), .A2(n33533), .A3(n33532), .A4(n33531), .ZN(
        n33545) );
  AOI22_X1 U4850 ( .A1(n7448), .A2(n34182), .B1(n7447), .B2(n32671), .ZN(
        n33538) );
  AOI22_X1 U4851 ( .A1(n7446), .A2(n34184), .B1(n7445), .B2(n34183), .ZN(
        n33537) );
  AOI22_X1 U4852 ( .A1(n7444), .A2(n32666), .B1(n7443), .B2(n34185), .ZN(
        n33536) );
  AOI22_X1 U4853 ( .A1(n7442), .A2(n32682), .B1(n7441), .B2(n32670), .ZN(
        n33535) );
  NAND4_X1 U4854 ( .A1(n33538), .A2(n33537), .A3(n33536), .A4(n33535), .ZN(
        n33544) );
  AOI22_X1 U4855 ( .A1(n7440), .A2(n34194), .B1(n7439), .B2(n32720), .ZN(
        n33542) );
  AOI22_X1 U4856 ( .A1(n7438), .A2(n32681), .B1(n7437), .B2(n32669), .ZN(
        n33541) );
  AOI22_X1 U4857 ( .A1(n7436), .A2(n34198), .B1(n7435), .B2(n32668), .ZN(
        n33540) );
  AOI22_X1 U4858 ( .A1(n7434), .A2(n34200), .B1(n7433), .B2(n32721), .ZN(
        n33539) );
  NAND4_X1 U4859 ( .A1(n33542), .A2(n33541), .A3(n33540), .A4(n33539), .ZN(
        n33543) );
  NOR4_X1 U4860 ( .A1(n33546), .A2(n33545), .A3(n33544), .A4(n33543), .ZN(
        n33547) );
  OAI22_X1 U4861 ( .A1(n33547), .A2(n32665), .B1(n34214), .B2(n32722), .ZN(
        n5813) );
  AOI22_X1 U4862 ( .A1(n7496), .A2(n34158), .B1(n7495), .B2(n32676), .ZN(
        n33551) );
  AOI22_X1 U4863 ( .A1(n7494), .A2(n32678), .B1(n7493), .B2(n32675), .ZN(
        n33550) );
  AOI22_X1 U4864 ( .A1(n7492), .A2(n32667), .B1(n7491), .B2(n34161), .ZN(
        n33549) );
  AOI22_X1 U4865 ( .A1(n7490), .A2(n32677), .B1(n7489), .B2(n32674), .ZN(
        n33548) );
  NAND4_X1 U4866 ( .A1(n33551), .A2(n33550), .A3(n33549), .A4(n33548), .ZN(
        n33567) );
  AOI22_X1 U4867 ( .A1(n7488), .A2(n34170), .B1(n7487), .B2(n32717), .ZN(
        n33555) );
  AOI22_X1 U4868 ( .A1(n7486), .A2(n32680), .B1(n7485), .B2(n32718), .ZN(
        n33554) );
  AOI22_X1 U4869 ( .A1(n7484), .A2(n32679), .B1(n7483), .B2(n32673), .ZN(
        n33553) );
  AOI22_X1 U4870 ( .A1(n7482), .A2(n32719), .B1(n7481), .B2(n32672), .ZN(
        n33552) );
  NAND4_X1 U4871 ( .A1(n33555), .A2(n33554), .A3(n33553), .A4(n33552), .ZN(
        n33566) );
  AOI22_X1 U4872 ( .A1(n7480), .A2(n34182), .B1(n7479), .B2(n32671), .ZN(
        n33559) );
  AOI22_X1 U4873 ( .A1(n7478), .A2(n34184), .B1(n7477), .B2(n34183), .ZN(
        n33558) );
  AOI22_X1 U4874 ( .A1(n7476), .A2(n32666), .B1(n7475), .B2(n34185), .ZN(
        n33557) );
  AOI22_X1 U4875 ( .A1(n7474), .A2(n32682), .B1(n7473), .B2(n32670), .ZN(
        n33556) );
  NAND4_X1 U4876 ( .A1(n33559), .A2(n33558), .A3(n33557), .A4(n33556), .ZN(
        n33565) );
  AOI22_X1 U4877 ( .A1(n7472), .A2(n34194), .B1(n7471), .B2(n32720), .ZN(
        n33563) );
  AOI22_X1 U4878 ( .A1(n7470), .A2(n32681), .B1(n7469), .B2(n32669), .ZN(
        n33562) );
  AOI22_X1 U4879 ( .A1(n7468), .A2(n34198), .B1(n7467), .B2(n32668), .ZN(
        n33561) );
  AOI22_X1 U4880 ( .A1(n7466), .A2(n34200), .B1(n7465), .B2(n34199), .ZN(
        n33560) );
  NAND4_X1 U4881 ( .A1(n33563), .A2(n33562), .A3(n33561), .A4(n33560), .ZN(
        n33564) );
  NOR4_X1 U4882 ( .A1(n33567), .A2(n33566), .A3(n33565), .A4(n33564), .ZN(
        n33568) );
  OAI22_X1 U4883 ( .A1(n33568), .A2(n32665), .B1(n34215), .B2(n32722), .ZN(
        n5814) );
  AOI22_X1 U4884 ( .A1(n7528), .A2(n34158), .B1(n7527), .B2(n32676), .ZN(
        n33572) );
  AOI22_X1 U4885 ( .A1(n7526), .A2(n32678), .B1(n7525), .B2(n32675), .ZN(
        n33571) );
  AOI22_X1 U4886 ( .A1(n7524), .A2(n32667), .B1(n7523), .B2(n34161), .ZN(
        n33570) );
  AOI22_X1 U4887 ( .A1(n7522), .A2(n32677), .B1(n7521), .B2(n32674), .ZN(
        n33569) );
  NAND4_X1 U4888 ( .A1(n33572), .A2(n33571), .A3(n33570), .A4(n33569), .ZN(
        n33588) );
  AOI22_X1 U4889 ( .A1(n7520), .A2(n34170), .B1(n7519), .B2(n32717), .ZN(
        n33576) );
  AOI22_X1 U4890 ( .A1(n7518), .A2(n32680), .B1(n7517), .B2(n32718), .ZN(
        n33575) );
  AOI22_X1 U4891 ( .A1(n7516), .A2(n32679), .B1(n7515), .B2(n32673), .ZN(
        n33574) );
  AOI22_X1 U4892 ( .A1(n7514), .A2(n34176), .B1(n7513), .B2(n32672), .ZN(
        n33573) );
  NAND4_X1 U4893 ( .A1(n33576), .A2(n33575), .A3(n33574), .A4(n33573), .ZN(
        n33587) );
  AOI22_X1 U4894 ( .A1(n7512), .A2(n34182), .B1(n7511), .B2(n32671), .ZN(
        n33580) );
  AOI22_X1 U4895 ( .A1(n7510), .A2(n34184), .B1(n7509), .B2(n34183), .ZN(
        n33579) );
  AOI22_X1 U4896 ( .A1(n7508), .A2(n32666), .B1(n7507), .B2(n34185), .ZN(
        n33578) );
  AOI22_X1 U4897 ( .A1(n7506), .A2(n32682), .B1(n7505), .B2(n32670), .ZN(
        n33577) );
  NAND4_X1 U4898 ( .A1(n33580), .A2(n33579), .A3(n33578), .A4(n33577), .ZN(
        n33586) );
  AOI22_X1 U4899 ( .A1(n7504), .A2(n34194), .B1(n7503), .B2(n32720), .ZN(
        n33584) );
  AOI22_X1 U4900 ( .A1(n7502), .A2(n32681), .B1(n7501), .B2(n32669), .ZN(
        n33583) );
  AOI22_X1 U4901 ( .A1(n7500), .A2(n34198), .B1(n7499), .B2(n32668), .ZN(
        n33582) );
  AOI22_X1 U4902 ( .A1(n7498), .A2(n34200), .B1(n7497), .B2(n34199), .ZN(
        n33581) );
  NAND4_X1 U4903 ( .A1(n33584), .A2(n33583), .A3(n33582), .A4(n33581), .ZN(
        n33585) );
  NOR4_X1 U4904 ( .A1(n33588), .A2(n33587), .A3(n33586), .A4(n33585), .ZN(
        n33589) );
  OAI22_X1 U4905 ( .A1(n33589), .A2(n32665), .B1(n34216), .B2(n32722), .ZN(
        n5815) );
  AOI22_X1 U4906 ( .A1(n7560), .A2(n34158), .B1(n7559), .B2(n32676), .ZN(
        n33593) );
  AOI22_X1 U4907 ( .A1(n7558), .A2(n32678), .B1(n7557), .B2(n32675), .ZN(
        n33592) );
  AOI22_X1 U4908 ( .A1(n7556), .A2(n32667), .B1(n7555), .B2(n34161), .ZN(
        n33591) );
  AOI22_X1 U4909 ( .A1(n7554), .A2(n32677), .B1(n7553), .B2(n32674), .ZN(
        n33590) );
  NAND4_X1 U4910 ( .A1(n33593), .A2(n33592), .A3(n33591), .A4(n33590), .ZN(
        n33609) );
  AOI22_X1 U4911 ( .A1(n7552), .A2(n34170), .B1(n7551), .B2(n32717), .ZN(
        n33597) );
  AOI22_X1 U4912 ( .A1(n7550), .A2(n32680), .B1(n7549), .B2(n32718), .ZN(
        n33596) );
  AOI22_X1 U4913 ( .A1(n7548), .A2(n32679), .B1(n7547), .B2(n32673), .ZN(
        n33595) );
  AOI22_X1 U4914 ( .A1(n7546), .A2(n34176), .B1(n7545), .B2(n32672), .ZN(
        n33594) );
  NAND4_X1 U4915 ( .A1(n33597), .A2(n33596), .A3(n33595), .A4(n33594), .ZN(
        n33608) );
  AOI22_X1 U4916 ( .A1(n7544), .A2(n34182), .B1(n7543), .B2(n32671), .ZN(
        n33601) );
  AOI22_X1 U4917 ( .A1(n7542), .A2(n34184), .B1(n7541), .B2(n34183), .ZN(
        n33600) );
  AOI22_X1 U4918 ( .A1(n7540), .A2(n32666), .B1(n7539), .B2(n34185), .ZN(
        n33599) );
  AOI22_X1 U4919 ( .A1(n7538), .A2(n32682), .B1(n7537), .B2(n32670), .ZN(
        n33598) );
  NAND4_X1 U4920 ( .A1(n33601), .A2(n33600), .A3(n33599), .A4(n33598), .ZN(
        n33607) );
  AOI22_X1 U4921 ( .A1(n7536), .A2(n34194), .B1(n7535), .B2(n32720), .ZN(
        n33605) );
  AOI22_X1 U4922 ( .A1(n7534), .A2(n32681), .B1(n7533), .B2(n32669), .ZN(
        n33604) );
  AOI22_X1 U4923 ( .A1(n7532), .A2(n34198), .B1(n7531), .B2(n32668), .ZN(
        n33603) );
  AOI22_X1 U4924 ( .A1(n7530), .A2(n34200), .B1(n7529), .B2(n32721), .ZN(
        n33602) );
  NAND4_X1 U4925 ( .A1(n33605), .A2(n33604), .A3(n33603), .A4(n33602), .ZN(
        n33606) );
  NOR4_X1 U4926 ( .A1(n33609), .A2(n33608), .A3(n33607), .A4(n33606), .ZN(
        n33610) );
  OAI22_X1 U4927 ( .A1(n33610), .A2(n32665), .B1(n32723), .B2(n32722), .ZN(
        n5816) );
  AOI22_X1 U4928 ( .A1(n7592), .A2(n34158), .B1(n7591), .B2(n32676), .ZN(
        n33614) );
  AOI22_X1 U4929 ( .A1(n7590), .A2(n32678), .B1(n7589), .B2(n32675), .ZN(
        n33613) );
  AOI22_X1 U4930 ( .A1(n7588), .A2(n32667), .B1(n7587), .B2(n34161), .ZN(
        n33612) );
  AOI22_X1 U4931 ( .A1(n7586), .A2(n32677), .B1(n7585), .B2(n32674), .ZN(
        n33611) );
  NAND4_X1 U4932 ( .A1(n33614), .A2(n33613), .A3(n33612), .A4(n33611), .ZN(
        n33630) );
  AOI22_X1 U4933 ( .A1(n7584), .A2(n34170), .B1(n7583), .B2(n32717), .ZN(
        n33618) );
  AOI22_X1 U4934 ( .A1(n7582), .A2(n32680), .B1(n7581), .B2(n32718), .ZN(
        n33617) );
  AOI22_X1 U4935 ( .A1(n7580), .A2(n32679), .B1(n7579), .B2(n32673), .ZN(
        n33616) );
  AOI22_X1 U4936 ( .A1(n7578), .A2(n34176), .B1(n7577), .B2(n32672), .ZN(
        n33615) );
  NAND4_X1 U4937 ( .A1(n33618), .A2(n33617), .A3(n33616), .A4(n33615), .ZN(
        n33629) );
  AOI22_X1 U4938 ( .A1(n7576), .A2(n34182), .B1(n7575), .B2(n32671), .ZN(
        n33622) );
  AOI22_X1 U4939 ( .A1(n7574), .A2(n34184), .B1(n7573), .B2(n34183), .ZN(
        n33621) );
  AOI22_X1 U4940 ( .A1(n7572), .A2(n32666), .B1(n7571), .B2(n34185), .ZN(
        n33620) );
  AOI22_X1 U4941 ( .A1(n7570), .A2(n32682), .B1(n7569), .B2(n32670), .ZN(
        n33619) );
  NAND4_X1 U4942 ( .A1(n33622), .A2(n33621), .A3(n33620), .A4(n33619), .ZN(
        n33628) );
  AOI22_X1 U4943 ( .A1(n7568), .A2(n34194), .B1(n7567), .B2(n32720), .ZN(
        n33626) );
  AOI22_X1 U4944 ( .A1(n7566), .A2(n32681), .B1(n7565), .B2(n32669), .ZN(
        n33625) );
  AOI22_X1 U4945 ( .A1(n7564), .A2(n34198), .B1(n7563), .B2(n32668), .ZN(
        n33624) );
  AOI22_X1 U4946 ( .A1(n7562), .A2(n34200), .B1(n7561), .B2(n34199), .ZN(
        n33623) );
  NAND4_X1 U4947 ( .A1(n33626), .A2(n33625), .A3(n33624), .A4(n33623), .ZN(
        n33627) );
  NOR4_X1 U4948 ( .A1(n33630), .A2(n33629), .A3(n33628), .A4(n33627), .ZN(
        n33631) );
  OAI22_X1 U4949 ( .A1(n33631), .A2(n32665), .B1(n20327), .B2(n32722), .ZN(
        n5817) );
  AOI22_X1 U4950 ( .A1(n7624), .A2(n34158), .B1(n7623), .B2(n32676), .ZN(
        n33635) );
  AOI22_X1 U4951 ( .A1(n7622), .A2(n32678), .B1(n7621), .B2(n32675), .ZN(
        n33634) );
  AOI22_X1 U4952 ( .A1(n7620), .A2(n32667), .B1(n7619), .B2(n34161), .ZN(
        n33633) );
  AOI22_X1 U4953 ( .A1(n7618), .A2(n32677), .B1(n7617), .B2(n32674), .ZN(
        n33632) );
  NAND4_X1 U4954 ( .A1(n33635), .A2(n33634), .A3(n33633), .A4(n33632), .ZN(
        n33651) );
  AOI22_X1 U4955 ( .A1(n7616), .A2(n34170), .B1(n7615), .B2(n34169), .ZN(
        n33639) );
  AOI22_X1 U4956 ( .A1(n7614), .A2(n32680), .B1(n7613), .B2(n34171), .ZN(
        n33638) );
  AOI22_X1 U4957 ( .A1(n7612), .A2(n32679), .B1(n7611), .B2(n32673), .ZN(
        n33637) );
  AOI22_X1 U4958 ( .A1(n7610), .A2(n34176), .B1(n7609), .B2(n32672), .ZN(
        n33636) );
  NAND4_X1 U4959 ( .A1(n33639), .A2(n33638), .A3(n33637), .A4(n33636), .ZN(
        n33650) );
  AOI22_X1 U4960 ( .A1(n7608), .A2(n34182), .B1(n7607), .B2(n32671), .ZN(
        n33643) );
  AOI22_X1 U4961 ( .A1(n7606), .A2(n34184), .B1(n7605), .B2(n34183), .ZN(
        n33642) );
  AOI22_X1 U4962 ( .A1(n7604), .A2(n32666), .B1(n7603), .B2(n34185), .ZN(
        n33641) );
  AOI22_X1 U4963 ( .A1(n7602), .A2(n32682), .B1(n7601), .B2(n32670), .ZN(
        n33640) );
  NAND4_X1 U4964 ( .A1(n33643), .A2(n33642), .A3(n33641), .A4(n33640), .ZN(
        n33649) );
  AOI22_X1 U4965 ( .A1(n7600), .A2(n34194), .B1(n7599), .B2(n34193), .ZN(
        n33647) );
  AOI22_X1 U4966 ( .A1(n7598), .A2(n32681), .B1(n7597), .B2(n32669), .ZN(
        n33646) );
  AOI22_X1 U4967 ( .A1(n7596), .A2(n34198), .B1(n7595), .B2(n32668), .ZN(
        n33645) );
  AOI22_X1 U4968 ( .A1(n7594), .A2(n34200), .B1(n7593), .B2(n34199), .ZN(
        n33644) );
  NAND4_X1 U4969 ( .A1(n33647), .A2(n33646), .A3(n33645), .A4(n33644), .ZN(
        n33648) );
  NOR4_X1 U4970 ( .A1(n33651), .A2(n33650), .A3(n33649), .A4(n33648), .ZN(
        n33652) );
  OAI22_X1 U4971 ( .A1(n33652), .A2(n32665), .B1(n14130), .B2(n32722), .ZN(
        n5818) );
  AOI22_X1 U4972 ( .A1(n7656), .A2(n34158), .B1(n7655), .B2(n32676), .ZN(
        n33656) );
  AOI22_X1 U4973 ( .A1(n7654), .A2(n32678), .B1(n7653), .B2(n32675), .ZN(
        n33655) );
  AOI22_X1 U4974 ( .A1(n7652), .A2(n32667), .B1(n7651), .B2(n34161), .ZN(
        n33654) );
  AOI22_X1 U4975 ( .A1(n7650), .A2(n32677), .B1(n7649), .B2(n32674), .ZN(
        n33653) );
  NAND4_X1 U4976 ( .A1(n33656), .A2(n33655), .A3(n33654), .A4(n33653), .ZN(
        n33672) );
  AOI22_X1 U4977 ( .A1(n7648), .A2(n34170), .B1(n7647), .B2(n34169), .ZN(
        n33660) );
  AOI22_X1 U4978 ( .A1(n7646), .A2(n32680), .B1(n7645), .B2(n34171), .ZN(
        n33659) );
  AOI22_X1 U4979 ( .A1(n7644), .A2(n32679), .B1(n7643), .B2(n32673), .ZN(
        n33658) );
  AOI22_X1 U4980 ( .A1(n7642), .A2(n34176), .B1(n7641), .B2(n32672), .ZN(
        n33657) );
  NAND4_X1 U4981 ( .A1(n33660), .A2(n33659), .A3(n33658), .A4(n33657), .ZN(
        n33671) );
  AOI22_X1 U4982 ( .A1(n7640), .A2(n34182), .B1(n7639), .B2(n32671), .ZN(
        n33664) );
  AOI22_X1 U4983 ( .A1(n7638), .A2(n34184), .B1(n7637), .B2(n34183), .ZN(
        n33663) );
  AOI22_X1 U4984 ( .A1(n7636), .A2(n32666), .B1(n7635), .B2(n34185), .ZN(
        n33662) );
  AOI22_X1 U4985 ( .A1(n7634), .A2(n32682), .B1(n7633), .B2(n32670), .ZN(
        n33661) );
  NAND4_X1 U4986 ( .A1(n33664), .A2(n33663), .A3(n33662), .A4(n33661), .ZN(
        n33670) );
  AOI22_X1 U4987 ( .A1(n7632), .A2(n34194), .B1(n7631), .B2(n34193), .ZN(
        n33668) );
  AOI22_X1 U4988 ( .A1(n7630), .A2(n32681), .B1(n7629), .B2(n32669), .ZN(
        n33667) );
  AOI22_X1 U4989 ( .A1(n7628), .A2(n34198), .B1(n7627), .B2(n32668), .ZN(
        n33666) );
  AOI22_X1 U4990 ( .A1(n7626), .A2(n34200), .B1(n7625), .B2(n34199), .ZN(
        n33665) );
  NAND4_X1 U4991 ( .A1(n33668), .A2(n33667), .A3(n33666), .A4(n33665), .ZN(
        n33669) );
  NOR4_X1 U4992 ( .A1(n33672), .A2(n33671), .A3(n33670), .A4(n33669), .ZN(
        n33673) );
  OAI22_X1 U4993 ( .A1(n33673), .A2(n32665), .B1(n14131), .B2(n32722), .ZN(
        n5819) );
  AOI22_X1 U4994 ( .A1(n7688), .A2(n32716), .B1(n7687), .B2(n32676), .ZN(
        n33677) );
  AOI22_X1 U4995 ( .A1(n7686), .A2(n32678), .B1(n7685), .B2(n32675), .ZN(
        n33676) );
  AOI22_X1 U4996 ( .A1(n7684), .A2(n32667), .B1(n7683), .B2(n34161), .ZN(
        n33675) );
  AOI22_X1 U4997 ( .A1(n7682), .A2(n32677), .B1(n7681), .B2(n32674), .ZN(
        n33674) );
  NAND4_X1 U4998 ( .A1(n33677), .A2(n33676), .A3(n33675), .A4(n33674), .ZN(
        n33693) );
  AOI22_X1 U4999 ( .A1(n7680), .A2(n34170), .B1(n7679), .B2(n34169), .ZN(
        n33681) );
  AOI22_X1 U5000 ( .A1(n7678), .A2(n32680), .B1(n7677), .B2(n34171), .ZN(
        n33680) );
  AOI22_X1 U5001 ( .A1(n7676), .A2(n32679), .B1(n7675), .B2(n32673), .ZN(
        n33679) );
  AOI22_X1 U5002 ( .A1(n7674), .A2(n34176), .B1(n7673), .B2(n32672), .ZN(
        n33678) );
  NAND4_X1 U5003 ( .A1(n33681), .A2(n33680), .A3(n33679), .A4(n33678), .ZN(
        n33692) );
  AOI22_X1 U5004 ( .A1(n7672), .A2(n34182), .B1(n7671), .B2(n32671), .ZN(
        n33685) );
  AOI22_X1 U5005 ( .A1(n7670), .A2(n34184), .B1(n7669), .B2(n34183), .ZN(
        n33684) );
  AOI22_X1 U5006 ( .A1(n7668), .A2(n32666), .B1(n7667), .B2(n34185), .ZN(
        n33683) );
  AOI22_X1 U5007 ( .A1(n7666), .A2(n32682), .B1(n7665), .B2(n32670), .ZN(
        n33682) );
  NAND4_X1 U5008 ( .A1(n33685), .A2(n33684), .A3(n33683), .A4(n33682), .ZN(
        n33691) );
  AOI22_X1 U5009 ( .A1(n7664), .A2(n34194), .B1(n7663), .B2(n34193), .ZN(
        n33689) );
  AOI22_X1 U5010 ( .A1(n7662), .A2(n32681), .B1(n7661), .B2(n32669), .ZN(
        n33688) );
  AOI22_X1 U5011 ( .A1(n7660), .A2(n34198), .B1(n7659), .B2(n32668), .ZN(
        n33687) );
  AOI22_X1 U5012 ( .A1(n7658), .A2(n34200), .B1(n7657), .B2(n32721), .ZN(
        n33686) );
  NAND4_X1 U5013 ( .A1(n33689), .A2(n33688), .A3(n33687), .A4(n33686), .ZN(
        n33690) );
  NOR4_X1 U5014 ( .A1(n33693), .A2(n33692), .A3(n33691), .A4(n33690), .ZN(
        n33694) );
  OAI22_X1 U5015 ( .A1(n33694), .A2(n32665), .B1(n14132), .B2(n32722), .ZN(
        n5820) );
  AOI22_X1 U5016 ( .A1(n7720), .A2(n32716), .B1(n7719), .B2(n32676), .ZN(
        n33698) );
  AOI22_X1 U5017 ( .A1(n7718), .A2(n32678), .B1(n7717), .B2(n32675), .ZN(
        n33697) );
  AOI22_X1 U5018 ( .A1(n7716), .A2(n32667), .B1(n7715), .B2(n34161), .ZN(
        n33696) );
  AOI22_X1 U5019 ( .A1(n7714), .A2(n32677), .B1(n7713), .B2(n32674), .ZN(
        n33695) );
  NAND4_X1 U5020 ( .A1(n33698), .A2(n33697), .A3(n33696), .A4(n33695), .ZN(
        n33714) );
  AOI22_X1 U5021 ( .A1(n7712), .A2(n34170), .B1(n7711), .B2(n34169), .ZN(
        n33702) );
  AOI22_X1 U5022 ( .A1(n7710), .A2(n32680), .B1(n7709), .B2(n34171), .ZN(
        n33701) );
  AOI22_X1 U5023 ( .A1(n7708), .A2(n32679), .B1(n7707), .B2(n32673), .ZN(
        n33700) );
  AOI22_X1 U5024 ( .A1(n7706), .A2(n32719), .B1(n7705), .B2(n32672), .ZN(
        n33699) );
  NAND4_X1 U5025 ( .A1(n33702), .A2(n33701), .A3(n33700), .A4(n33699), .ZN(
        n33713) );
  AOI22_X1 U5026 ( .A1(n7704), .A2(n34182), .B1(n7703), .B2(n32671), .ZN(
        n33706) );
  AOI22_X1 U5027 ( .A1(n7702), .A2(n34184), .B1(n7701), .B2(n34183), .ZN(
        n33705) );
  AOI22_X1 U5028 ( .A1(n7700), .A2(n32666), .B1(n7699), .B2(n34185), .ZN(
        n33704) );
  AOI22_X1 U5029 ( .A1(n7698), .A2(n32682), .B1(n7697), .B2(n32670), .ZN(
        n33703) );
  NAND4_X1 U5030 ( .A1(n33706), .A2(n33705), .A3(n33704), .A4(n33703), .ZN(
        n33712) );
  AOI22_X1 U5031 ( .A1(n7696), .A2(n34194), .B1(n7695), .B2(n34193), .ZN(
        n33710) );
  AOI22_X1 U5032 ( .A1(n7694), .A2(n32681), .B1(n7693), .B2(n32669), .ZN(
        n33709) );
  AOI22_X1 U5033 ( .A1(n7692), .A2(n34198), .B1(n7691), .B2(n32668), .ZN(
        n33708) );
  AOI22_X1 U5034 ( .A1(n7690), .A2(n34200), .B1(n7689), .B2(n34199), .ZN(
        n33707) );
  NAND4_X1 U5035 ( .A1(n33710), .A2(n33709), .A3(n33708), .A4(n33707), .ZN(
        n33711) );
  NOR4_X1 U5036 ( .A1(n33714), .A2(n33713), .A3(n33712), .A4(n33711), .ZN(
        n33715) );
  OAI22_X1 U5037 ( .A1(n33715), .A2(n32665), .B1(n32730), .B2(n32722), .ZN(
        n5821) );
  AOI22_X1 U5038 ( .A1(n7752), .A2(n32716), .B1(n7751), .B2(n32676), .ZN(
        n33719) );
  AOI22_X1 U5039 ( .A1(n7750), .A2(n32678), .B1(n7749), .B2(n32675), .ZN(
        n33718) );
  AOI22_X1 U5040 ( .A1(n7748), .A2(n32667), .B1(n7747), .B2(n34161), .ZN(
        n33717) );
  AOI22_X1 U5041 ( .A1(n7746), .A2(n32677), .B1(n7745), .B2(n32674), .ZN(
        n33716) );
  NAND4_X1 U5042 ( .A1(n33719), .A2(n33718), .A3(n33717), .A4(n33716), .ZN(
        n33735) );
  AOI22_X1 U5043 ( .A1(n7744), .A2(n34170), .B1(n7743), .B2(n34169), .ZN(
        n33723) );
  AOI22_X1 U5044 ( .A1(n7742), .A2(n32680), .B1(n7741), .B2(n34171), .ZN(
        n33722) );
  AOI22_X1 U5045 ( .A1(n7740), .A2(n32679), .B1(n7739), .B2(n32673), .ZN(
        n33721) );
  AOI22_X1 U5046 ( .A1(n7738), .A2(n32719), .B1(n7737), .B2(n32672), .ZN(
        n33720) );
  NAND4_X1 U5047 ( .A1(n33723), .A2(n33722), .A3(n33721), .A4(n33720), .ZN(
        n33734) );
  AOI22_X1 U5048 ( .A1(n7736), .A2(n34182), .B1(n7735), .B2(n32671), .ZN(
        n33727) );
  AOI22_X1 U5049 ( .A1(n7734), .A2(n34184), .B1(n7733), .B2(n34183), .ZN(
        n33726) );
  AOI22_X1 U5050 ( .A1(n7732), .A2(n32666), .B1(n7731), .B2(n34185), .ZN(
        n33725) );
  AOI22_X1 U5051 ( .A1(n7730), .A2(n32682), .B1(n7729), .B2(n32670), .ZN(
        n33724) );
  NAND4_X1 U5052 ( .A1(n33727), .A2(n33726), .A3(n33725), .A4(n33724), .ZN(
        n33733) );
  AOI22_X1 U5053 ( .A1(n7728), .A2(n34194), .B1(n7727), .B2(n34193), .ZN(
        n33731) );
  AOI22_X1 U5054 ( .A1(n7726), .A2(n32681), .B1(n7725), .B2(n32669), .ZN(
        n33730) );
  AOI22_X1 U5055 ( .A1(n7724), .A2(n34198), .B1(n7723), .B2(n32668), .ZN(
        n33729) );
  AOI22_X1 U5056 ( .A1(n7722), .A2(n34200), .B1(n7721), .B2(n32721), .ZN(
        n33728) );
  NAND4_X1 U5057 ( .A1(n33731), .A2(n33730), .A3(n33729), .A4(n33728), .ZN(
        n33732) );
  NOR4_X1 U5058 ( .A1(n33735), .A2(n33734), .A3(n33733), .A4(n33732), .ZN(
        n33736) );
  OAI22_X1 U5059 ( .A1(n33736), .A2(n32665), .B1(n14134), .B2(n32722), .ZN(
        n5822) );
  AOI22_X1 U5060 ( .A1(n7784), .A2(n32716), .B1(n7783), .B2(n32676), .ZN(
        n33740) );
  AOI22_X1 U5061 ( .A1(n7782), .A2(n32678), .B1(n7781), .B2(n32675), .ZN(
        n33739) );
  AOI22_X1 U5062 ( .A1(n7780), .A2(n32667), .B1(n7779), .B2(n34161), .ZN(
        n33738) );
  AOI22_X1 U5063 ( .A1(n7778), .A2(n32677), .B1(n7777), .B2(n32674), .ZN(
        n33737) );
  NAND4_X1 U5064 ( .A1(n33740), .A2(n33739), .A3(n33738), .A4(n33737), .ZN(
        n33756) );
  AOI22_X1 U5065 ( .A1(n7776), .A2(n34170), .B1(n7775), .B2(n34169), .ZN(
        n33744) );
  AOI22_X1 U5066 ( .A1(n7774), .A2(n32680), .B1(n7773), .B2(n32718), .ZN(
        n33743) );
  AOI22_X1 U5067 ( .A1(n7772), .A2(n32679), .B1(n7771), .B2(n32673), .ZN(
        n33742) );
  AOI22_X1 U5068 ( .A1(n7770), .A2(n32719), .B1(n7769), .B2(n32672), .ZN(
        n33741) );
  NAND4_X1 U5069 ( .A1(n33744), .A2(n33743), .A3(n33742), .A4(n33741), .ZN(
        n33755) );
  AOI22_X1 U5070 ( .A1(n7768), .A2(n34182), .B1(n7767), .B2(n32671), .ZN(
        n33748) );
  AOI22_X1 U5071 ( .A1(n7766), .A2(n34184), .B1(n7765), .B2(n34183), .ZN(
        n33747) );
  AOI22_X1 U5072 ( .A1(n7764), .A2(n32666), .B1(n7763), .B2(n34185), .ZN(
        n33746) );
  AOI22_X1 U5073 ( .A1(n7762), .A2(n32682), .B1(n7761), .B2(n32670), .ZN(
        n33745) );
  NAND4_X1 U5074 ( .A1(n33748), .A2(n33747), .A3(n33746), .A4(n33745), .ZN(
        n33754) );
  AOI22_X1 U5075 ( .A1(n7760), .A2(n34194), .B1(n7759), .B2(n34193), .ZN(
        n33752) );
  AOI22_X1 U5076 ( .A1(n7758), .A2(n32681), .B1(n7757), .B2(n32669), .ZN(
        n33751) );
  AOI22_X1 U5077 ( .A1(n7756), .A2(n34198), .B1(n7755), .B2(n32668), .ZN(
        n33750) );
  AOI22_X1 U5078 ( .A1(n7754), .A2(n34200), .B1(n7753), .B2(n32721), .ZN(
        n33749) );
  NAND4_X1 U5079 ( .A1(n33752), .A2(n33751), .A3(n33750), .A4(n33749), .ZN(
        n33753) );
  NOR4_X1 U5080 ( .A1(n33756), .A2(n33755), .A3(n33754), .A4(n33753), .ZN(
        n33757) );
  OAI22_X1 U5081 ( .A1(n33757), .A2(n32665), .B1(n14135), .B2(n32722), .ZN(
        n5823) );
  AOI22_X1 U5082 ( .A1(n7816), .A2(n32716), .B1(n7815), .B2(n32676), .ZN(
        n33761) );
  AOI22_X1 U5083 ( .A1(n7814), .A2(n32678), .B1(n7813), .B2(n32675), .ZN(
        n33760) );
  AOI22_X1 U5084 ( .A1(n7812), .A2(n32667), .B1(n7811), .B2(n34161), .ZN(
        n33759) );
  AOI22_X1 U5085 ( .A1(n7810), .A2(n32677), .B1(n7809), .B2(n32674), .ZN(
        n33758) );
  NAND4_X1 U5086 ( .A1(n33761), .A2(n33760), .A3(n33759), .A4(n33758), .ZN(
        n33777) );
  AOI22_X1 U5087 ( .A1(n7808), .A2(n34170), .B1(n7807), .B2(n32717), .ZN(
        n33765) );
  AOI22_X1 U5088 ( .A1(n7806), .A2(n32680), .B1(n7805), .B2(n32718), .ZN(
        n33764) );
  AOI22_X1 U5089 ( .A1(n7804), .A2(n32679), .B1(n7803), .B2(n32673), .ZN(
        n33763) );
  AOI22_X1 U5090 ( .A1(n7802), .A2(n32719), .B1(n7801), .B2(n32672), .ZN(
        n33762) );
  NAND4_X1 U5091 ( .A1(n33765), .A2(n33764), .A3(n33763), .A4(n33762), .ZN(
        n33776) );
  AOI22_X1 U5092 ( .A1(n7800), .A2(n34182), .B1(n7799), .B2(n32671), .ZN(
        n33769) );
  AOI22_X1 U5093 ( .A1(n7798), .A2(n34184), .B1(n7797), .B2(n34183), .ZN(
        n33768) );
  AOI22_X1 U5094 ( .A1(n7796), .A2(n32666), .B1(n7795), .B2(n34185), .ZN(
        n33767) );
  AOI22_X1 U5095 ( .A1(n7794), .A2(n32682), .B1(n7793), .B2(n32670), .ZN(
        n33766) );
  NAND4_X1 U5096 ( .A1(n33769), .A2(n33768), .A3(n33767), .A4(n33766), .ZN(
        n33775) );
  AOI22_X1 U5097 ( .A1(n7792), .A2(n34194), .B1(n7791), .B2(n32720), .ZN(
        n33773) );
  AOI22_X1 U5098 ( .A1(n7790), .A2(n32681), .B1(n7789), .B2(n32669), .ZN(
        n33772) );
  AOI22_X1 U5099 ( .A1(n7788), .A2(n34198), .B1(n7787), .B2(n32668), .ZN(
        n33771) );
  AOI22_X1 U5100 ( .A1(n7786), .A2(n34200), .B1(n7785), .B2(n32721), .ZN(
        n33770) );
  NAND4_X1 U5101 ( .A1(n33773), .A2(n33772), .A3(n33771), .A4(n33770), .ZN(
        n33774) );
  NOR4_X1 U5102 ( .A1(n33777), .A2(n33776), .A3(n33775), .A4(n33774), .ZN(
        n33778) );
  OAI22_X1 U5103 ( .A1(n33778), .A2(n32665), .B1(n14136), .B2(n32722), .ZN(
        n5824) );
  AOI22_X1 U5104 ( .A1(n7848), .A2(n32716), .B1(n7847), .B2(n32676), .ZN(
        n33782) );
  AOI22_X1 U5105 ( .A1(n7846), .A2(n32678), .B1(n7845), .B2(n32675), .ZN(
        n33781) );
  AOI22_X1 U5106 ( .A1(n7844), .A2(n32667), .B1(n7843), .B2(n34161), .ZN(
        n33780) );
  AOI22_X1 U5107 ( .A1(n7842), .A2(n32677), .B1(n7841), .B2(n32674), .ZN(
        n33779) );
  NAND4_X1 U5108 ( .A1(n33782), .A2(n33781), .A3(n33780), .A4(n33779), .ZN(
        n33798) );
  AOI22_X1 U5109 ( .A1(n7840), .A2(n34170), .B1(n7839), .B2(n32717), .ZN(
        n33786) );
  AOI22_X1 U5110 ( .A1(n7838), .A2(n32680), .B1(n7837), .B2(n32718), .ZN(
        n33785) );
  AOI22_X1 U5111 ( .A1(n7836), .A2(n32679), .B1(n7835), .B2(n32673), .ZN(
        n33784) );
  AOI22_X1 U5112 ( .A1(n7834), .A2(n32719), .B1(n7833), .B2(n32672), .ZN(
        n33783) );
  NAND4_X1 U5113 ( .A1(n33786), .A2(n33785), .A3(n33784), .A4(n33783), .ZN(
        n33797) );
  AOI22_X1 U5114 ( .A1(n7832), .A2(n34182), .B1(n7831), .B2(n32671), .ZN(
        n33790) );
  AOI22_X1 U5115 ( .A1(n7830), .A2(n34184), .B1(n7829), .B2(n34183), .ZN(
        n33789) );
  AOI22_X1 U5116 ( .A1(n7828), .A2(n32666), .B1(n7827), .B2(n34185), .ZN(
        n33788) );
  AOI22_X1 U5117 ( .A1(n7826), .A2(n32682), .B1(n7825), .B2(n32670), .ZN(
        n33787) );
  NAND4_X1 U5118 ( .A1(n33790), .A2(n33789), .A3(n33788), .A4(n33787), .ZN(
        n33796) );
  AOI22_X1 U5119 ( .A1(n7824), .A2(n34194), .B1(n7823), .B2(n32720), .ZN(
        n33794) );
  AOI22_X1 U5120 ( .A1(n7822), .A2(n32681), .B1(n7821), .B2(n32669), .ZN(
        n33793) );
  AOI22_X1 U5121 ( .A1(n7820), .A2(n34198), .B1(n7819), .B2(n32668), .ZN(
        n33792) );
  AOI22_X1 U5122 ( .A1(n7818), .A2(n34200), .B1(n7817), .B2(n32721), .ZN(
        n33791) );
  NAND4_X1 U5123 ( .A1(n33794), .A2(n33793), .A3(n33792), .A4(n33791), .ZN(
        n33795) );
  NOR4_X1 U5124 ( .A1(n33798), .A2(n33797), .A3(n33796), .A4(n33795), .ZN(
        n33799) );
  OAI22_X1 U5125 ( .A1(n33799), .A2(n32665), .B1(n14137), .B2(n32722), .ZN(
        n5825) );
  AOI22_X1 U5126 ( .A1(n7880), .A2(n32716), .B1(n7879), .B2(n32676), .ZN(
        n33803) );
  AOI22_X1 U5127 ( .A1(n7878), .A2(n32678), .B1(n7877), .B2(n32675), .ZN(
        n33802) );
  AOI22_X1 U5128 ( .A1(n7876), .A2(n32667), .B1(n7875), .B2(n34161), .ZN(
        n33801) );
  AOI22_X1 U5129 ( .A1(n7874), .A2(n32677), .B1(n7873), .B2(n32674), .ZN(
        n33800) );
  NAND4_X1 U5130 ( .A1(n33803), .A2(n33802), .A3(n33801), .A4(n33800), .ZN(
        n33819) );
  AOI22_X1 U5131 ( .A1(n7872), .A2(n34170), .B1(n7871), .B2(n32717), .ZN(
        n33807) );
  AOI22_X1 U5132 ( .A1(n7870), .A2(n32680), .B1(n7869), .B2(n32718), .ZN(
        n33806) );
  AOI22_X1 U5133 ( .A1(n7868), .A2(n32679), .B1(n7867), .B2(n32673), .ZN(
        n33805) );
  AOI22_X1 U5134 ( .A1(n7866), .A2(n32719), .B1(n7865), .B2(n32672), .ZN(
        n33804) );
  NAND4_X1 U5135 ( .A1(n33807), .A2(n33806), .A3(n33805), .A4(n33804), .ZN(
        n33818) );
  AOI22_X1 U5136 ( .A1(n7864), .A2(n34182), .B1(n7863), .B2(n32671), .ZN(
        n33811) );
  AOI22_X1 U5137 ( .A1(n7862), .A2(n34184), .B1(n7861), .B2(n34183), .ZN(
        n33810) );
  AOI22_X1 U5138 ( .A1(n7860), .A2(n32666), .B1(n7859), .B2(n34185), .ZN(
        n33809) );
  AOI22_X1 U5139 ( .A1(n7858), .A2(n32682), .B1(n7857), .B2(n32670), .ZN(
        n33808) );
  NAND4_X1 U5140 ( .A1(n33811), .A2(n33810), .A3(n33809), .A4(n33808), .ZN(
        n33817) );
  AOI22_X1 U5141 ( .A1(n7856), .A2(n34194), .B1(n7855), .B2(n32720), .ZN(
        n33815) );
  AOI22_X1 U5142 ( .A1(n7854), .A2(n32681), .B1(n7853), .B2(n32669), .ZN(
        n33814) );
  AOI22_X1 U5143 ( .A1(n7852), .A2(n34198), .B1(n7851), .B2(n32668), .ZN(
        n33813) );
  AOI22_X1 U5144 ( .A1(n7850), .A2(n34200), .B1(n7849), .B2(n32721), .ZN(
        n33812) );
  NAND4_X1 U5145 ( .A1(n33815), .A2(n33814), .A3(n33813), .A4(n33812), .ZN(
        n33816) );
  NOR4_X1 U5146 ( .A1(n33819), .A2(n33818), .A3(n33817), .A4(n33816), .ZN(
        n33820) );
  OAI22_X1 U5147 ( .A1(n33820), .A2(n32665), .B1(n32729), .B2(n32722), .ZN(
        n5826) );
  AOI22_X1 U5148 ( .A1(n7912), .A2(n32716), .B1(n7911), .B2(n32676), .ZN(
        n33824) );
  AOI22_X1 U5149 ( .A1(n7910), .A2(n32678), .B1(n7909), .B2(n32675), .ZN(
        n33823) );
  AOI22_X1 U5150 ( .A1(n7908), .A2(n32667), .B1(n7907), .B2(n34161), .ZN(
        n33822) );
  AOI22_X1 U5151 ( .A1(n7906), .A2(n32677), .B1(n7905), .B2(n32674), .ZN(
        n33821) );
  NAND4_X1 U5152 ( .A1(n33824), .A2(n33823), .A3(n33822), .A4(n33821), .ZN(
        n33840) );
  AOI22_X1 U5153 ( .A1(n7904), .A2(n34170), .B1(n7903), .B2(n32717), .ZN(
        n33828) );
  AOI22_X1 U5154 ( .A1(n7902), .A2(n32680), .B1(n7901), .B2(n32718), .ZN(
        n33827) );
  AOI22_X1 U5155 ( .A1(n7900), .A2(n32679), .B1(n7899), .B2(n32673), .ZN(
        n33826) );
  AOI22_X1 U5156 ( .A1(n7898), .A2(n32719), .B1(n7897), .B2(n32672), .ZN(
        n33825) );
  NAND4_X1 U5157 ( .A1(n33828), .A2(n33827), .A3(n33826), .A4(n33825), .ZN(
        n33839) );
  AOI22_X1 U5158 ( .A1(n7896), .A2(n34182), .B1(n7895), .B2(n32671), .ZN(
        n33832) );
  AOI22_X1 U5159 ( .A1(n7894), .A2(n34184), .B1(n7893), .B2(n34183), .ZN(
        n33831) );
  AOI22_X1 U5160 ( .A1(n7892), .A2(n32666), .B1(n7891), .B2(n34185), .ZN(
        n33830) );
  AOI22_X1 U5161 ( .A1(n7890), .A2(n32682), .B1(n7889), .B2(n32670), .ZN(
        n33829) );
  NAND4_X1 U5162 ( .A1(n33832), .A2(n33831), .A3(n33830), .A4(n33829), .ZN(
        n33838) );
  AOI22_X1 U5163 ( .A1(n7888), .A2(n34194), .B1(n7887), .B2(n32720), .ZN(
        n33836) );
  AOI22_X1 U5164 ( .A1(n7886), .A2(n32681), .B1(n7885), .B2(n32669), .ZN(
        n33835) );
  AOI22_X1 U5165 ( .A1(n7884), .A2(n34198), .B1(n7883), .B2(n32668), .ZN(
        n33834) );
  AOI22_X1 U5166 ( .A1(n7882), .A2(n34200), .B1(n7881), .B2(n32721), .ZN(
        n33833) );
  NAND4_X1 U5167 ( .A1(n33836), .A2(n33835), .A3(n33834), .A4(n33833), .ZN(
        n33837) );
  NOR4_X1 U5168 ( .A1(n33840), .A2(n33839), .A3(n33838), .A4(n33837), .ZN(
        n33841) );
  OAI22_X1 U5169 ( .A1(n33841), .A2(n32665), .B1(n32728), .B2(n32722), .ZN(
        n5827) );
  AOI22_X1 U5170 ( .A1(n7944), .A2(n32716), .B1(n7943), .B2(n32676), .ZN(
        n33845) );
  AOI22_X1 U5171 ( .A1(n7942), .A2(n32678), .B1(n7941), .B2(n32675), .ZN(
        n33844) );
  AOI22_X1 U5172 ( .A1(n7940), .A2(n32667), .B1(n7939), .B2(n34161), .ZN(
        n33843) );
  AOI22_X1 U5173 ( .A1(n7938), .A2(n32677), .B1(n7937), .B2(n32674), .ZN(
        n33842) );
  NAND4_X1 U5174 ( .A1(n33845), .A2(n33844), .A3(n33843), .A4(n33842), .ZN(
        n33861) );
  AOI22_X1 U5175 ( .A1(n7936), .A2(n34170), .B1(n7935), .B2(n32717), .ZN(
        n33849) );
  AOI22_X1 U5176 ( .A1(n7934), .A2(n32680), .B1(n7933), .B2(n32718), .ZN(
        n33848) );
  AOI22_X1 U5177 ( .A1(n7932), .A2(n32679), .B1(n7931), .B2(n32673), .ZN(
        n33847) );
  AOI22_X1 U5178 ( .A1(n7930), .A2(n32719), .B1(n7929), .B2(n32672), .ZN(
        n33846) );
  NAND4_X1 U5179 ( .A1(n33849), .A2(n33848), .A3(n33847), .A4(n33846), .ZN(
        n33860) );
  AOI22_X1 U5180 ( .A1(n7928), .A2(n34182), .B1(n7927), .B2(n32671), .ZN(
        n33853) );
  AOI22_X1 U5181 ( .A1(n7926), .A2(n34184), .B1(n7925), .B2(n34183), .ZN(
        n33852) );
  AOI22_X1 U5182 ( .A1(n7924), .A2(n32666), .B1(n7923), .B2(n34185), .ZN(
        n33851) );
  AOI22_X1 U5183 ( .A1(n7922), .A2(n32682), .B1(n7921), .B2(n32670), .ZN(
        n33850) );
  NAND4_X1 U5184 ( .A1(n33853), .A2(n33852), .A3(n33851), .A4(n33850), .ZN(
        n33859) );
  AOI22_X1 U5185 ( .A1(n7920), .A2(n34194), .B1(n7919), .B2(n32720), .ZN(
        n33857) );
  AOI22_X1 U5186 ( .A1(n7918), .A2(n32681), .B1(n7917), .B2(n32669), .ZN(
        n33856) );
  AOI22_X1 U5187 ( .A1(n7916), .A2(n34198), .B1(n7915), .B2(n32668), .ZN(
        n33855) );
  AOI22_X1 U5188 ( .A1(n7914), .A2(n34200), .B1(n7913), .B2(n32721), .ZN(
        n33854) );
  NAND4_X1 U5189 ( .A1(n33857), .A2(n33856), .A3(n33855), .A4(n33854), .ZN(
        n33858) );
  NOR4_X1 U5190 ( .A1(n33861), .A2(n33860), .A3(n33859), .A4(n33858), .ZN(
        n33862) );
  OAI22_X1 U5191 ( .A1(n33862), .A2(n32665), .B1(n14140), .B2(n32722), .ZN(
        n5828) );
  AOI22_X1 U5192 ( .A1(n7976), .A2(n32716), .B1(n7975), .B2(n32676), .ZN(
        n33866) );
  AOI22_X1 U5193 ( .A1(n7974), .A2(n32678), .B1(n7973), .B2(n32675), .ZN(
        n33865) );
  AOI22_X1 U5194 ( .A1(n7972), .A2(n32667), .B1(n7971), .B2(n34161), .ZN(
        n33864) );
  AOI22_X1 U5195 ( .A1(n7970), .A2(n32677), .B1(n7969), .B2(n32674), .ZN(
        n33863) );
  NAND4_X1 U5196 ( .A1(n33866), .A2(n33865), .A3(n33864), .A4(n33863), .ZN(
        n33882) );
  AOI22_X1 U5197 ( .A1(n7968), .A2(n34170), .B1(n7967), .B2(n32717), .ZN(
        n33870) );
  AOI22_X1 U5198 ( .A1(n7966), .A2(n32680), .B1(n7965), .B2(n32718), .ZN(
        n33869) );
  AOI22_X1 U5199 ( .A1(n7964), .A2(n32679), .B1(n7963), .B2(n32673), .ZN(
        n33868) );
  AOI22_X1 U5200 ( .A1(n7962), .A2(n32719), .B1(n7961), .B2(n32672), .ZN(
        n33867) );
  NAND4_X1 U5201 ( .A1(n33870), .A2(n33869), .A3(n33868), .A4(n33867), .ZN(
        n33881) );
  AOI22_X1 U5202 ( .A1(n7960), .A2(n34182), .B1(n7959), .B2(n32671), .ZN(
        n33874) );
  AOI22_X1 U5203 ( .A1(n7958), .A2(n34184), .B1(n7957), .B2(n34183), .ZN(
        n33873) );
  AOI22_X1 U5204 ( .A1(n7956), .A2(n32666), .B1(n7955), .B2(n34185), .ZN(
        n33872) );
  AOI22_X1 U5205 ( .A1(n7954), .A2(n32682), .B1(n7953), .B2(n32670), .ZN(
        n33871) );
  NAND4_X1 U5206 ( .A1(n33874), .A2(n33873), .A3(n33872), .A4(n33871), .ZN(
        n33880) );
  AOI22_X1 U5207 ( .A1(n7952), .A2(n34194), .B1(n7951), .B2(n32720), .ZN(
        n33878) );
  AOI22_X1 U5208 ( .A1(n7950), .A2(n32681), .B1(n7949), .B2(n32669), .ZN(
        n33877) );
  AOI22_X1 U5209 ( .A1(n7948), .A2(n34198), .B1(n7947), .B2(n32668), .ZN(
        n33876) );
  AOI22_X1 U5210 ( .A1(n7946), .A2(n34200), .B1(n7945), .B2(n32721), .ZN(
        n33875) );
  NAND4_X1 U5211 ( .A1(n33878), .A2(n33877), .A3(n33876), .A4(n33875), .ZN(
        n33879) );
  NOR4_X1 U5212 ( .A1(n33882), .A2(n33881), .A3(n33880), .A4(n33879), .ZN(
        n33883) );
  OAI22_X1 U5213 ( .A1(n33883), .A2(n32665), .B1(n14141), .B2(n32722), .ZN(
        n5829) );
  AOI22_X1 U5214 ( .A1(n8008), .A2(n32716), .B1(n8007), .B2(n32676), .ZN(
        n33887) );
  AOI22_X1 U5215 ( .A1(n8006), .A2(n32678), .B1(n8005), .B2(n32675), .ZN(
        n33886) );
  AOI22_X1 U5216 ( .A1(n8004), .A2(n32667), .B1(n8003), .B2(n34161), .ZN(
        n33885) );
  AOI22_X1 U5217 ( .A1(n8002), .A2(n32677), .B1(n8001), .B2(n32674), .ZN(
        n33884) );
  NAND4_X1 U5218 ( .A1(n33887), .A2(n33886), .A3(n33885), .A4(n33884), .ZN(
        n33903) );
  AOI22_X1 U5219 ( .A1(n8000), .A2(n34170), .B1(n7999), .B2(n32717), .ZN(
        n33891) );
  AOI22_X1 U5220 ( .A1(n7998), .A2(n32680), .B1(n7997), .B2(n32718), .ZN(
        n33890) );
  AOI22_X1 U5221 ( .A1(n7996), .A2(n32679), .B1(n7995), .B2(n32673), .ZN(
        n33889) );
  AOI22_X1 U5222 ( .A1(n7994), .A2(n32719), .B1(n7993), .B2(n32672), .ZN(
        n33888) );
  NAND4_X1 U5223 ( .A1(n33891), .A2(n33890), .A3(n33889), .A4(n33888), .ZN(
        n33902) );
  AOI22_X1 U5224 ( .A1(n7992), .A2(n34182), .B1(n7991), .B2(n32671), .ZN(
        n33895) );
  AOI22_X1 U5225 ( .A1(n7990), .A2(n34184), .B1(n7989), .B2(n34183), .ZN(
        n33894) );
  AOI22_X1 U5226 ( .A1(n7988), .A2(n32666), .B1(n7987), .B2(n34185), .ZN(
        n33893) );
  AOI22_X1 U5227 ( .A1(n7986), .A2(n32682), .B1(n7985), .B2(n32670), .ZN(
        n33892) );
  NAND4_X1 U5228 ( .A1(n33895), .A2(n33894), .A3(n33893), .A4(n33892), .ZN(
        n33901) );
  AOI22_X1 U5229 ( .A1(n7984), .A2(n34194), .B1(n7983), .B2(n32720), .ZN(
        n33899) );
  AOI22_X1 U5230 ( .A1(n7982), .A2(n32681), .B1(n7981), .B2(n32669), .ZN(
        n33898) );
  AOI22_X1 U5231 ( .A1(n7980), .A2(n34198), .B1(n7979), .B2(n32668), .ZN(
        n33897) );
  AOI22_X1 U5232 ( .A1(n7978), .A2(n34200), .B1(n7977), .B2(n32721), .ZN(
        n33896) );
  NAND4_X1 U5233 ( .A1(n33899), .A2(n33898), .A3(n33897), .A4(n33896), .ZN(
        n33900) );
  NOR4_X1 U5234 ( .A1(n33903), .A2(n33902), .A3(n33901), .A4(n33900), .ZN(
        n33904) );
  OAI22_X1 U5235 ( .A1(n33904), .A2(n32665), .B1(n14142), .B2(n32722), .ZN(
        n5830) );
  AOI22_X1 U5236 ( .A1(n8040), .A2(n32716), .B1(n8039), .B2(n32676), .ZN(
        n33908) );
  AOI22_X1 U5237 ( .A1(n8038), .A2(n32678), .B1(n8037), .B2(n32675), .ZN(
        n33907) );
  AOI22_X1 U5238 ( .A1(n8036), .A2(n32667), .B1(n8035), .B2(n34161), .ZN(
        n33906) );
  AOI22_X1 U5239 ( .A1(n8034), .A2(n32677), .B1(n8033), .B2(n32674), .ZN(
        n33905) );
  NAND4_X1 U5240 ( .A1(n33908), .A2(n33907), .A3(n33906), .A4(n33905), .ZN(
        n33924) );
  AOI22_X1 U5241 ( .A1(n8032), .A2(n34170), .B1(n8031), .B2(n32717), .ZN(
        n33912) );
  AOI22_X1 U5242 ( .A1(n8030), .A2(n32680), .B1(n8029), .B2(n32718), .ZN(
        n33911) );
  AOI22_X1 U5243 ( .A1(n8028), .A2(n32679), .B1(n8027), .B2(n32673), .ZN(
        n33910) );
  AOI22_X1 U5244 ( .A1(n8026), .A2(n32719), .B1(n8025), .B2(n32672), .ZN(
        n33909) );
  NAND4_X1 U5245 ( .A1(n33912), .A2(n33911), .A3(n33910), .A4(n33909), .ZN(
        n33923) );
  AOI22_X1 U5246 ( .A1(n8024), .A2(n34182), .B1(n8023), .B2(n32671), .ZN(
        n33916) );
  AOI22_X1 U5247 ( .A1(n8022), .A2(n34184), .B1(n8021), .B2(n34183), .ZN(
        n33915) );
  AOI22_X1 U5248 ( .A1(n8020), .A2(n32666), .B1(n8019), .B2(n34185), .ZN(
        n33914) );
  AOI22_X1 U5249 ( .A1(n8018), .A2(n32682), .B1(n8017), .B2(n32670), .ZN(
        n33913) );
  NAND4_X1 U5250 ( .A1(n33916), .A2(n33915), .A3(n33914), .A4(n33913), .ZN(
        n33922) );
  AOI22_X1 U5251 ( .A1(n8016), .A2(n34194), .B1(n8015), .B2(n32720), .ZN(
        n33920) );
  AOI22_X1 U5252 ( .A1(n8014), .A2(n32681), .B1(n8013), .B2(n32669), .ZN(
        n33919) );
  AOI22_X1 U5253 ( .A1(n8012), .A2(n34198), .B1(n8011), .B2(n32668), .ZN(
        n33918) );
  AOI22_X1 U5254 ( .A1(n8010), .A2(n34200), .B1(n8009), .B2(n32721), .ZN(
        n33917) );
  NAND4_X1 U5255 ( .A1(n33920), .A2(n33919), .A3(n33918), .A4(n33917), .ZN(
        n33921) );
  NOR4_X1 U5256 ( .A1(n33924), .A2(n33923), .A3(n33922), .A4(n33921), .ZN(
        n33925) );
  OAI22_X1 U5257 ( .A1(n33925), .A2(n32665), .B1(n14143), .B2(n32722), .ZN(
        n5831) );
  AOI22_X1 U5258 ( .A1(n8072), .A2(n32716), .B1(n8071), .B2(n32676), .ZN(
        n33929) );
  AOI22_X1 U5259 ( .A1(n8070), .A2(n32678), .B1(n8069), .B2(n32675), .ZN(
        n33928) );
  AOI22_X1 U5260 ( .A1(n8068), .A2(n32667), .B1(n8067), .B2(n34161), .ZN(
        n33927) );
  AOI22_X1 U5261 ( .A1(n8066), .A2(n32677), .B1(n8065), .B2(n32674), .ZN(
        n33926) );
  NAND4_X1 U5262 ( .A1(n33929), .A2(n33928), .A3(n33927), .A4(n33926), .ZN(
        n33945) );
  AOI22_X1 U5263 ( .A1(n8064), .A2(n34170), .B1(n8063), .B2(n32717), .ZN(
        n33933) );
  AOI22_X1 U5264 ( .A1(n8062), .A2(n32680), .B1(n8061), .B2(n32718), .ZN(
        n33932) );
  AOI22_X1 U5265 ( .A1(n8060), .A2(n32679), .B1(n8059), .B2(n32673), .ZN(
        n33931) );
  AOI22_X1 U5266 ( .A1(n8058), .A2(n32719), .B1(n8057), .B2(n32672), .ZN(
        n33930) );
  NAND4_X1 U5267 ( .A1(n33933), .A2(n33932), .A3(n33931), .A4(n33930), .ZN(
        n33944) );
  AOI22_X1 U5268 ( .A1(n8056), .A2(n34182), .B1(n8055), .B2(n32671), .ZN(
        n33937) );
  AOI22_X1 U5269 ( .A1(n8054), .A2(n34184), .B1(n8053), .B2(n34183), .ZN(
        n33936) );
  AOI22_X1 U5270 ( .A1(n8052), .A2(n32666), .B1(n8051), .B2(n34185), .ZN(
        n33935) );
  AOI22_X1 U5271 ( .A1(n8050), .A2(n32682), .B1(n8049), .B2(n32670), .ZN(
        n33934) );
  NAND4_X1 U5272 ( .A1(n33937), .A2(n33936), .A3(n33935), .A4(n33934), .ZN(
        n33943) );
  AOI22_X1 U5273 ( .A1(n8048), .A2(n34194), .B1(n8047), .B2(n32720), .ZN(
        n33941) );
  AOI22_X1 U5274 ( .A1(n8046), .A2(n32681), .B1(n8045), .B2(n32669), .ZN(
        n33940) );
  AOI22_X1 U5275 ( .A1(n8044), .A2(n34198), .B1(n8043), .B2(n32668), .ZN(
        n33939) );
  AOI22_X1 U5276 ( .A1(n8042), .A2(n34200), .B1(n8041), .B2(n32721), .ZN(
        n33938) );
  NAND4_X1 U5277 ( .A1(n33941), .A2(n33940), .A3(n33939), .A4(n33938), .ZN(
        n33942) );
  NOR4_X1 U5278 ( .A1(n33945), .A2(n33944), .A3(n33943), .A4(n33942), .ZN(
        n33946) );
  OAI22_X1 U5279 ( .A1(n33946), .A2(n32665), .B1(n14144), .B2(n32722), .ZN(
        n5832) );
  AOI22_X1 U5280 ( .A1(n8104), .A2(n32716), .B1(n8103), .B2(n32676), .ZN(
        n33950) );
  AOI22_X1 U5281 ( .A1(n8102), .A2(n32678), .B1(n8101), .B2(n32675), .ZN(
        n33949) );
  AOI22_X1 U5282 ( .A1(n8100), .A2(n32667), .B1(n8099), .B2(n34161), .ZN(
        n33948) );
  AOI22_X1 U5283 ( .A1(n8098), .A2(n32677), .B1(n8097), .B2(n32674), .ZN(
        n33947) );
  NAND4_X1 U5284 ( .A1(n33950), .A2(n33949), .A3(n33948), .A4(n33947), .ZN(
        n33966) );
  AOI22_X1 U5285 ( .A1(n8096), .A2(n34170), .B1(n8095), .B2(n32717), .ZN(
        n33954) );
  AOI22_X1 U5286 ( .A1(n8094), .A2(n32680), .B1(n8093), .B2(n32718), .ZN(
        n33953) );
  AOI22_X1 U5287 ( .A1(n8092), .A2(n32679), .B1(n8091), .B2(n32673), .ZN(
        n33952) );
  AOI22_X1 U5288 ( .A1(n8090), .A2(n32719), .B1(n8089), .B2(n32672), .ZN(
        n33951) );
  NAND4_X1 U5289 ( .A1(n33954), .A2(n33953), .A3(n33952), .A4(n33951), .ZN(
        n33965) );
  AOI22_X1 U5290 ( .A1(n8088), .A2(n34182), .B1(n8087), .B2(n32671), .ZN(
        n33958) );
  AOI22_X1 U5291 ( .A1(n8086), .A2(n34184), .B1(n8085), .B2(n34183), .ZN(
        n33957) );
  AOI22_X1 U5292 ( .A1(n8084), .A2(n32666), .B1(n8083), .B2(n34185), .ZN(
        n33956) );
  AOI22_X1 U5293 ( .A1(n8082), .A2(n32682), .B1(n8081), .B2(n32670), .ZN(
        n33955) );
  NAND4_X1 U5294 ( .A1(n33958), .A2(n33957), .A3(n33956), .A4(n33955), .ZN(
        n33964) );
  AOI22_X1 U5295 ( .A1(n8080), .A2(n34194), .B1(n8079), .B2(n32720), .ZN(
        n33962) );
  AOI22_X1 U5296 ( .A1(n8078), .A2(n32681), .B1(n8077), .B2(n32669), .ZN(
        n33961) );
  AOI22_X1 U5297 ( .A1(n8076), .A2(n34198), .B1(n8075), .B2(n32668), .ZN(
        n33960) );
  AOI22_X1 U5298 ( .A1(n8074), .A2(n34200), .B1(n8073), .B2(n32721), .ZN(
        n33959) );
  NAND4_X1 U5299 ( .A1(n33962), .A2(n33961), .A3(n33960), .A4(n33959), .ZN(
        n33963) );
  NOR4_X1 U5300 ( .A1(n33966), .A2(n33965), .A3(n33964), .A4(n33963), .ZN(
        n33967) );
  OAI22_X1 U5301 ( .A1(n33967), .A2(n32665), .B1(n14145), .B2(n32722), .ZN(
        n5833) );
  AOI22_X1 U5302 ( .A1(n8136), .A2(n32716), .B1(n8135), .B2(n32676), .ZN(
        n33971) );
  AOI22_X1 U5303 ( .A1(n8134), .A2(n32678), .B1(n8133), .B2(n32675), .ZN(
        n33970) );
  AOI22_X1 U5304 ( .A1(n8132), .A2(n32667), .B1(n8131), .B2(n34161), .ZN(
        n33969) );
  AOI22_X1 U5305 ( .A1(n8130), .A2(n32677), .B1(n8129), .B2(n32674), .ZN(
        n33968) );
  NAND4_X1 U5306 ( .A1(n33971), .A2(n33970), .A3(n33969), .A4(n33968), .ZN(
        n33987) );
  AOI22_X1 U5307 ( .A1(n8128), .A2(n34170), .B1(n8127), .B2(n32717), .ZN(
        n33975) );
  AOI22_X1 U5308 ( .A1(n8126), .A2(n32680), .B1(n8125), .B2(n32718), .ZN(
        n33974) );
  AOI22_X1 U5309 ( .A1(n8124), .A2(n32679), .B1(n8123), .B2(n32673), .ZN(
        n33973) );
  AOI22_X1 U5310 ( .A1(n8122), .A2(n32719), .B1(n8121), .B2(n32672), .ZN(
        n33972) );
  NAND4_X1 U5311 ( .A1(n33975), .A2(n33974), .A3(n33973), .A4(n33972), .ZN(
        n33986) );
  AOI22_X1 U5312 ( .A1(n8120), .A2(n34182), .B1(n8119), .B2(n32671), .ZN(
        n33979) );
  AOI22_X1 U5313 ( .A1(n8118), .A2(n34184), .B1(n8117), .B2(n34183), .ZN(
        n33978) );
  AOI22_X1 U5314 ( .A1(n8116), .A2(n32666), .B1(n8115), .B2(n34185), .ZN(
        n33977) );
  AOI22_X1 U5315 ( .A1(n8114), .A2(n32682), .B1(n8113), .B2(n32670), .ZN(
        n33976) );
  NAND4_X1 U5316 ( .A1(n33979), .A2(n33978), .A3(n33977), .A4(n33976), .ZN(
        n33985) );
  AOI22_X1 U5317 ( .A1(n8112), .A2(n34194), .B1(n8111), .B2(n32720), .ZN(
        n33983) );
  AOI22_X1 U5318 ( .A1(n8110), .A2(n32681), .B1(n8109), .B2(n32669), .ZN(
        n33982) );
  AOI22_X1 U5319 ( .A1(n8108), .A2(n34198), .B1(n8107), .B2(n32668), .ZN(
        n33981) );
  AOI22_X1 U5320 ( .A1(n8106), .A2(n34200), .B1(n8105), .B2(n32721), .ZN(
        n33980) );
  NAND4_X1 U5321 ( .A1(n33983), .A2(n33982), .A3(n33981), .A4(n33980), .ZN(
        n33984) );
  NOR4_X1 U5322 ( .A1(n33987), .A2(n33986), .A3(n33985), .A4(n33984), .ZN(
        n33988) );
  OAI22_X1 U5323 ( .A1(n33988), .A2(n32665), .B1(n32727), .B2(n32722), .ZN(
        n5834) );
  AOI22_X1 U5324 ( .A1(n8168), .A2(n32716), .B1(n8167), .B2(n32676), .ZN(
        n33992) );
  AOI22_X1 U5325 ( .A1(n8166), .A2(n32678), .B1(n8165), .B2(n32675), .ZN(
        n33991) );
  AOI22_X1 U5326 ( .A1(n8164), .A2(n32667), .B1(n8163), .B2(n34161), .ZN(
        n33990) );
  AOI22_X1 U5327 ( .A1(n8162), .A2(n32677), .B1(n8161), .B2(n32674), .ZN(
        n33989) );
  NAND4_X1 U5328 ( .A1(n33992), .A2(n33991), .A3(n33990), .A4(n33989), .ZN(
        n34008) );
  AOI22_X1 U5329 ( .A1(n8160), .A2(n34170), .B1(n8159), .B2(n32717), .ZN(
        n33996) );
  AOI22_X1 U5330 ( .A1(n8158), .A2(n32680), .B1(n8157), .B2(n32718), .ZN(
        n33995) );
  AOI22_X1 U5331 ( .A1(n8156), .A2(n32679), .B1(n8155), .B2(n32673), .ZN(
        n33994) );
  AOI22_X1 U5332 ( .A1(n8154), .A2(n32719), .B1(n8153), .B2(n32672), .ZN(
        n33993) );
  NAND4_X1 U5333 ( .A1(n33996), .A2(n33995), .A3(n33994), .A4(n33993), .ZN(
        n34007) );
  AOI22_X1 U5334 ( .A1(n8152), .A2(n34182), .B1(n8151), .B2(n32671), .ZN(
        n34000) );
  AOI22_X1 U5335 ( .A1(n8150), .A2(n34184), .B1(n8149), .B2(n34183), .ZN(
        n33999) );
  AOI22_X1 U5336 ( .A1(n8148), .A2(n32666), .B1(n8147), .B2(n34185), .ZN(
        n33998) );
  AOI22_X1 U5337 ( .A1(n8146), .A2(n32682), .B1(n8145), .B2(n32670), .ZN(
        n33997) );
  NAND4_X1 U5338 ( .A1(n34000), .A2(n33999), .A3(n33998), .A4(n33997), .ZN(
        n34006) );
  AOI22_X1 U5339 ( .A1(n8144), .A2(n34194), .B1(n8143), .B2(n32720), .ZN(
        n34004) );
  AOI22_X1 U5340 ( .A1(n8142), .A2(n32681), .B1(n8141), .B2(n32669), .ZN(
        n34003) );
  AOI22_X1 U5341 ( .A1(n8140), .A2(n34198), .B1(n8139), .B2(n32668), .ZN(
        n34002) );
  AOI22_X1 U5342 ( .A1(n8138), .A2(n34200), .B1(n8137), .B2(n32721), .ZN(
        n34001) );
  NAND4_X1 U5343 ( .A1(n34004), .A2(n34003), .A3(n34002), .A4(n34001), .ZN(
        n34005) );
  NOR4_X1 U5344 ( .A1(n34008), .A2(n34007), .A3(n34006), .A4(n34005), .ZN(
        n34009) );
  OAI22_X1 U5345 ( .A1(n34009), .A2(n32665), .B1(n32726), .B2(n32722), .ZN(
        n5835) );
  AOI22_X1 U5346 ( .A1(n8200), .A2(n32716), .B1(n8199), .B2(n32676), .ZN(
        n34013) );
  AOI22_X1 U5347 ( .A1(n8198), .A2(n32678), .B1(n8197), .B2(n32675), .ZN(
        n34012) );
  AOI22_X1 U5348 ( .A1(n8196), .A2(n32667), .B1(n8195), .B2(n34161), .ZN(
        n34011) );
  AOI22_X1 U5349 ( .A1(n8194), .A2(n32677), .B1(n8193), .B2(n32674), .ZN(
        n34010) );
  NAND4_X1 U5350 ( .A1(n34013), .A2(n34012), .A3(n34011), .A4(n34010), .ZN(
        n34029) );
  AOI22_X1 U5351 ( .A1(n8192), .A2(n34170), .B1(n8191), .B2(n34169), .ZN(
        n34017) );
  AOI22_X1 U5352 ( .A1(n8190), .A2(n32680), .B1(n8189), .B2(n34171), .ZN(
        n34016) );
  AOI22_X1 U5353 ( .A1(n8188), .A2(n32679), .B1(n8187), .B2(n32673), .ZN(
        n34015) );
  AOI22_X1 U5354 ( .A1(n8186), .A2(n32719), .B1(n8185), .B2(n32672), .ZN(
        n34014) );
  NAND4_X1 U5355 ( .A1(n34017), .A2(n34016), .A3(n34015), .A4(n34014), .ZN(
        n34028) );
  AOI22_X1 U5356 ( .A1(n8184), .A2(n34182), .B1(n8183), .B2(n32671), .ZN(
        n34021) );
  AOI22_X1 U5357 ( .A1(n8182), .A2(n34184), .B1(n8181), .B2(n34183), .ZN(
        n34020) );
  AOI22_X1 U5358 ( .A1(n8180), .A2(n32666), .B1(n8179), .B2(n34185), .ZN(
        n34019) );
  AOI22_X1 U5359 ( .A1(n8178), .A2(n32682), .B1(n8177), .B2(n32670), .ZN(
        n34018) );
  NAND4_X1 U5360 ( .A1(n34021), .A2(n34020), .A3(n34019), .A4(n34018), .ZN(
        n34027) );
  AOI22_X1 U5361 ( .A1(n8176), .A2(n34194), .B1(n8175), .B2(n34193), .ZN(
        n34025) );
  AOI22_X1 U5362 ( .A1(n8174), .A2(n32681), .B1(n8173), .B2(n32669), .ZN(
        n34024) );
  AOI22_X1 U5363 ( .A1(n8172), .A2(n34198), .B1(n8171), .B2(n32668), .ZN(
        n34023) );
  AOI22_X1 U5364 ( .A1(n8170), .A2(n34200), .B1(n8169), .B2(n34199), .ZN(
        n34022) );
  NAND4_X1 U5365 ( .A1(n34025), .A2(n34024), .A3(n34023), .A4(n34022), .ZN(
        n34026) );
  NOR4_X1 U5366 ( .A1(n34029), .A2(n34028), .A3(n34027), .A4(n34026), .ZN(
        n34030) );
  OAI22_X1 U5367 ( .A1(n34030), .A2(n32665), .B1(n14148), .B2(n32722), .ZN(
        n5836) );
  AOI22_X1 U5368 ( .A1(n8232), .A2(n32716), .B1(n8231), .B2(n32676), .ZN(
        n34034) );
  AOI22_X1 U5369 ( .A1(n8230), .A2(n32678), .B1(n8229), .B2(n32675), .ZN(
        n34033) );
  AOI22_X1 U5370 ( .A1(n8228), .A2(n32667), .B1(n8227), .B2(n34161), .ZN(
        n34032) );
  AOI22_X1 U5371 ( .A1(n8226), .A2(n32677), .B1(n8225), .B2(n32674), .ZN(
        n34031) );
  NAND4_X1 U5372 ( .A1(n34034), .A2(n34033), .A3(n34032), .A4(n34031), .ZN(
        n34050) );
  AOI22_X1 U5373 ( .A1(n8224), .A2(n34170), .B1(n8223), .B2(n34169), .ZN(
        n34038) );
  AOI22_X1 U5374 ( .A1(n8222), .A2(n32680), .B1(n8221), .B2(n34171), .ZN(
        n34037) );
  AOI22_X1 U5375 ( .A1(n8220), .A2(n32679), .B1(n8219), .B2(n32673), .ZN(
        n34036) );
  AOI22_X1 U5376 ( .A1(n8218), .A2(n32719), .B1(n8217), .B2(n32672), .ZN(
        n34035) );
  NAND4_X1 U5377 ( .A1(n34038), .A2(n34037), .A3(n34036), .A4(n34035), .ZN(
        n34049) );
  AOI22_X1 U5378 ( .A1(n8216), .A2(n34182), .B1(n8215), .B2(n32671), .ZN(
        n34042) );
  AOI22_X1 U5379 ( .A1(n8214), .A2(n34184), .B1(n8213), .B2(n34183), .ZN(
        n34041) );
  AOI22_X1 U5380 ( .A1(n8212), .A2(n32666), .B1(n8211), .B2(n34185), .ZN(
        n34040) );
  AOI22_X1 U5381 ( .A1(n8210), .A2(n32682), .B1(n8209), .B2(n32670), .ZN(
        n34039) );
  NAND4_X1 U5382 ( .A1(n34042), .A2(n34041), .A3(n34040), .A4(n34039), .ZN(
        n34048) );
  AOI22_X1 U5383 ( .A1(n8208), .A2(n34194), .B1(n8207), .B2(n34193), .ZN(
        n34046) );
  AOI22_X1 U5384 ( .A1(n8206), .A2(n32681), .B1(n8205), .B2(n32669), .ZN(
        n34045) );
  AOI22_X1 U5385 ( .A1(n8204), .A2(n34198), .B1(n8203), .B2(n32668), .ZN(
        n34044) );
  AOI22_X1 U5386 ( .A1(n8202), .A2(n34200), .B1(n8201), .B2(n34199), .ZN(
        n34043) );
  NAND4_X1 U5387 ( .A1(n34046), .A2(n34045), .A3(n34044), .A4(n34043), .ZN(
        n34047) );
  NOR4_X1 U5388 ( .A1(n34050), .A2(n34049), .A3(n34048), .A4(n34047), .ZN(
        n34051) );
  OAI22_X1 U5389 ( .A1(n34051), .A2(n32665), .B1(n14149), .B2(n32722), .ZN(
        n5837) );
  AOI22_X1 U5390 ( .A1(n8264), .A2(n34158), .B1(n8263), .B2(n32676), .ZN(
        n34055) );
  AOI22_X1 U5391 ( .A1(n8262), .A2(n32678), .B1(n8261), .B2(n32675), .ZN(
        n34054) );
  AOI22_X1 U5392 ( .A1(n8260), .A2(n32667), .B1(n8259), .B2(n34161), .ZN(
        n34053) );
  AOI22_X1 U5393 ( .A1(n8258), .A2(n32677), .B1(n8257), .B2(n32674), .ZN(
        n34052) );
  NAND4_X1 U5394 ( .A1(n34055), .A2(n34054), .A3(n34053), .A4(n34052), .ZN(
        n34071) );
  AOI22_X1 U5395 ( .A1(n8256), .A2(n34170), .B1(n8255), .B2(n34169), .ZN(
        n34059) );
  AOI22_X1 U5396 ( .A1(n8254), .A2(n32680), .B1(n8253), .B2(n34171), .ZN(
        n34058) );
  AOI22_X1 U5397 ( .A1(n8252), .A2(n32679), .B1(n8251), .B2(n32673), .ZN(
        n34057) );
  AOI22_X1 U5398 ( .A1(n8250), .A2(n32719), .B1(n8249), .B2(n32672), .ZN(
        n34056) );
  NAND4_X1 U5399 ( .A1(n34059), .A2(n34058), .A3(n34057), .A4(n34056), .ZN(
        n34070) );
  AOI22_X1 U5400 ( .A1(n8248), .A2(n34182), .B1(n8247), .B2(n32671), .ZN(
        n34063) );
  AOI22_X1 U5401 ( .A1(n8246), .A2(n34184), .B1(n8245), .B2(n34183), .ZN(
        n34062) );
  AOI22_X1 U5402 ( .A1(n8244), .A2(n34186), .B1(n8243), .B2(n34185), .ZN(
        n34061) );
  AOI22_X1 U5403 ( .A1(n8242), .A2(n32682), .B1(n8241), .B2(n32670), .ZN(
        n34060) );
  NAND4_X1 U5404 ( .A1(n34063), .A2(n34062), .A3(n34061), .A4(n34060), .ZN(
        n34069) );
  AOI22_X1 U5405 ( .A1(n8240), .A2(n34194), .B1(n8239), .B2(n34193), .ZN(
        n34067) );
  AOI22_X1 U5406 ( .A1(n8238), .A2(n32681), .B1(n8237), .B2(n32669), .ZN(
        n34066) );
  AOI22_X1 U5407 ( .A1(n8236), .A2(n34198), .B1(n8235), .B2(n32668), .ZN(
        n34065) );
  AOI22_X1 U5408 ( .A1(n8234), .A2(n34200), .B1(n8233), .B2(n34199), .ZN(
        n34064) );
  NAND4_X1 U5409 ( .A1(n34067), .A2(n34066), .A3(n34065), .A4(n34064), .ZN(
        n34068) );
  NOR4_X1 U5410 ( .A1(n34071), .A2(n34070), .A3(n34069), .A4(n34068), .ZN(
        n34072) );
  OAI22_X1 U5411 ( .A1(n34072), .A2(n34210), .B1(n14150), .B2(n32722), .ZN(
        n5838) );
  AOI22_X1 U5412 ( .A1(n8296), .A2(n32716), .B1(n8295), .B2(n32676), .ZN(
        n34076) );
  AOI22_X1 U5413 ( .A1(n8294), .A2(n32678), .B1(n8293), .B2(n32675), .ZN(
        n34075) );
  AOI22_X1 U5414 ( .A1(n8292), .A2(n34162), .B1(n8291), .B2(n34161), .ZN(
        n34074) );
  AOI22_X1 U5415 ( .A1(n8290), .A2(n32677), .B1(n8289), .B2(n32674), .ZN(
        n34073) );
  NAND4_X1 U5416 ( .A1(n34076), .A2(n34075), .A3(n34074), .A4(n34073), .ZN(
        n34092) );
  AOI22_X1 U5417 ( .A1(n8288), .A2(n34170), .B1(n8287), .B2(n34169), .ZN(
        n34080) );
  AOI22_X1 U5418 ( .A1(n8286), .A2(n32680), .B1(n8285), .B2(n34171), .ZN(
        n34079) );
  AOI22_X1 U5419 ( .A1(n8284), .A2(n32679), .B1(n8283), .B2(n32673), .ZN(
        n34078) );
  AOI22_X1 U5420 ( .A1(n8282), .A2(n32719), .B1(n8281), .B2(n32672), .ZN(
        n34077) );
  NAND4_X1 U5421 ( .A1(n34080), .A2(n34079), .A3(n34078), .A4(n34077), .ZN(
        n34091) );
  AOI22_X1 U5422 ( .A1(n8280), .A2(n34182), .B1(n8279), .B2(n32671), .ZN(
        n34084) );
  AOI22_X1 U5423 ( .A1(n8278), .A2(n34184), .B1(n8277), .B2(n34183), .ZN(
        n34083) );
  AOI22_X1 U5424 ( .A1(n8276), .A2(n34186), .B1(n8275), .B2(n34185), .ZN(
        n34082) );
  AOI22_X1 U5425 ( .A1(n8274), .A2(n32682), .B1(n8273), .B2(n32670), .ZN(
        n34081) );
  NAND4_X1 U5426 ( .A1(n34084), .A2(n34083), .A3(n34082), .A4(n34081), .ZN(
        n34090) );
  AOI22_X1 U5427 ( .A1(n8272), .A2(n34194), .B1(n8271), .B2(n34193), .ZN(
        n34088) );
  AOI22_X1 U5428 ( .A1(n8270), .A2(n32681), .B1(n8269), .B2(n32669), .ZN(
        n34087) );
  AOI22_X1 U5429 ( .A1(n8268), .A2(n34198), .B1(n8267), .B2(n32668), .ZN(
        n34086) );
  AOI22_X1 U5430 ( .A1(n8266), .A2(n34200), .B1(n8265), .B2(n34199), .ZN(
        n34085) );
  NAND4_X1 U5431 ( .A1(n34088), .A2(n34087), .A3(n34086), .A4(n34085), .ZN(
        n34089) );
  NOR4_X1 U5432 ( .A1(n34092), .A2(n34091), .A3(n34090), .A4(n34089), .ZN(
        n34093) );
  OAI22_X1 U5433 ( .A1(n34093), .A2(n34210), .B1(n14151), .B2(n32722), .ZN(
        n5839) );
  AOI22_X1 U5434 ( .A1(n8328), .A2(n32716), .B1(n8327), .B2(n32676), .ZN(
        n34097) );
  AOI22_X1 U5435 ( .A1(n8326), .A2(n32678), .B1(n8325), .B2(n32675), .ZN(
        n34096) );
  AOI22_X1 U5436 ( .A1(n8324), .A2(n34162), .B1(n8323), .B2(n34161), .ZN(
        n34095) );
  AOI22_X1 U5437 ( .A1(n8322), .A2(n32677), .B1(n8321), .B2(n32674), .ZN(
        n34094) );
  NAND4_X1 U5438 ( .A1(n34097), .A2(n34096), .A3(n34095), .A4(n34094), .ZN(
        n34113) );
  AOI22_X1 U5439 ( .A1(n8320), .A2(n34170), .B1(n8319), .B2(n32717), .ZN(
        n34101) );
  AOI22_X1 U5440 ( .A1(n8318), .A2(n32680), .B1(n8317), .B2(n32718), .ZN(
        n34100) );
  AOI22_X1 U5441 ( .A1(n8316), .A2(n32679), .B1(n8315), .B2(n32673), .ZN(
        n34099) );
  AOI22_X1 U5442 ( .A1(n8314), .A2(n34176), .B1(n8313), .B2(n32672), .ZN(
        n34098) );
  NAND4_X1 U5443 ( .A1(n34101), .A2(n34100), .A3(n34099), .A4(n34098), .ZN(
        n34112) );
  AOI22_X1 U5444 ( .A1(n8312), .A2(n34182), .B1(n8311), .B2(n32671), .ZN(
        n34105) );
  AOI22_X1 U5445 ( .A1(n8310), .A2(n34184), .B1(n8309), .B2(n34183), .ZN(
        n34104) );
  AOI22_X1 U5446 ( .A1(n8308), .A2(n34186), .B1(n8307), .B2(n34185), .ZN(
        n34103) );
  AOI22_X1 U5447 ( .A1(n8306), .A2(n32682), .B1(n8305), .B2(n32670), .ZN(
        n34102) );
  NAND4_X1 U5448 ( .A1(n34105), .A2(n34104), .A3(n34103), .A4(n34102), .ZN(
        n34111) );
  AOI22_X1 U5449 ( .A1(n8304), .A2(n34194), .B1(n8303), .B2(n32720), .ZN(
        n34109) );
  AOI22_X1 U5450 ( .A1(n8302), .A2(n32681), .B1(n8301), .B2(n32669), .ZN(
        n34108) );
  AOI22_X1 U5451 ( .A1(n8300), .A2(n34198), .B1(n8299), .B2(n32668), .ZN(
        n34107) );
  AOI22_X1 U5452 ( .A1(n8298), .A2(n34200), .B1(n8297), .B2(n32721), .ZN(
        n34106) );
  NAND4_X1 U5453 ( .A1(n34109), .A2(n34108), .A3(n34107), .A4(n34106), .ZN(
        n34110) );
  NOR4_X1 U5454 ( .A1(n34113), .A2(n34112), .A3(n34111), .A4(n34110), .ZN(
        n34114) );
  OAI22_X1 U5455 ( .A1(n34114), .A2(n34210), .B1(n14152), .B2(n32722), .ZN(
        n5840) );
  AOI22_X1 U5456 ( .A1(n8360), .A2(n34158), .B1(n8359), .B2(n32676), .ZN(
        n34118) );
  AOI22_X1 U5457 ( .A1(n8358), .A2(n32678), .B1(n8357), .B2(n32675), .ZN(
        n34117) );
  AOI22_X1 U5458 ( .A1(n8356), .A2(n32667), .B1(n8355), .B2(n34161), .ZN(
        n34116) );
  AOI22_X1 U5459 ( .A1(n8354), .A2(n32677), .B1(n8353), .B2(n32674), .ZN(
        n34115) );
  NAND4_X1 U5460 ( .A1(n34118), .A2(n34117), .A3(n34116), .A4(n34115), .ZN(
        n34134) );
  AOI22_X1 U5461 ( .A1(n8352), .A2(n34170), .B1(n8351), .B2(n32717), .ZN(
        n34122) );
  AOI22_X1 U5462 ( .A1(n8350), .A2(n32680), .B1(n8349), .B2(n34171), .ZN(
        n34121) );
  AOI22_X1 U5463 ( .A1(n8348), .A2(n32679), .B1(n8347), .B2(n32673), .ZN(
        n34120) );
  AOI22_X1 U5464 ( .A1(n8346), .A2(n34176), .B1(n8345), .B2(n32672), .ZN(
        n34119) );
  NAND4_X1 U5465 ( .A1(n34122), .A2(n34121), .A3(n34120), .A4(n34119), .ZN(
        n34133) );
  AOI22_X1 U5466 ( .A1(n8344), .A2(n34182), .B1(n8343), .B2(n32671), .ZN(
        n34126) );
  AOI22_X1 U5467 ( .A1(n8342), .A2(n34184), .B1(n8341), .B2(n34183), .ZN(
        n34125) );
  AOI22_X1 U5468 ( .A1(n8340), .A2(n34186), .B1(n8339), .B2(n34185), .ZN(
        n34124) );
  AOI22_X1 U5469 ( .A1(n8338), .A2(n32682), .B1(n8337), .B2(n32670), .ZN(
        n34123) );
  NAND4_X1 U5470 ( .A1(n34126), .A2(n34125), .A3(n34124), .A4(n34123), .ZN(
        n34132) );
  AOI22_X1 U5471 ( .A1(n8336), .A2(n34194), .B1(n8335), .B2(n32720), .ZN(
        n34130) );
  AOI22_X1 U5472 ( .A1(n8334), .A2(n32681), .B1(n8333), .B2(n32669), .ZN(
        n34129) );
  AOI22_X1 U5473 ( .A1(n8332), .A2(n34198), .B1(n8331), .B2(n32668), .ZN(
        n34128) );
  AOI22_X1 U5474 ( .A1(n8330), .A2(n34200), .B1(n8329), .B2(n32721), .ZN(
        n34127) );
  NAND4_X1 U5475 ( .A1(n34130), .A2(n34129), .A3(n34128), .A4(n34127), .ZN(
        n34131) );
  NOR4_X1 U5476 ( .A1(n34134), .A2(n34133), .A3(n34132), .A4(n34131), .ZN(
        n34135) );
  OAI22_X1 U5477 ( .A1(n34135), .A2(n34210), .B1(n14153), .B2(n32722), .ZN(
        n5841) );
  AOI22_X1 U5478 ( .A1(n8392), .A2(n32716), .B1(n8391), .B2(n32676), .ZN(
        n34139) );
  AOI22_X1 U5479 ( .A1(n8390), .A2(n32678), .B1(n8389), .B2(n32675), .ZN(
        n34138) );
  AOI22_X1 U5480 ( .A1(n8388), .A2(n34162), .B1(n8387), .B2(n34161), .ZN(
        n34137) );
  AOI22_X1 U5481 ( .A1(n8386), .A2(n32677), .B1(n8385), .B2(n32674), .ZN(
        n34136) );
  NAND4_X1 U5482 ( .A1(n34139), .A2(n34138), .A3(n34137), .A4(n34136), .ZN(
        n34155) );
  AOI22_X1 U5483 ( .A1(n8384), .A2(n34170), .B1(n8383), .B2(n32717), .ZN(
        n34143) );
  AOI22_X1 U5484 ( .A1(n8382), .A2(n32680), .B1(n8381), .B2(n32718), .ZN(
        n34142) );
  AOI22_X1 U5485 ( .A1(n8380), .A2(n32679), .B1(n8379), .B2(n32673), .ZN(
        n34141) );
  AOI22_X1 U5486 ( .A1(n8378), .A2(n34176), .B1(n8377), .B2(n32672), .ZN(
        n34140) );
  NAND4_X1 U5487 ( .A1(n34143), .A2(n34142), .A3(n34141), .A4(n34140), .ZN(
        n34154) );
  AOI22_X1 U5488 ( .A1(n8376), .A2(n34182), .B1(n8375), .B2(n32671), .ZN(
        n34147) );
  AOI22_X1 U5489 ( .A1(n8374), .A2(n34184), .B1(n8373), .B2(n34183), .ZN(
        n34146) );
  AOI22_X1 U5490 ( .A1(n8372), .A2(n32666), .B1(n8371), .B2(n34185), .ZN(
        n34145) );
  AOI22_X1 U5491 ( .A1(n8370), .A2(n32682), .B1(n8369), .B2(n32670), .ZN(
        n34144) );
  NAND4_X1 U5492 ( .A1(n34147), .A2(n34146), .A3(n34145), .A4(n34144), .ZN(
        n34153) );
  AOI22_X1 U5493 ( .A1(n8368), .A2(n34194), .B1(n8367), .B2(n32720), .ZN(
        n34151) );
  AOI22_X1 U5494 ( .A1(n8366), .A2(n32681), .B1(n8365), .B2(n32669), .ZN(
        n34150) );
  AOI22_X1 U5495 ( .A1(n8364), .A2(n34198), .B1(n8363), .B2(n32668), .ZN(
        n34149) );
  AOI22_X1 U5496 ( .A1(n8362), .A2(n34200), .B1(n8361), .B2(n32721), .ZN(
        n34148) );
  NAND4_X1 U5497 ( .A1(n34151), .A2(n34150), .A3(n34149), .A4(n34148), .ZN(
        n34152) );
  NOR4_X1 U5498 ( .A1(n34155), .A2(n34154), .A3(n34153), .A4(n34152), .ZN(
        n34156) );
  OAI22_X1 U5499 ( .A1(n34156), .A2(n32665), .B1(n14154), .B2(n32722), .ZN(
        n5842) );
  AOI22_X1 U5500 ( .A1(n8424), .A2(n32716), .B1(n8423), .B2(n32676), .ZN(
        n34168) );
  AOI22_X1 U5501 ( .A1(n8422), .A2(n32678), .B1(n8421), .B2(n32675), .ZN(
        n34167) );
  AOI22_X1 U5502 ( .A1(n8420), .A2(n34162), .B1(n8419), .B2(n34161), .ZN(
        n34166) );
  AOI22_X1 U5503 ( .A1(n8418), .A2(n32677), .B1(n8417), .B2(n32674), .ZN(
        n34165) );
  NAND4_X1 U5504 ( .A1(n34168), .A2(n34167), .A3(n34166), .A4(n34165), .ZN(
        n34208) );
  AOI22_X1 U5505 ( .A1(n8416), .A2(n34170), .B1(n8415), .B2(n32717), .ZN(
        n34180) );
  AOI22_X1 U5506 ( .A1(n8414), .A2(n32680), .B1(n8413), .B2(n32718), .ZN(
        n34179) );
  AOI22_X1 U5507 ( .A1(n8412), .A2(n32679), .B1(n8411), .B2(n32673), .ZN(
        n34178) );
  AOI22_X1 U5508 ( .A1(n8410), .A2(n34176), .B1(n8409), .B2(n32672), .ZN(
        n34177) );
  NAND4_X1 U5509 ( .A1(n34180), .A2(n34179), .A3(n34178), .A4(n34177), .ZN(
        n34207) );
  AOI22_X1 U5510 ( .A1(n8408), .A2(n34182), .B1(n8407), .B2(n32671), .ZN(
        n34192) );
  AOI22_X1 U5511 ( .A1(n8406), .A2(n34184), .B1(n8405), .B2(n34183), .ZN(
        n34191) );
  AOI22_X1 U5512 ( .A1(n8404), .A2(n32666), .B1(n8403), .B2(n34185), .ZN(
        n34190) );
  AOI22_X1 U5513 ( .A1(n8402), .A2(n32682), .B1(n8401), .B2(n32670), .ZN(
        n34189) );
  NAND4_X1 U5514 ( .A1(n34192), .A2(n34191), .A3(n34190), .A4(n34189), .ZN(
        n34206) );
  AOI22_X1 U5515 ( .A1(n8400), .A2(n34194), .B1(n8399), .B2(n32720), .ZN(
        n34204) );
  AOI22_X1 U5516 ( .A1(n8398), .A2(n32681), .B1(n8397), .B2(n32669), .ZN(
        n34203) );
  AOI22_X1 U5517 ( .A1(n8396), .A2(n34198), .B1(n8395), .B2(n32668), .ZN(
        n34202) );
  AOI22_X1 U5518 ( .A1(n8394), .A2(n34200), .B1(n8393), .B2(n32721), .ZN(
        n34201) );
  NAND4_X1 U5519 ( .A1(n34204), .A2(n34203), .A3(n34202), .A4(n34201), .ZN(
        n34205) );
  NOR4_X1 U5520 ( .A1(n34208), .A2(n34207), .A3(n34206), .A4(n34205), .ZN(
        n34211) );
  OAI22_X1 U5521 ( .A1(n34211), .A2(n32665), .B1(n14155), .B2(n32722), .ZN(
        n5843) );
  NAND2_X1 U5522 ( .A1(EN), .A2(RD2), .ZN(n34212) );
  NAND2_X1 U5523 ( .A1(RST), .A2(n34212), .ZN(n5845) );
  INV_X1 U5524 ( .A(n34213), .ZN(n5913) );
endmodule


module SNPS_CLOCK_GATE_HIGH_DLX_WIDTH32_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net247640, n2, n3;
  assign net247640 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net247640), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_DLX_WIDTH32_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net247640, n2, n3;
  assign net247640 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net247640), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_DLX_WIDTH32_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net247640, n2, n3;
  assign net247640 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net247640), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_DLX_WIDTH32_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net247640, n2, n3;
  assign net247640 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net247640), .A2(TE), .ZN(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_DLX_WIDTH32_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net247640, n2, n3;
  assign net247640 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
  OR2_X1 U1 ( .A1(net247640), .A2(TE), .ZN(n3) );
endmodule


module DLX_WIDTH32 ( CLK, RST, IRAM_EN, IRAM_ADDR, IRAM_DATA, DRAM_EN, DRAM_RW, 
        DRAM_ADDR, DRAM_DATA_IN, DRAM_DATA_OUT );
  output [5:0] IRAM_ADDR;
  input [31:0] IRAM_DATA;
  output [5:0] DRAM_ADDR;
  input [31:0] DRAM_DATA_IN;
  output [31:0] DRAM_DATA_OUT;
  input CLK, RST;
  output IRAM_EN, DRAM_EN, DRAM_RW;
  wire   w_RF_RD1, w_RF_RD2, w_MuxIMM_SEL, w_SIGN_EN, w_MuxA_SEL, w_MuxB_SEL,
         w_EQ_COND, w_JUMP_EN, w_RF_WE3, w_RF_WE4, w_SIGN_LD_EN, w_RF_WE,
         \IR/n61 , \IR/n60 , \IR/n59 , \IR/n58 , \IR/n57 , \CU/n140 ,
         \CU/n139 , \CU/n138 , \CU/n142 , \CU/aluOpcodei[4] ,
         \CU/aluOpcodei[3] , \CU/aluOpcodei[2] , \CU/aluOpcodei[1] ,
         \CU/aluOpcodei[0] , \CU/cw[3] , \CU/cw[6] , \CU/cw[17] , \CU/cw[18] ,
         \CU/cw[20] , \CU/cw[21] , \CU/aluOpcode2[4] , \CU/aluOpcode2[3] ,
         \CU/aluOpcode2[2] , \CU/aluOpcode2[1] , \CU/aluOpcode2[0] ,
         \CU/aluOpcode1[4] , \CU/aluOpcode1[3] , \CU/aluOpcode1[2] ,
         \CU/aluOpcode1[1] , \CU/aluOpcode1[0] , \CU/cw4[2] , \CU/cw4[1] ,
         \CU/cw4[0] , \CU/cw3[7] , \CU/cw3[6] , \CU/cw3[5] , \CU/cw3[4] ,
         \CU/cw3[3] , \CU/cw3[2] , \CU/cw3[1] , \CU/cw3[0] , \CU/cw3_9 ,
         \CU/cw3_10 , \CU/cw3_11 , \CU/cw2[15] , \CU/cw2[14] , \CU/cw2[13] ,
         \CU/cw2[12] , \CU/cw2[11] , \CU/cw2[10] , \CU/cw2[9] , \CU/cw2[8] ,
         \CU/cw2[7] , \CU/cw2[6] , \CU/cw2[5] , \CU/cw2[4] , \CU/cw2[3] ,
         \CU/cw2[2] , \CU/cw2[1] , \CU/cw2[0] , \CU/cw1[20] , \CU/cw1[19] ,
         \CU/cw1[18] , \CU/cw1[17] , \CU/cw1[15] , \CU/cw1[14] , \CU/cw1[13] ,
         \CU/cw1[12] , \CU/cw1[11] , \CU/cw1[10] , \CU/cw1[9] , \CU/cw1[8] ,
         \CU/cw1[7] , \CU/cw1[6] , \CU/cw1[5] , \CU/cw1[4] , \CU/cw1[3] ,
         \CU/cw1[2] , \CU/cw1[1] , \CU/cw1[0] , \DP/IMMS26[25] ,
         \DP/IMMS26[24] , \DP/IMMS26[23] , \DP/IMMS26[22] , \DP/IMMS26[21] ,
         \DP/RD4[0] , \DP/RD4[1] , \DP/RD4[2] , \DP/RD4[3] , \DP/RD4[4] ,
         \DP/RegB_IN[31] , \DP/RegB_IN[30] , \DP/RegB_IN[29] ,
         \DP/RegB_IN[28] , \DP/RegB_IN[27] , \DP/RegB_IN[26] ,
         \DP/RegB_IN[25] , \DP/RegB_IN[24] , \DP/RegB_IN[23] ,
         \DP/RegB_IN[22] , \DP/RegB_IN[21] , \DP/RegB_IN[20] ,
         \DP/RegB_IN[19] , \DP/RegB_IN[18] , \DP/RegB_IN[17] ,
         \DP/RegB_IN[16] , \DP/RegB_IN[15] , \DP/RegB_IN[14] ,
         \DP/RegB_IN[13] , \DP/RegB_IN[12] , \DP/RegB_IN[11] ,
         \DP/RegB_IN[10] , \DP/RegB_IN[9] , \DP/RegB_IN[8] , \DP/RegB_IN[7] ,
         \DP/RegB_IN[6] , \DP/RegB_IN[5] , \DP/RegB_IN[4] , \DP/RegB_IN[3] ,
         \DP/RegB_IN[2] , \DP/RegB_IN[1] , \DP/RegB_IN[0] , \DP/RegA_IN[31] ,
         \DP/RegA_IN[30] , \DP/RegA_IN[29] , \DP/RegA_IN[28] ,
         \DP/RegA_IN[27] , \DP/RegA_IN[26] , \DP/RegA_IN[25] ,
         \DP/RegA_IN[24] , \DP/RegA_IN[23] , \DP/RegA_IN[22] ,
         \DP/RegA_IN[21] , \DP/RegA_IN[20] , \DP/RegA_IN[19] ,
         \DP/RegA_IN[18] , \DP/RegA_IN[17] , \DP/RegA_IN[16] ,
         \DP/RegA_IN[15] , \DP/RegA_IN[14] , \DP/RegA_IN[13] ,
         \DP/RegA_IN[12] , \DP/RegA_IN[11] , \DP/RegA_IN[10] , \DP/RegA_IN[9] ,
         \DP/RegA_IN[8] , \DP/RegA_IN[7] , \DP/RegA_IN[6] , \DP/RegA_IN[5] ,
         \DP/RegA_IN[4] , \DP/RegA_IN[3] , \DP/RegA_IN[2] , \DP/RegA_IN[1] ,
         \DP/RegA_IN[0] , \DP/NPC[1] , \DP/NPC[0] , \DP/RegRD2/n14 ,
         \DP/RegRD2/n13 , \DP/RegRD2/n12 , \DP/RegRD2/n11 , \DP/RegRD2/n10 ,
         \DP/RegRD2/n7 , \DP/ALU0/n109 , \DP/ALU0/n112 , \DP/ALU0/n114 ,
         \DP/ALU0/N27 , \DP/ALU0/N20 , \DP/ALU0/S_B_LHI[15] ,
         \DP/ALU0/S_B_LHI[14] , \DP/ALU0/S_B_LHI[13] , \DP/ALU0/S_B_LHI[12] ,
         \DP/ALU0/S_B_LHI[11] , \DP/ALU0/S_B_LHI[10] , \DP/ALU0/S_B_LHI[9] ,
         \DP/ALU0/S_B_LHI[8] , \DP/ALU0/S_B_LHI[7] , \DP/ALU0/S_B_LHI[6] ,
         \DP/ALU0/S_B_LHI[5] , \DP/ALU0/S_B_LHI[4] , \DP/ALU0/S_B_LHI[3] ,
         \DP/ALU0/S_B_LHI[2] , \DP/ALU0/S_B_LHI[1] , \DP/ALU0/S_B_LHI[0] ,
         \DP/ALU0/S_B_MULT[15] , \DP/ALU0/S_B_MULT[14] ,
         \DP/ALU0/S_B_MULT[13] , \DP/ALU0/S_B_MULT[12] ,
         \DP/ALU0/S_B_MULT[11] , \DP/ALU0/S_B_MULT[10] , \DP/ALU0/S_B_MULT[9] ,
         \DP/ALU0/S_B_MULT[8] , \DP/ALU0/S_B_MULT[7] , \DP/ALU0/S_B_MULT[6] ,
         \DP/ALU0/S_B_MULT[5] , \DP/ALU0/S_B_MULT[4] , \DP/ALU0/S_B_MULT[3] ,
         \DP/ALU0/S_B_MULT[2] , \DP/ALU0/S_B_MULT[1] , \DP/ALU0/S_B_MULT[0] ,
         \DP/ALU0/s_A_MULT[15] , \DP/ALU0/s_A_MULT[14] ,
         \DP/ALU0/s_A_MULT[13] , \DP/ALU0/s_A_MULT[12] ,
         \DP/ALU0/s_A_MULT[11] , \DP/ALU0/s_A_MULT[10] , \DP/ALU0/s_A_MULT[9] ,
         \DP/ALU0/s_A_MULT[8] , \DP/ALU0/s_A_MULT[7] , \DP/ALU0/s_A_MULT[6] ,
         \DP/ALU0/s_A_MULT[5] , \DP/ALU0/s_A_MULT[4] , \DP/ALU0/s_A_MULT[3] ,
         \DP/ALU0/s_A_MULT[2] , \DP/ALU0/s_A_MULT[1] , \DP/ALU0/s_A_MULT[0] ,
         \DP/ALU0/s_SHIFT[1] , \DP/ALU0/s_SHIFT[0] , \DP/ALU0/S_B_SHIFT[4] ,
         \DP/ALU0/S_B_SHIFT[3] , \DP/ALU0/S_B_SHIFT[2] ,
         \DP/ALU0/S_B_SHIFT[1] , \DP/ALU0/S_B_SHIFT[0] ,
         \DP/ALU0/s_A_SHIFT[31] , \DP/ALU0/s_A_SHIFT[30] ,
         \DP/ALU0/s_A_SHIFT[29] , \DP/ALU0/s_A_SHIFT[28] ,
         \DP/ALU0/s_A_SHIFT[27] , \DP/ALU0/s_A_SHIFT[26] ,
         \DP/ALU0/s_A_SHIFT[25] , \DP/ALU0/s_A_SHIFT[24] ,
         \DP/ALU0/s_A_SHIFT[23] , \DP/ALU0/s_A_SHIFT[22] ,
         \DP/ALU0/s_A_SHIFT[21] , \DP/ALU0/s_A_SHIFT[20] ,
         \DP/ALU0/s_A_SHIFT[19] , \DP/ALU0/s_A_SHIFT[18] ,
         \DP/ALU0/s_A_SHIFT[17] , \DP/ALU0/s_A_SHIFT[16] ,
         \DP/ALU0/s_A_SHIFT[15] , \DP/ALU0/s_A_SHIFT[14] ,
         \DP/ALU0/s_A_SHIFT[13] , \DP/ALU0/s_A_SHIFT[12] ,
         \DP/ALU0/s_A_SHIFT[11] , \DP/ALU0/s_A_SHIFT[10] ,
         \DP/ALU0/s_A_SHIFT[9] , \DP/ALU0/s_A_SHIFT[8] ,
         \DP/ALU0/s_A_SHIFT[7] , \DP/ALU0/s_A_SHIFT[6] ,
         \DP/ALU0/s_A_SHIFT[5] , \DP/ALU0/s_A_SHIFT[4] ,
         \DP/ALU0/s_A_SHIFT[3] , \DP/ALU0/s_A_SHIFT[2] ,
         \DP/ALU0/s_A_SHIFT[1] , \DP/ALU0/s_A_SHIFT[0] , \DP/ALU0/s_LOGIC[3] ,
         \DP/ALU0/s_LOGIC[2] , \DP/ALU0/S_B_LOGIC[31] ,
         \DP/ALU0/S_B_LOGIC[30] , \DP/ALU0/S_B_LOGIC[29] ,
         \DP/ALU0/S_B_LOGIC[28] , \DP/ALU0/S_B_LOGIC[27] ,
         \DP/ALU0/S_B_LOGIC[26] , \DP/ALU0/S_B_LOGIC[25] ,
         \DP/ALU0/S_B_LOGIC[24] , \DP/ALU0/S_B_LOGIC[23] ,
         \DP/ALU0/S_B_LOGIC[22] , \DP/ALU0/S_B_LOGIC[21] ,
         \DP/ALU0/S_B_LOGIC[20] , \DP/ALU0/S_B_LOGIC[19] ,
         \DP/ALU0/S_B_LOGIC[18] , \DP/ALU0/S_B_LOGIC[17] ,
         \DP/ALU0/S_B_LOGIC[16] , \DP/ALU0/S_B_LOGIC[15] ,
         \DP/ALU0/S_B_LOGIC[14] , \DP/ALU0/S_B_LOGIC[13] ,
         \DP/ALU0/S_B_LOGIC[12] , \DP/ALU0/S_B_LOGIC[11] ,
         \DP/ALU0/S_B_LOGIC[10] , \DP/ALU0/S_B_LOGIC[9] ,
         \DP/ALU0/S_B_LOGIC[8] , \DP/ALU0/S_B_LOGIC[7] ,
         \DP/ALU0/S_B_LOGIC[6] , \DP/ALU0/S_B_LOGIC[5] ,
         \DP/ALU0/S_B_LOGIC[4] , \DP/ALU0/S_B_LOGIC[3] ,
         \DP/ALU0/S_B_LOGIC[2] , \DP/ALU0/S_B_LOGIC[1] ,
         \DP/ALU0/S_B_LOGIC[0] , \DP/ALU0/s_A_LOGIC[31] ,
         \DP/ALU0/s_A_LOGIC[30] , \DP/ALU0/s_A_LOGIC[29] ,
         \DP/ALU0/s_A_LOGIC[28] , \DP/ALU0/s_A_LOGIC[27] ,
         \DP/ALU0/s_A_LOGIC[26] , \DP/ALU0/s_A_LOGIC[25] ,
         \DP/ALU0/s_A_LOGIC[24] , \DP/ALU0/s_A_LOGIC[23] ,
         \DP/ALU0/s_A_LOGIC[22] , \DP/ALU0/s_A_LOGIC[21] ,
         \DP/ALU0/s_A_LOGIC[20] , \DP/ALU0/s_A_LOGIC[19] ,
         \DP/ALU0/s_A_LOGIC[18] , \DP/ALU0/s_A_LOGIC[17] ,
         \DP/ALU0/s_A_LOGIC[16] , \DP/ALU0/s_A_LOGIC[15] ,
         \DP/ALU0/s_A_LOGIC[14] , \DP/ALU0/s_A_LOGIC[13] ,
         \DP/ALU0/s_A_LOGIC[12] , \DP/ALU0/s_A_LOGIC[11] ,
         \DP/ALU0/s_A_LOGIC[10] , \DP/ALU0/s_A_LOGIC[9] ,
         \DP/ALU0/s_A_LOGIC[8] , \DP/ALU0/s_A_LOGIC[7] ,
         \DP/ALU0/s_A_LOGIC[6] , \DP/ALU0/s_A_LOGIC[5] ,
         \DP/ALU0/s_A_LOGIC[4] , \DP/ALU0/s_A_LOGIC[3] ,
         \DP/ALU0/s_A_LOGIC[2] , \DP/ALU0/s_A_LOGIC[1] ,
         \DP/ALU0/s_A_LOGIC[0] , \DP/ALU0/s_ADD_SUB , \DP/ALU0/S_B_ADDER[31] ,
         \DP/ALU0/S_B_ADDER[30] , \DP/ALU0/S_B_ADDER[29] ,
         \DP/ALU0/S_B_ADDER[28] , \DP/ALU0/S_B_ADDER[27] ,
         \DP/ALU0/S_B_ADDER[26] , \DP/ALU0/S_B_ADDER[25] ,
         \DP/ALU0/S_B_ADDER[24] , \DP/ALU0/S_B_ADDER[23] ,
         \DP/ALU0/S_B_ADDER[22] , \DP/ALU0/S_B_ADDER[21] ,
         \DP/ALU0/S_B_ADDER[20] , \DP/ALU0/S_B_ADDER[19] ,
         \DP/ALU0/S_B_ADDER[18] , \DP/ALU0/S_B_ADDER[17] ,
         \DP/ALU0/S_B_ADDER[16] , \DP/ALU0/S_B_ADDER[15] ,
         \DP/ALU0/S_B_ADDER[14] , \DP/ALU0/S_B_ADDER[13] ,
         \DP/ALU0/S_B_ADDER[12] , \DP/ALU0/S_B_ADDER[11] ,
         \DP/ALU0/S_B_ADDER[10] , \DP/ALU0/S_B_ADDER[9] ,
         \DP/ALU0/S_B_ADDER[8] , \DP/ALU0/S_B_ADDER[7] ,
         \DP/ALU0/S_B_ADDER[6] , \DP/ALU0/S_B_ADDER[5] ,
         \DP/ALU0/S_B_ADDER[4] , \DP/ALU0/S_B_ADDER[3] ,
         \DP/ALU0/S_B_ADDER[2] , \DP/ALU0/S_B_ADDER[1] ,
         \DP/ALU0/S_B_ADDER[0] , \DP/ALU0/s_A_ADDER[31] ,
         \DP/ALU0/s_A_ADDER[30] , \DP/ALU0/s_A_ADDER[29] ,
         \DP/ALU0/s_A_ADDER[28] , \DP/ALU0/s_A_ADDER[27] ,
         \DP/ALU0/s_A_ADDER[26] , \DP/ALU0/s_A_ADDER[25] ,
         \DP/ALU0/s_A_ADDER[24] , \DP/ALU0/s_A_ADDER[23] ,
         \DP/ALU0/s_A_ADDER[22] , \DP/ALU0/s_A_ADDER[21] ,
         \DP/ALU0/s_A_ADDER[20] , \DP/ALU0/s_A_ADDER[19] ,
         \DP/ALU0/s_A_ADDER[18] , \DP/ALU0/s_A_ADDER[17] ,
         \DP/ALU0/s_A_ADDER[16] , \DP/ALU0/s_A_ADDER[15] ,
         \DP/ALU0/s_A_ADDER[14] , \DP/ALU0/s_A_ADDER[13] ,
         \DP/ALU0/s_A_ADDER[12] , \DP/ALU0/s_A_ADDER[11] ,
         \DP/ALU0/s_A_ADDER[10] , \DP/ALU0/s_A_ADDER[9] ,
         \DP/ALU0/s_A_ADDER[8] , \DP/ALU0/s_A_ADDER[7] ,
         \DP/ALU0/s_A_ADDER[6] , \DP/ALU0/s_A_ADDER[5] ,
         \DP/ALU0/s_A_ADDER[4] , \DP/ALU0/s_A_ADDER[3] ,
         \DP/ALU0/s_A_ADDER[2] , \DP/ALU0/s_A_ADDER[1] ,
         \DP/ALU0/s_A_ADDER[0] , \DP/ALU0/s_SIGN , \DP/RegALU3/n97 ,
         \DP/RegALU3/n96 , \DP/RegALU3/n94 , \DP/RegALU3/n93 ,
         \DP/RegALU3/n92 , \DP/RegALU3/n91 , \DP/RegALU3/n90 ,
         \DP/RegALU3/n89 , \DP/RegALU3/n88 , \DP/RegALU3/n87 ,
         \DP/RegALU3/n86 , \DP/RegALU3/n85 , \DP/RegALU3/n84 ,
         \DP/RegALU3/n83 , \DP/RegALU3/n82 , \DP/RegALU3/n81 ,
         \DP/RegALU3/n80 , \DP/RegALU3/n79 , \DP/RegALU3/n78 ,
         \DP/RegALU3/n77 , \DP/RegALU3/n76 , \DP/RegALU3/n75 ,
         \DP/RegALU3/n74 , \DP/RegALU3/n73 , \DP/RegALU3/n72 ,
         \DP/RegALU3/n71 , \DP/RegALU3/n70 , \DP/RegALU3/n69 ,
         \DP/RegALU3/n68 , \DP/RegRD3/n14 , \DP/RegRD3/n13 , \DP/RegRD3/n12 ,
         \DP/RegRD3/n11 , \DP/RegRD3/n10 , \DP/RegRD4/n14 , \DP/RegRD4/n13 ,
         \DP/RegRD4/n12 , \DP/RegRD4/n11 , \DP/RegRD4/n10 , \DP/RegRD4/n7 ,
         n897, n1176, n3015, n3018, n3019, n3020, n3021, n3022, n3024, n3025,
         n3026, n3027, n3028, n3029, n3032, n3033, n3034, n3036, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3061, n3062, n3064, n3065, n3067, n3068, n3070, n3071, n3073, n3074,
         n3076, n3077, n3079, n3080, n3082, n3083, n3085, n3086, n3088, n3089,
         n3091, n3092, n3094, n3095, n3098, n3099, n3101, n3102, n3104, n3105,
         n3107, n3108, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, \intadd_0/B[26] , \intadd_0/B[25] , \intadd_0/B[24] ,
         \intadd_0/B[23] , \intadd_0/B[22] , \intadd_0/B[21] ,
         \intadd_0/B[20] , \intadd_0/B[19] , \intadd_0/B[18] ,
         \intadd_0/B[17] , \intadd_0/B[16] , \intadd_0/B[15] ,
         \intadd_0/B[14] , \intadd_0/B[13] , \intadd_0/B[12] ,
         \intadd_0/B[11] , \intadd_0/B[10] , \intadd_0/B[9] , \intadd_0/B[8] ,
         \intadd_0/B[7] , \intadd_0/B[6] , \intadd_0/B[5] , \intadd_0/B[4] ,
         \intadd_0/B[3] , \intadd_0/B[2] , \intadd_0/B[1] , \intadd_0/B[0] ,
         \intadd_0/CI , \intadd_0/SUM[26] , \intadd_0/SUM[25] ,
         \intadd_0/SUM[24] , \intadd_0/SUM[23] , \intadd_0/SUM[22] ,
         \intadd_0/SUM[21] , \intadd_0/SUM[20] , \intadd_0/SUM[19] ,
         \intadd_0/SUM[18] , \intadd_0/SUM[17] , \intadd_0/SUM[16] ,
         \intadd_0/SUM[15] , \intadd_0/SUM[14] , \intadd_0/SUM[13] ,
         \intadd_0/SUM[12] , \intadd_0/SUM[11] , \intadd_0/SUM[10] ,
         \intadd_0/SUM[9] , \intadd_0/SUM[8] , \intadd_0/SUM[7] ,
         \intadd_0/SUM[6] , \intadd_0/SUM[5] , \intadd_0/SUM[4] ,
         \intadd_0/SUM[3] , \intadd_0/SUM[2] , \intadd_0/SUM[1] ,
         \intadd_0/SUM[0] , \intadd_0/n27 , \intadd_0/n26 , \intadd_0/n25 ,
         \intadd_0/n24 , \intadd_0/n23 , \intadd_0/n22 , \intadd_0/n21 ,
         \intadd_0/n20 , \intadd_0/n19 , \intadd_0/n18 , \intadd_0/n17 ,
         \intadd_0/n16 , \intadd_0/n15 , \intadd_0/n14 , \intadd_0/n13 ,
         \intadd_0/n12 , \intadd_0/n11 , \intadd_0/n10 , \intadd_0/n9 ,
         \intadd_0/n8 , \intadd_0/n7 , \intadd_0/n6 , \intadd_0/n5 ,
         \intadd_0/n4 , \intadd_0/n3 , \intadd_0/n2 , \intadd_0/n1 ,
         \intadd_1/A[12] , \intadd_1/A[11] , \intadd_1/A[0] , \intadd_1/B[12] ,
         \intadd_1/B[11] , \intadd_1/B[10] , \intadd_1/B[9] , \intadd_1/B[8] ,
         \intadd_1/B[7] , \intadd_1/B[6] , \intadd_1/B[5] , \intadd_1/B[4] ,
         \intadd_1/B[3] , \intadd_1/B[2] , \intadd_1/B[1] , \intadd_1/CI ,
         \intadd_1/SUM[12] , \intadd_1/SUM[11] , \intadd_1/SUM[10] ,
         \intadd_1/SUM[9] , \intadd_1/SUM[8] , \intadd_1/SUM[7] ,
         \intadd_1/SUM[6] , \intadd_1/SUM[5] , \intadd_1/SUM[4] ,
         \intadd_1/SUM[3] , \intadd_1/SUM[2] , \intadd_1/SUM[1] ,
         \intadd_1/SUM[0] , \intadd_1/n13 , \intadd_1/n12 , \intadd_1/n11 ,
         \intadd_1/n10 , \intadd_1/n9 , \intadd_1/n8 , \intadd_1/n7 ,
         \intadd_1/n6 , \intadd_1/n5 , \intadd_1/n4 , \intadd_1/n3 ,
         \intadd_1/n2 , \intadd_1/n1 , \intadd_2/A[12] , \intadd_2/A[11] ,
         \intadd_2/A[10] , \intadd_2/A[9] , \intadd_2/A[8] , \intadd_2/A[7] ,
         \intadd_2/A[6] , \intadd_2/A[5] , \intadd_2/A[4] , \intadd_2/A[3] ,
         \intadd_2/A[2] , \intadd_2/A[1] , \intadd_2/A[0] , \intadd_2/B[12] ,
         \intadd_2/B[11] , \intadd_2/B[10] , \intadd_2/B[9] , \intadd_2/B[8] ,
         \intadd_2/B[7] , \intadd_2/B[6] , \intadd_2/B[5] , \intadd_2/B[4] ,
         \intadd_2/B[3] , \intadd_2/B[2] , \intadd_2/B[1] , \intadd_2/B[0] ,
         \intadd_2/CI , \intadd_2/SUM[12] , \intadd_2/SUM[11] ,
         \intadd_2/SUM[10] , \intadd_2/SUM[9] , \intadd_2/SUM[8] ,
         \intadd_2/SUM[7] , \intadd_2/SUM[6] , \intadd_2/SUM[5] ,
         \intadd_2/SUM[4] , \intadd_2/SUM[3] , \intadd_2/SUM[2] ,
         \intadd_2/SUM[1] , \intadd_2/SUM[0] , \intadd_2/n13 , \intadd_2/n12 ,
         \intadd_2/n11 , \intadd_2/n10 , \intadd_2/n9 , \intadd_2/n8 ,
         \intadd_2/n7 , \intadd_2/n6 , \intadd_2/n5 , \intadd_2/n4 ,
         \intadd_2/n3 , \intadd_2/n2 , \intadd_2/n1 , \intadd_3/A[12] ,
         \intadd_3/A[11] , \intadd_3/A[10] , \intadd_3/A[9] , \intadd_3/A[8] ,
         \intadd_3/A[7] , \intadd_3/A[6] , \intadd_3/A[5] , \intadd_3/A[4] ,
         \intadd_3/A[3] , \intadd_3/A[2] , \intadd_3/A[1] , \intadd_3/A[0] ,
         \intadd_3/B[12] , \intadd_3/B[11] , \intadd_3/B[0] ,
         \intadd_3/SUM[1] , \intadd_3/SUM[0] , \intadd_3/n13 , \intadd_3/n12 ,
         \intadd_3/n11 , \intadd_3/n10 , \intadd_3/n9 , \intadd_3/n8 ,
         \intadd_3/n7 , \intadd_3/n6 , \intadd_3/n5 , \intadd_3/n4 ,
         \intadd_3/n3 , \intadd_3/n2 , \intadd_3/n1 , \intadd_4/A[12] ,
         \intadd_4/A[11] , \intadd_4/A[0] , \intadd_4/B[12] , \intadd_4/B[11] ,
         \intadd_4/B[10] , \intadd_4/B[9] , \intadd_4/B[8] , \intadd_4/B[7] ,
         \intadd_4/B[6] , \intadd_4/B[5] , \intadd_4/B[4] , \intadd_4/B[3] ,
         \intadd_4/B[2] , \intadd_4/B[1] , \intadd_4/CI , \intadd_4/SUM[12] ,
         \intadd_4/SUM[11] , \intadd_4/SUM[10] , \intadd_4/SUM[9] ,
         \intadd_4/SUM[8] , \intadd_4/SUM[7] , \intadd_4/SUM[6] ,
         \intadd_4/SUM[5] , \intadd_4/SUM[4] , \intadd_4/SUM[3] ,
         \intadd_4/SUM[2] , \intadd_4/SUM[1] , \intadd_4/SUM[0] ,
         \intadd_4/n13 , \intadd_4/n12 , \intadd_4/n11 , \intadd_4/n10 ,
         \intadd_4/n9 , \intadd_4/n8 , \intadd_4/n7 , \intadd_4/n6 ,
         \intadd_4/n5 , \intadd_4/n4 , \intadd_4/n3 , \intadd_4/n2 ,
         \intadd_4/n1 , \intadd_5/A[12] , \intadd_5/A[11] , \intadd_5/A[10] ,
         \intadd_5/A[9] , \intadd_5/A[8] , \intadd_5/A[7] , \intadd_5/A[6] ,
         \intadd_5/A[5] , \intadd_5/A[4] , \intadd_5/A[3] , \intadd_5/A[2] ,
         \intadd_5/A[1] , \intadd_5/A[0] , \intadd_5/B[12] , \intadd_5/B[0] ,
         \intadd_5/SUM[12] , \intadd_5/SUM[11] , \intadd_5/SUM[10] ,
         \intadd_5/SUM[9] , \intadd_5/SUM[8] , \intadd_5/SUM[7] ,
         \intadd_5/SUM[6] , \intadd_5/SUM[5] , \intadd_5/SUM[4] ,
         \intadd_5/SUM[3] , \intadd_5/SUM[2] , \intadd_5/SUM[1] ,
         \intadd_5/SUM[0] , \intadd_5/n13 , \intadd_5/n12 , \intadd_5/n11 ,
         \intadd_5/n10 , \intadd_5/n9 , \intadd_5/n8 , \intadd_5/n7 ,
         \intadd_5/n6 , \intadd_5/n5 , \intadd_5/n4 , \intadd_5/n3 ,
         \intadd_5/n2 , \intadd_5/n1 , \intadd_6/A[12] , \intadd_6/A[11] ,
         \intadd_6/A[0] , \intadd_6/B[12] , \intadd_6/B[11] , \intadd_6/B[10] ,
         \intadd_6/B[9] , \intadd_6/B[8] , \intadd_6/B[7] , \intadd_6/B[6] ,
         \intadd_6/B[5] , \intadd_6/B[4] , \intadd_6/B[3] , \intadd_6/B[2] ,
         \intadd_6/B[1] , \intadd_6/CI , \intadd_6/SUM[12] ,
         \intadd_6/SUM[11] , \intadd_6/SUM[10] , \intadd_6/SUM[9] ,
         \intadd_6/SUM[8] , \intadd_6/SUM[7] , \intadd_6/SUM[6] ,
         \intadd_6/SUM[5] , \intadd_6/SUM[4] , \intadd_6/SUM[3] ,
         \intadd_6/SUM[2] , \intadd_6/SUM[1] , \intadd_6/SUM[0] ,
         \intadd_6/n13 , \intadd_6/n12 , \intadd_6/n11 , \intadd_6/n10 ,
         \intadd_6/n9 , \intadd_6/n8 , \intadd_6/n7 , \intadd_6/n6 ,
         \intadd_6/n5 , \intadd_6/n4 , \intadd_6/n3 , \intadd_6/n2 ,
         \intadd_6/n1 , \intadd_7/A[12] , \intadd_7/A[11] , \intadd_7/A[10] ,
         \intadd_7/A[9] , \intadd_7/A[8] , \intadd_7/A[7] , \intadd_7/A[6] ,
         \intadd_7/A[5] , \intadd_7/A[4] , \intadd_7/A[3] , \intadd_7/A[2] ,
         \intadd_7/A[1] , \intadd_7/A[0] , \intadd_7/B[12] , \intadd_7/B[11] ,
         \intadd_7/B[10] , \intadd_7/B[9] , \intadd_7/B[8] , \intadd_7/B[7] ,
         \intadd_7/B[6] , \intadd_7/B[5] , \intadd_7/B[4] , \intadd_7/B[3] ,
         \intadd_7/B[2] , \intadd_7/B[1] , \intadd_7/B[0] , \intadd_7/CI ,
         \intadd_7/SUM[12] , \intadd_7/SUM[11] , \intadd_7/SUM[10] ,
         \intadd_7/SUM[9] , \intadd_7/SUM[8] , \intadd_7/SUM[7] ,
         \intadd_7/SUM[6] , \intadd_7/SUM[5] , \intadd_7/SUM[4] ,
         \intadd_7/SUM[3] , \intadd_7/SUM[2] , \intadd_7/SUM[1] ,
         \intadd_7/SUM[0] , \intadd_7/n13 , \intadd_7/n12 , \intadd_7/n11 ,
         \intadd_7/n10 , \intadd_7/n9 , \intadd_7/n8 , \intadd_7/n7 ,
         \intadd_7/n6 , \intadd_7/n5 , \intadd_7/n4 , \intadd_7/n3 ,
         \intadd_7/n2 , \intadd_7/n1 , n3190, n3191, n3214, n3247, n3248,
         n3249, n3253, n3254, n3260, n3270, n3273, n4923, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5158,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5402, n5463, n7226, n7227, n7228, n7229,
         n7230, n7286, n7478, n7489, \intadd_8/B[3] , \intadd_8/B[2] ,
         \intadd_8/B[1] , \intadd_8/CI , \intadd_8/SUM[3] , \intadd_8/SUM[2] ,
         \intadd_8/SUM[1] , \intadd_8/SUM[0] , \intadd_8/n4 , \intadd_8/n3 ,
         \intadd_8/n2 , \intadd_8/n1 , n7564, n7616, n7617, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7660, n7661, n7662, n7663, n7667,
         n7676, n7679, n9277, n9315, n18754, n19108, n20899, n22592, n26670,
         n32415, n32429, n37948, n40059, n40060, n40065, n43886, n43968,
         n43969, n45959, n47726, n47727, n49659, n49781, n49808, n49809,
         n49810, n49811, n49814, n49815, n49819, n49832, n49834, n49838,
         n49839, n49842, n49843, n49844, n49845, n49849, n49853, n49857,
         n49866, n49869, n49872, n49907, n49908, n49909, n49913, n49917,
         n49937, n49938, n49939, n49940, n49942, n49951, n49952, n49955,
         n49958, n51524, n51525, n51527, n51529, n51531, n51532, n51533,
         n51535, n51536, n51537, n51572, n51619, n51623, n51641, n51642,
         n51643, n51644, n51646, n51647, n51648, n51649, n51651, n51652,
         n51653, n51654, n51655, n51656, n51658, n51659, n51660, n51661,
         n51662, n51663, n51664, n51665, n51666, n51667, n51668, n51669,
         n51670, n51671, n51672, n51673, n51674, n51675, n51676, n51677,
         n51678, n51680, n51681, n51682, n51683, n51684, n51685, n51686,
         n51687, n51688, n51689, n51690, n51691, n51692, n51693, n51694,
         n51695, n51696, n51697, n51698, n51699, n51773, n51774, n51775,
         n51776, n51777, n51778, n51779, n51780, n51781, n51782, n51783,
         n51784, n51785, n51786, n51787, n51788, n51789, n51790, n51791,
         n51792, n51793, n51794, n51795, n51796, n51797, n51798, n51799,
         n51800, n51801, n51802, n51803, n53259, n53260, n53261, n53262,
         n53263, n53264, n53265, n53266, n53267, n53268, n53269, n53270,
         n53271, n53272, n53273, n53274, n53275, n53276, n53277, n53278,
         n53279, n53280, n53281, n53282, n53283, n53284, n53285, n53286,
         n53287, n53288, n53289, n53290, n53291, n53292, n53293, n53294,
         n53295, n53296, n53297, n53298, n53299, n53300, n53301, n53302,
         n53303, n53304, n53305, n53306, n53307, n53308, n53309, n53310,
         n53311, n53312, n53313, n53314, n53315, n53316, n53317, n53318,
         n53319, n53320, n53321, n53322, n53323, n53324, n53325, n53326,
         n53327, n53328, n53329, n53330, n53331, n53332, n53333, n53334,
         n53335, n53336, n53337, n53338, n53339, n53340, n53341, n53342,
         n53343, n53344, n53345, n53346, n53347, n53348, n53349, n53350,
         n53351, n53352, n53353, n53354, n53355, n53356, n53357, n53358,
         n53359, n53360, n53361, n53362, n53363, n53364, n53365, n53366,
         n53367, n53368, n53369, n53370, n53371, n53372, n53373, n53374,
         n53375, n53376, n53377, n53378, n53379, n53380, n53381, n53382,
         n53383, n53384, n53385, n53386, n53387, n53388, n53389, n53390,
         n53391, n53392, n53393, n53394, n53395, n53396, n53397, n53398,
         n53399, n53400, n53401, n53402, n53403, n53404, n53405, n53406,
         n53407, n53408, n53409, n53410, n53411, n53412, n53413, n53414,
         n53419, n53420, n53421, n53422, n53423, n53424, n53425, n53426,
         n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434,
         n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442,
         n53443, n53444, n53445, n53446, n53447, n53448, n53449, n53450,
         n53451, n53452, n53453, n53454, n53455, n53456, n53457, n53458,
         n53459, n53460, n53461, n53462, n53463, n53464, n53465, n53466,
         n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474,
         n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482,
         n53483, n53484, n53485, n53486, n53487, n53488, n53489, n53490,
         n53491, n53492, n53493, n53494, n53495, n53496, n53497, n53498,
         n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506,
         n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514,
         n53515, n53548, n53549, n53550, n53551, n53552, n53553, n53554,
         n53555, n53556, n53557, n53558, n53559, n53560, n53561, n53562,
         n53563, n53564, n53565, n53566, n53567, n53568, n53569, n53570,
         n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578,
         n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586,
         n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594,
         n53595, n53596, n53601, n53603, n53604, n53605, n53606, n53607,
         n53608, n53609, n53610, n53611, n53612, n53613, n53614, n53615,
         n53616, n53617, n53618, n53619, n53620, n53621, n53622, n53623,
         n53624, n53625, n53626, n53627, n53628, n53630, n53631, n53632,
         n53633, n53634, n53635, n53637, n53638, n53639, n53640, n53641,
         n53642, n53643, n53644, n53645, n53646, n53647, n53648, n53649,
         n53650, n53651, n53652, n53653, n53654, n53655, n53656, n53657,
         n53658, n53659, n53660, n53661, n53662, n53663, n53664, n53665,
         n53666, n53667, n53668, n53669, n53670, n53671, n53672, n53673,
         n53674, n53675, n53676, n53677, n53678, n53679, n53680, n53681,
         n53682, n53683, n53684, n53685, n53686, n53687, n53688, n53689,
         n53690, n53691, n53692, n53693, n53694, n53695, n53696, n53697,
         n53698, n53699, n53700, n53701, n53702, n53703, n53704, n53705,
         n53706, n53707, n53708, n53709, n53710, n53711, n53712, n53713,
         n53714, n53715, n53716, n53717, n53718, n53719, n53720, n53721,
         n53722, n53723, n53724, n53725, n53726, n53727, n53728, n53729,
         n53730, n53731, n53732, n53733, n53734, n53735, n53736, n53737,
         n53738, n53739, n53740, n53741, n53742, n53743, n53744, n53745,
         n53746, n53747, n53748, n53749, n53750, n53751, n53752, n53753,
         n53754, n53755, n53756, n53757, n53758, n53759, n53760, n53761,
         n53762, n53763, n53764, n53765, n53766, n53767, n53768, n53769,
         n53770, n53771, n53772, n53773, n53774, n53775, n53776, n53777,
         n53778, n53779, n53780, n53781, n53782, n53783, n53784, n53785,
         n53786, n53787, n53788, n53789, n53790, n53791, n53792, n53793,
         n53794, n53795, n53796, n53797, n53798, n53799, n53800, n53801,
         n53802, n53803, n53804, n53805, n53806, n53807, n53808, n53809,
         n53810, n53811, n53812, n53813, n53814, n53815, n53816, n53817,
         n53818, n53819, n53820, n53821, n53822, n53823, n53824, n53825,
         n53826, n53827, n53828, n53829, n53830, n53831, n53832, n53833,
         n53834, n53835, n53836, n53837, n53838, n53839, n53840, n53841,
         n53842, n53843, n53844, n53845, n53846, n53847, n53848, n53849,
         n53850, n53851, n53852, n53853, n53854, n53855, n53856, n53857,
         n53858, n53859, n53860, n53861, n53862, n53863, n53864, n53865,
         n53866, n53867, n53868, n53869, n53870, n53871, n53872, n53873,
         n53874, n53875, n53876, n53877, n53878, n53879, n53880, n53881,
         n53882, n53883, n53884, n53885, n53886, n53887, n53888, n53889,
         n53890, n53891, n53892, n53893, n53894, n53895, n53896, n53897,
         n53898, n53899, n53900, n53901, n53902, n53903, n53904, n53905,
         n53906, n53907, n53908, n53909, n53910, n53911, n53912, n53913,
         n53914, n53915, n53916, n53917, n53918, n53919, n53920, n53921,
         n53922, n53923, n53924, n53925, n53926, n53927, n53928, n53929,
         n53930, n53931, n53932, n53933, n53934, n53935, n53936, n53937,
         n53938, n53939, n53940, n53941, n53942, n53943, n53944, n53945,
         n53946, n53947, n53948, n53949, n53950, n53951, n53952, n53953,
         n53954, n53955, n53956, n53957, n53958, n53959, n53960, n53961,
         n53962, n53963, n53964, n53965, n53966, n53967, n53968, n53969,
         n53970, n53971, n53972, n53973, n53974, n53975, n53976, n53977,
         n53978, n53979, n53980, n53981, n53982, n53983, n53984, n53985,
         n53986, n53987, n53988, n53989, n53990, n53991, n53992, n53993,
         n53994, n53995, n53996, n53997, n53998, n53999, n54000, n54001,
         n54002, n54003, n54004, n54005, n54006, n54007, n54008, n54009,
         n54010, n54011, n54012, n54013, n54014, n54015, n54016, n54017,
         n54018, n54019, n54020, n54021, n54022, n54023, n54024, n54025,
         n54026, n54027, n54028, n54029, n54030, n54031, n54032, n54033,
         n54034, n54035, n54036, n54037, n54038, n54039, n54040, n54041,
         n54042, n54043, n54044, n54045, n54046, n54047, n54048, n54049,
         n54050, n54051, n54052, n54053, n54054, n54055, n54056, n54057,
         n54058, n54059, n54060, n54061, n54062, n54063, n54064, n54065,
         n54066, n54067, n54068, n54069, n54070, n54071, n54072, n54073,
         n54074, n54075, n54076, n54077, n54078, n54079, n54080, n54081,
         n54082, n54083, n54084, n54085, n54086, n54087, n54088, n54089,
         n54090, n54091, n54092, n54093, n54094, n54095, n54096, n54097,
         n54098, n54099, n54100, n54101, n54102, n54103, n54104, n54105,
         n54106, n54107, n54108, n54109, n54110, n54111, n54112, n54113,
         n54114, n54115, n54116, n54117, n54118, n54119, n54120, n54121,
         n54122, n54123, n54124, n54125, n54126, n54127, n54128, n54129,
         n54130, n54131, n54132, n54133, n54134, n54135, n54136, n54137,
         n54138, n54139, n54140, n54141, n54142, n54143, n54144, n54145,
         n54146, n54147, n54148, n54149, n54150, n54151, n54152, n54153,
         n54154, n54155, n54156, n54157, n54158, n54159, n54160, n54161,
         n54162, n54163, n54164, n54165, n54166, n54167, n54168, n54169,
         n54170, n54171, n54172, n54173, n54174, n54175, n54176, n54177,
         n54178, n54179, n54180, n54181, n54182, n54183, n54184, n54185,
         n54186, n54187, n54188, n54189, n54190, n54191, n54192, n54193,
         n54194, n54195, n54196, n54197, n54198, n54199, n54200, n54201,
         n54202, n54203, n54204, n54205, n54206, n54207, n54208, n54209,
         n54210, n54211, n54212, n54213, n54214, n54215, n54216, n54217,
         n54218, n54219, n54220, n54221, n54222, n54223, n54224, n54225,
         n54226, n54227, n54228, n54229, n54230, n54231, n54232, n54233,
         n54234, n54235, n54236, n54237, n54238, n54239, n54240, n54241,
         n54242, n54243, n54244, n54245, n54246, n54247, n54248, n54249,
         n54250, n54251, n54252, n54253, n54254, n54255, n54256, n54257,
         n54258, n54259, n54260, n54261, n54262, n54263, n54264, n54265,
         n54266, n54267, n54268, n54269, n54270, n54271, n54272, n54273,
         n54274, n54275, n54276, n54277, n54278, n54279, n54280, n54281,
         n54282, n54283, n54284, n54285, n54286, n54287, n54288, n54289,
         n54290, n54291, n54292, n54293, n54294, n54295, n54296, n54297,
         n54298, n54299, n54300, n54301, n54302, n54303, n54304, n54305,
         n54306, n54307, n54308, n54309, n54310, n54311, n54312, n54313,
         n54314, n54315, n54316, n54317, n54318, n54319, n54320, n54321,
         n54322, n54323, n54324, n54325, n54326, n54327, n54328, n54329,
         n54330, n54331, n54332, n54333, n54334, n54335, n54336, n54337,
         n54338, n54339, n54340, n54341, n54342, n54343, n54344, n54345,
         n54346, n54347, n54348, n54349, n54350, n54351, n54352, n54353,
         n54354, n54355, n54356, n54357, n54358, n54359, n54360, n54361,
         n54362, n54363, n54364, n54365, n54366, n54367, n54368, n54369,
         n54370, n54371, n54372, n54373, n54374, n54375, n54376, n54377,
         n54378, n54379, n54380, n54381, n54382, n54383, n54384, n54385,
         n54386, n54387, n54388, n54389, n54390, n54391, n54392, n54393,
         n54394, n54395, n54396, n54397, n54398, n54399, n54400, n54401,
         n54402, n54403, n54404, n54405, n54406, n54407, n54408, n54409,
         n54410, n54411, n54412, n54413, n54414, n54415, n54416, n54417,
         n54418, n54419, n54420, n54421, n54422, n54423, n54424, n54425,
         n54426, n54427, n54428, n54429, n54430, n54431, n54432, n54433,
         n54434, n54435, n54436, n54437, n54438, n54439, n54440, n54441,
         n54442, n54443, n54444, n54445, n54446, n54447, n54448, n54449,
         n54450, n54451, n54452, n54453, n54454, n54455, n54456, n54457,
         n54458, n54459, n54460, n54461, n54462, n54463, n54464, n54465,
         n54466, n54467, n54468, n54469, n54470, n54471, n54472, n54473,
         n54474, n54475, n54476, n54477, n54478, n54479, n54480, n54481,
         n54482, n54483, n54484, n54485, n54486, n54487, n54488, n54489,
         n54490, n54491, n54492, n54493, n54494, n54495, n54496, n54497,
         n54498, n54499, n54500, n54501, n54502, n54503, n54504, n54505,
         n54506, n54507, n54508, n54509, n54510, n54511, n54512, n54513,
         n54514, n54515, n54516, n54517, n54518, n54519, n54520, n54521,
         n54522, n54523, n54524, n54525, n54526, n54527, n54528, n54529,
         n54530, n54531, n54532, n54533, n54534, n54535, n54536, n54537,
         n54538, n54539, n54540, n54541, n54542, n54543, n54544, n54545,
         n54546, n54547, n54548, n54549, n54550, n54551, n54552, n54553,
         n54554, n54555, n54556, n54557, n54558, n54559, n54560, n54561,
         n54562, n54563, n54564, n54565, n54566, n54567, n54568, n54569,
         n54570, n54571, n54572, n54573, n54574, n54575, n54576, n54577,
         n54578, n54579, n54580, n54581, n54582, n54583, n54584, n54585,
         n54586, n54587, n54588, n54589, n54590, n54591, n54592, n54593,
         n54594, n54595, n54596, n54597, n54598, n54599, n54600, n54601,
         n54602, n54603, n54604, n54605, n54606, n54607, n54608, n54609,
         n54610, n54611, n54612, n54613, n54614, n54615, n54616, n54617,
         n54618, n54619, n54620, n54621, n54622, n54623, n54624, n54625,
         n54626, n54627, n54628, n54629, n54630, n54631, n54632, n54633,
         n54634, n54635, n54636, n54637, n54638, n54639, n54640, n54641,
         n54642, n54643, n54644, n54645, n54646, n54647, n54648, n54649,
         n54650, n54651, n54652, n54653, n54654, n54655, n54656, n54657,
         n54658, n54659, n54660, n54661, n54662, n54663, n54664, n54665,
         n54666, n54667, n54668, n54669, n54670, n54671, n54672, n54673,
         n54674, n54675, n54676, n54677, n54678, n54679, n54680, n54681,
         n54682, n54683, n54684, n54685, n54686, n54687, n54688, n54689,
         n54690, n54691, n54692, n54693, n54694, n54695, n54696, n54697,
         n54698, n54699, n54700, n54701, n54702, n54703, n54704, n54705,
         n54706, n54707, n54708, n54709, n54710, n54711, n54712, n54713,
         n54714, n54715, n54716, n54717, n54718, n54719, n54720, n54721,
         n54722, n54723, n54724, n54725, n54726, n54727, n54728, n54729,
         n54730, n54731, n54732, n54733, n54734, n54735, n54736, n54737,
         n54738, n54739, n54740, n54741, n54742, n54743, n54744, n54745,
         n54746, n54747, n54748, n54749, n54750, n54751, n54752, n54753,
         n54754, n54755, n54756, n54757, n54758, n54759, n54760, n54761,
         n54762, n54763, n54764, n54765, n54766, n54767, n54768, n54769,
         n54770, n54771, n54772, n54773, n54774, n54775, n54776, n54777,
         n54778, n54779, n54780, n54781, n54782, n54783, n54784, n54785,
         n54786, n54787, n54788, n54789, n54790, n54791, n54792, n54793,
         n54794, n54795, n54796, n54797, n54798, n54799, n54800, n54801,
         n54802, n54803, n54804, n54805, n54806, n54807, n54808, n54809,
         n54810, n54811, n54812, n54813, n54814, n54815, n54816, n54817,
         n54818, n54819, n54820, n54821, n54822, n54823, n54824, n54825,
         n54826, n54827, n54828, n54829, n54830, n54831, n54832, n54833,
         n54834, n54835, n54836, n54837, n54838, n54839, n54840, n54841,
         n54842, n54843, n54844, n54845, n54846, n54847, n54848, n54849,
         n54850, n54851, n54852, n54853, n54854, n54855, n54856, n54857,
         n54858, n54859, n54860, n54861, n54862, n54863, n54864, n54865,
         n54866, n54867, n54868, n54869, n54870, n54871, n54872, n54873,
         n54874, n54875, n54876, n54877, n54878, n54879, n54880, n54881,
         n54882, n54883, n54884, n54885, n54886, n54887, n54888, n54889,
         n54890, n54891, n54892, n54893, n54894, n54895, n54896, n54897,
         n54898, n54899, n54900, n54901, n54902, n54903, n54904, n54905,
         n54906, n54907, n54908, n54909, n54910, n54911, n54912, n54913,
         n54914, n54915, n54916, n54917, n54918, n54919, n54920, n54921,
         n54922, n54923, n54924, n54925, n54926, n54927, n54928, n54929,
         n54930, n54931, n54932, n54933, n54934, n54935, n54936, n54937,
         n54938, n54939, n54940, n54941, n54942, n54943, n54944, n54945,
         n54946, n54947, n54948, n54949, n54950, n54951, n54952, n54953,
         n54954, n54955, n54956, n54957, n54958, n54959, n54960, n54961,
         n54962, n54963, n54964, n54965, n54966, n54967, n54968, n54969,
         n54970, n54971, n54972, n54973, n54974, n54975, n54976, n54977,
         n54978, n54979, n54980, n54981, n54982, n54983, n54984, n54985,
         n54986, n54987, n54988, n54989, n54990, n54991, n54992, n54993,
         n54994, n54995, n54996, n54997, n54998, n54999, n55000, n55001,
         n55002, n55003, n55004, n55005, n55006, n55007, n55008, n55009,
         n55010, n55011, n55012, n55013, n55014, n55015, n55016, n55017,
         n55018, n55019, n55020, n55021, n55022, n55023, n55024, n55025,
         n55026, n55027, n55028, n55029, n55030, n55031, n55032, n55033,
         n55034, n55035, n55036, n55037, n55038, n55039, n55040, n55041,
         n55042, n55043, n55044, n55045, n55046, n55047, n55048, n55049,
         n55050, n55051, n55052, n55053, n55054, n55055, n55056, n55057,
         n55058, n55059, n55060, n55061, n55062, n55063, n55064, n55065,
         n55066, n55067, n55068, n55069, n55070, n55071, n55072, n55073,
         n55074, n55075, n55076, n55077, n55078, n55079, n55080, n55081,
         n55082, n55083, n55084, n55085, n55086, n55087, n55088, n55089,
         n55090, n55091, n55092, n55093, n55094, n55095, n55096, n55097,
         n55098, n55099, n55100, n55101, n55102, n55103, n55104, n55105,
         n55106, n55107, n55108, n55109, n55110, n55111, n55112, n55113,
         n55114, n55115, n55116, n55117, n55118, n55119, n55120, n55121,
         n55122, n55123, n55124, n55125, n55126, n55127, n55128, n55129,
         n55130, n55131, n55132, n55133, n55134, n55135, n55136, n55137,
         n55138, n55139, n55140, n55141, n55142, n55143, n55144, n55145,
         n55146, n55147, n55148, n55149, n55150, n55151, n55152, n55153,
         n55154, n55155, n55156, n55157, n55158, n55159, n55160, n55161,
         n55162, n55163, n55164, n55165, n55166, n55167, n55168, n55169,
         n55170, n55171, n55172, n55173, n55174, n55175, n55176, n55177,
         n55178, n55179, n55180, n55181, n55182, n55183, n55184, n55185,
         n55186, n55187, n55188, n55189, n55190, n55191, n55192, n55193,
         n55194, n55195, n55196, n55197, n55198, n55199, n55200, n55201,
         n55202, n55203, n55204, n55205, n55206, n55207, n55208, n55209,
         n55210, n55211, n55212, n55213, n55214, n55215, n55216, n55217,
         n55218, n55219, n55220, n55221, n55222, n55223, n55224, n55225,
         n55226, n55227, n55228, n55229, n55230, n55231, n55232, n55233,
         n55234, n55235, n55236, n55237, n55238, n55239, n55240, n55241,
         n55242, n55243, n55244, n55245, n55246, n55247, n55248, n55249,
         n55250, n55251, n55252, n55253, n55254, n55255, n55256, n55257,
         n55258, n55259, n55260, n55261, n55262, n55263, n55264, n55265,
         n55266, n55267, n55268, n55269, n55270, n55271, n55272, n55273,
         n55274, n55275, n55276, n55277, n55278, n55279, n55280, n55281,
         n55282, n55283, n55284, n55285, n55286, n55287, n55288, n55289,
         n55290, n55291, n55292, n55293, n55294, n55295, n55296, n55297,
         n55298, n55299, n55300, n55301, n55302, n55303, n55304, n55305,
         n55306, n55307, n55308, n55309, n55310, n55311, n55312, n55313,
         n55314, n55315, n55316, n55317, n55318, n55319, n55320, n55321,
         n55322, n55323, n55324, n55325, n55326, n55327, n55328, n55329,
         n55330, n55331, n55332, n55333, n55334, n55335, n55336, n55337,
         n55338, n55339, n55340, n55341, n55342, n55343, n55344, n55345,
         n55346, n55347, n55348, n55349, n55350, n55351, n55352, n55353,
         n55354, n55355, n55356, n55357, n55358, n55359, n55360, n55361,
         n55362;
  wire   [31:6] w_PC_OUT;
  wire   [31:0] w_IR_OUT;
  wire   [4:0] w_ALU_OPCODE;
  wire   [2:0] w_MuxLD_SEL;
  wire   [2:0] w_MuxSW_SEL;
  wire   [4:0] w_RS2;
  assign IRAM_ADDR[1] = \DP/NPC[1] ;
  assign IRAM_ADDR[0] = \DP/NPC[0] ;

  DFF_X1 \PC/DOUT_reg[4]  ( .D(n5089), .CK(n5185), .Q(IRAM_ADDR[4]), .QN(n3270) );
  DFF_X1 \PC/DOUT_reg[16]  ( .D(n5090), .CK(n5185), .QN(n53690) );
  DFF_X1 \PC/DOUT_reg[21]  ( .D(n5091), .CK(n5185), .Q(w_PC_OUT[21]) );
  DFF_X1 \PC/DOUT_reg[14]  ( .D(n5092), .CK(n5185), .Q(n53594), .QN(n53675) );
  DFF_X1 \PC/DOUT_reg[22]  ( .D(n5093), .CK(n5185), .QN(n53655) );
  DFF_X1 \PC/DOUT_reg[10]  ( .D(n5094), .CK(n5185), .QN(n53656) );
  DFF_X1 \PC/DOUT_reg[26]  ( .D(n5095), .CK(n5185), .QN(n53674) );
  DFF_X1 \PC/DOUT_reg[5]  ( .D(n5097), .CK(n5185), .Q(IRAM_ADDR[5]), .QN(n7230) );
  DFF_X1 \PC/DOUT_reg[19]  ( .D(n5098), .CK(n5185), .Q(w_PC_OUT[19]) );
  DFF_X1 \PC/DOUT_reg[28]  ( .D(n5099), .CK(n5185), .Q(n53601), .QN(n53676) );
  DFF_X1 \PC/DOUT_reg[30]  ( .D(n5100), .CK(n5185), .QN(n49845) );
  DFF_X1 \PC/DOUT_reg[1]  ( .D(n5101), .CK(n5185), .Q(\DP/NPC[1] ), .QN(n7227)
         );
  DFF_X1 \PC/DOUT_reg[2]  ( .D(n5102), .CK(n5185), .Q(IRAM_ADDR[2]), .QN(n7228) );
  DFF_X1 \PC/DOUT_reg[17]  ( .D(n5103), .CK(n5185), .Q(w_PC_OUT[17]) );
  DFF_X1 \PC/DOUT_reg[12]  ( .D(n5104), .CK(n5185), .QN(n53659) );
  DFF_X1 \PC/DOUT_reg[15]  ( .D(n5105), .CK(n5185), .Q(w_PC_OUT[15]) );
  DFF_X1 \PC/DOUT_reg[13]  ( .D(n5106), .CK(n5185), .Q(w_PC_OUT[13]) );
  DFF_X1 \PC/DOUT_reg[23]  ( .D(n5107), .CK(n5185), .Q(w_PC_OUT[23]), .QN(
        n53792) );
  DFF_X1 \PC/DOUT_reg[24]  ( .D(n5108), .CK(n5185), .QN(n53700) );
  DFF_X1 \PC/DOUT_reg[29]  ( .D(n5109), .CK(n5185), .Q(w_PC_OUT[29]), .QN(
        n53776) );
  DFF_X1 \PC/DOUT_reg[27]  ( .D(n5110), .CK(n5185), .Q(w_PC_OUT[27]) );
  DFF_X1 \PC/DOUT_reg[20]  ( .D(n5111), .CK(n5185), .QN(n53658) );
  DFF_X1 \PC/DOUT_reg[18]  ( .D(n5112), .CK(n5185), .QN(n53691) );
  DFF_X1 \PC/DOUT_reg[0]  ( .D(n5113), .CK(n5185), .Q(\DP/NPC[0] ), .QN(n7226)
         );
  DFF_X1 \PC/DOUT_reg[11]  ( .D(n5114), .CK(n5185), .Q(w_PC_OUT[11]), .QN(
        n53785) );
  DFF_X1 \PC/DOUT_reg[8]  ( .D(n5115), .CK(n5185), .QN(n53657) );
  DFF_X1 \PC/DOUT_reg[25]  ( .D(n5116), .CK(n5185), .Q(w_PC_OUT[25]), .QN(
        n53744) );
  DFF_X1 \PC/DOUT_reg[31]  ( .D(n5117), .CK(n5185), .Q(w_PC_OUT[31]) );
  DFF_X1 \PC/DOUT_reg[3]  ( .D(n5118), .CK(n5185), .Q(IRAM_ADDR[3]), .QN(n7229) );
  DFF_X1 \PC/DOUT_reg[7]  ( .D(n5120), .CK(n5185), .Q(w_PC_OUT[7]) );
  DFF_X1 \IR/DOUT_reg[31]  ( .D(n5123), .CK(n5185), .Q(w_IR_OUT[31]), .QN(
        n53653) );
  DFFR_X1 \CU/cw2_reg[18]  ( .D(\CU/cw1[18] ), .CK(CLK), .RN(RST), .Q(
        w_MuxIMM_SEL) );
  DFFR_X1 \CU/cw3_reg[15]  ( .D(\CU/cw2[15] ), .CK(CLK), .RN(RST), .Q(
        w_MuxA_SEL), .QN(n53763) );
  DFFR_X1 \CU/cw3_reg[14]  ( .D(\CU/cw2[14] ), .CK(CLK), .RN(RST), .Q(
        w_MuxB_SEL), .QN(n53762) );
  DFFR_X1 \CU/aluOpcode3_reg[0]  ( .D(\CU/aluOpcode2[0] ), .CK(CLK), .RN(RST), 
        .Q(w_ALU_OPCODE[0]), .QN(n53646) );
  DFFR_X1 \CU/aluOpcode2_reg[0]  ( .D(\CU/aluOpcode1[0] ), .CK(CLK), .RN(RST), 
        .Q(\CU/aluOpcode2[0] ) );
  DFFR_X1 \CU/aluOpcode3_reg[1]  ( .D(\CU/aluOpcode2[1] ), .CK(CLK), .RN(RST), 
        .Q(w_ALU_OPCODE[1]), .QN(n53679) );
  DFFR_X1 \CU/aluOpcode2_reg[1]  ( .D(\CU/aluOpcode1[1] ), .CK(CLK), .RN(RST), 
        .Q(\CU/aluOpcode2[1] ) );
  DFFR_X1 \CU/aluOpcode3_reg[2]  ( .D(\CU/aluOpcode2[2] ), .CK(CLK), .RN(RST), 
        .Q(w_ALU_OPCODE[2]), .QN(n53680) );
  DFFR_X1 \CU/aluOpcode2_reg[2]  ( .D(\CU/aluOpcode1[2] ), .CK(CLK), .RN(RST), 
        .Q(\CU/aluOpcode2[2] ) );
  DFFR_X1 \CU/aluOpcode3_reg[3]  ( .D(\CU/aluOpcode2[3] ), .CK(CLK), .RN(RST), 
        .Q(w_ALU_OPCODE[3]) );
  DFFR_X1 \CU/aluOpcode2_reg[3]  ( .D(\CU/aluOpcode1[3] ), .CK(CLK), .RN(RST), 
        .Q(\CU/aluOpcode2[3] ) );
  DFFR_X1 \CU/aluOpcode3_reg[4]  ( .D(\CU/aluOpcode2[4] ), .CK(CLK), .RN(RST), 
        .Q(w_ALU_OPCODE[4]), .QN(n53692) );
  DFFR_X1 \CU/aluOpcode2_reg[4]  ( .D(\CU/aluOpcode1[4] ), .CK(CLK), .RN(RST), 
        .Q(\CU/aluOpcode2[4] ) );
  DFFR_X1 \CU/aluOpcode1_reg[0]  ( .D(\CU/aluOpcodei[0] ), .CK(CLK), .RN(RST), 
        .Q(\CU/aluOpcode1[0] ) );
  DFFR_X1 \CU/aluOpcode1_reg[1]  ( .D(\CU/aluOpcodei[1] ), .CK(CLK), .RN(RST), 
        .Q(\CU/aluOpcode1[1] ) );
  DFFR_X1 \CU/aluOpcode1_reg[2]  ( .D(\CU/aluOpcodei[2] ), .CK(CLK), .RN(RST), 
        .Q(\CU/aluOpcode1[2] ) );
  DFFR_X1 \CU/aluOpcode1_reg[3]  ( .D(\CU/aluOpcodei[3] ), .CK(CLK), .RN(RST), 
        .Q(\CU/aluOpcode1[3] ) );
  DFFR_X1 \CU/aluOpcode1_reg[4]  ( .D(\CU/aluOpcodei[4] ), .CK(CLK), .RN(RST), 
        .Q(\CU/aluOpcode1[4] ) );
  DFFR_X1 \CU/cw5_reg[1]  ( .D(\CU/cw4[1] ), .CK(CLK), .RN(RST), .Q(w_RF_WE)
         );
  DFFR_X1 \CU/cw4_reg[0]  ( .D(\CU/cw3[0] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw4[0] ) );
  DFFR_X1 \CU/cw4_reg[1]  ( .D(\CU/cw3[1] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw4[1] ) );
  DFFR_X1 \CU/cw4_reg[2]  ( .D(\CU/cw3[2] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw4[2] ) );
  DFFR_X1 \CU/cw4_reg[3]  ( .D(\CU/cw3[3] ), .CK(CLK), .RN(RST), .Q(
        w_MuxSW_SEL[0]) );
  DFFR_X1 \CU/cw4_reg[4]  ( .D(\CU/cw3[4] ), .CK(CLK), .RN(RST), .Q(
        w_MuxSW_SEL[1]), .QN(n53752) );
  DFFR_X1 \CU/cw4_reg[5]  ( .D(\CU/cw3[5] ), .CK(CLK), .RN(RST), .Q(
        w_MuxSW_SEL[2]), .QN(n53677) );
  DFFR_X1 \CU/cw4_reg[6]  ( .D(\CU/cw3[6] ), .CK(CLK), .RN(RST), .Q(
        w_MuxLD_SEL[0]) );
  DFFR_X1 \CU/cw4_reg[7]  ( .D(\CU/cw3[7] ), .CK(CLK), .RN(RST), .Q(
        w_MuxLD_SEL[1]), .QN(n53701) );
  DFFR_X1 \CU/cw4_reg[8]  ( .D(w_RF_WE3), .CK(CLK), .RN(RST), .Q(w_RF_WE4), 
        .QN(n53654) );
  DFFR_X1 \CU/cw4_reg[9]  ( .D(\CU/cw3_9 ), .CK(CLK), .RN(RST), .Q(
        w_SIGN_LD_EN) );
  DFFR_X1 \CU/cw4_reg[10]  ( .D(\CU/cw3_10 ), .CK(CLK), .RN(RST), .Q(DRAM_RW)
         );
  DFFR_X1 \CU/cw4_reg[11]  ( .D(\CU/cw3_11 ), .CK(CLK), .RN(RST), .Q(DRAM_EN), 
        .QN(n3021) );
  DFFR_X1 \CU/cw3_reg[0]  ( .D(\CU/cw2[0] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw3[0] ) );
  DFFR_X1 \CU/cw3_reg[1]  ( .D(\CU/cw2[1] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw3[1] ) );
  DFFR_X1 \CU/cw3_reg[2]  ( .D(\CU/cw2[2] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw3[2] ) );
  DFFR_X1 \CU/cw3_reg[3]  ( .D(\CU/cw2[3] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw3[3] ) );
  DFFR_X1 \CU/cw3_reg[4]  ( .D(\CU/cw2[4] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw3[4] ) );
  DFFR_X1 \CU/cw3_reg[5]  ( .D(\CU/cw2[5] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw3[5] ) );
  DFFR_X1 \CU/cw3_reg[6]  ( .D(\CU/cw2[6] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw3[6] ) );
  DFFR_X1 \CU/cw3_reg[7]  ( .D(\CU/cw2[7] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw3[7] ) );
  DFFR_X1 \CU/cw3_reg[8]  ( .D(\CU/cw2[8] ), .CK(CLK), .RN(RST), .Q(w_RF_WE3)
         );
  DFFR_X1 \CU/cw3_reg[9]  ( .D(\CU/cw2[9] ), .CK(CLK), .RN(RST), .Q(\CU/cw3_9 ) );
  DFFR_X1 \CU/cw3_reg[10]  ( .D(\CU/cw2[10] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw3_10 ) );
  DFFR_X1 \CU/cw3_reg[11]  ( .D(\CU/cw2[11] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw3_11 ), .QN(n3020) );
  DFFR_X1 \CU/cw3_reg[12]  ( .D(\CU/cw2[12] ), .CK(CLK), .RN(RST), .Q(
        w_JUMP_EN) );
  DFFR_X1 \CU/cw3_reg[13]  ( .D(\CU/cw2[13] ), .CK(CLK), .RN(RST), .Q(
        w_EQ_COND) );
  DFFR_X1 \CU/cw2_reg[0]  ( .D(\CU/cw1[0] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[0] ) );
  DFFR_X1 \CU/cw2_reg[1]  ( .D(\CU/cw1[1] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[1] ) );
  DFFR_X1 \CU/cw2_reg[2]  ( .D(\CU/cw1[2] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[2] ) );
  DFFR_X1 \CU/cw2_reg[3]  ( .D(\CU/cw1[3] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[3] ) );
  DFFR_X1 \CU/cw2_reg[4]  ( .D(\CU/cw1[4] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[4] ) );
  DFFR_X1 \CU/cw2_reg[5]  ( .D(\CU/cw1[5] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[5] ) );
  DFFR_X1 \CU/cw2_reg[6]  ( .D(\CU/cw1[6] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[6] ) );
  DFFR_X1 \CU/cw2_reg[7]  ( .D(\CU/cw1[7] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[7] ) );
  DFFR_X1 \CU/cw2_reg[8]  ( .D(\CU/cw1[8] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[8] ) );
  DFFR_X1 \CU/cw2_reg[9]  ( .D(\CU/cw1[9] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[9] ) );
  DFFR_X1 \CU/cw2_reg[10]  ( .D(\CU/cw1[10] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[10] ) );
  DFFR_X1 \CU/cw2_reg[11]  ( .D(\CU/cw1[11] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[11] ), .QN(n3019) );
  DFFR_X1 \CU/cw2_reg[12]  ( .D(\CU/cw1[12] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[12] ) );
  DFFR_X1 \CU/cw2_reg[13]  ( .D(\CU/cw1[13] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[13] ) );
  DFFR_X1 \CU/cw2_reg[14]  ( .D(\CU/cw1[14] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[14] ) );
  DFFR_X1 \CU/cw2_reg[15]  ( .D(\CU/cw1[15] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw2[15] ) );
  DFFR_X1 \CU/cw2_reg[17]  ( .D(\CU/cw1[17] ), .CK(CLK), .RN(RST), .Q(
        w_SIGN_EN) );
  DFFR_X1 \CU/cw2_reg[19]  ( .D(\CU/cw1[19] ), .CK(CLK), .RN(RST), .Q(w_RF_RD2) );
  DFFR_X1 \CU/cw2_reg[20]  ( .D(\CU/cw1[20] ), .CK(CLK), .RN(RST), .Q(w_RF_RD1) );
  DFFR_X1 \CU/cw1_reg[0]  ( .D(n45959), .CK(CLK), .RN(RST), .Q(\CU/cw1[0] ) );
  DFFR_X1 \CU/cw1_reg[1]  ( .D(\CU/n142 ), .CK(CLK), .RN(RST), .Q(\CU/cw1[1] )
         );
  DFFR_X1 \CU/cw1_reg[2]  ( .D(n49781), .CK(CLK), .RN(RST), .Q(\CU/cw1[2] ) );
  DFFR_X1 \CU/cw1_reg[3]  ( .D(\CU/cw[3] ), .CK(CLK), .RN(RST), .Q(\CU/cw1[3] ) );
  DFFR_X1 \CU/cw1_reg[4]  ( .D(\CU/n140 ), .CK(CLK), .RN(RST), .Q(\CU/cw1[4] )
         );
  DFFR_X1 \CU/cw1_reg[5]  ( .D(\CU/n139 ), .CK(CLK), .RN(RST), .Q(\CU/cw1[5] )
         );
  DFFR_X1 \CU/cw1_reg[6]  ( .D(\CU/cw[6] ), .CK(CLK), .RN(RST), .Q(\CU/cw1[6] ) );
  DFFR_X1 \CU/cw1_reg[7]  ( .D(n3024), .CK(CLK), .RN(RST), .Q(\CU/cw1[7] ) );
  DFFR_X1 \CU/cw1_reg[8]  ( .D(n3022), .CK(CLK), .RN(RST), .Q(\CU/cw1[8] ) );
  DFFR_X1 \CU/cw1_reg[10]  ( .D(n32415), .CK(CLK), .RN(RST), .Q(\CU/cw1[10] )
         );
  DFFR_X1 \CU/cw1_reg[11]  ( .D(\CU/cw[21] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw1[11] ) );
  DFFR_X1 \CU/cw1_reg[12]  ( .D(n32429), .CK(CLK), .RN(RST), .Q(\CU/cw1[12] )
         );
  DFFR_X1 \CU/cw1_reg[13]  ( .D(\CU/n138 ), .CK(CLK), .RN(RST), .Q(
        \CU/cw1[13] ) );
  DFFR_X1 \CU/cw1_reg[14]  ( .D(n3025), .CK(CLK), .RN(RST), .Q(\CU/cw1[14] )
         );
  DFFR_X1 \CU/cw1_reg[17]  ( .D(\CU/cw[17] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw1[17] ) );
  DFFR_X1 \CU/cw1_reg[18]  ( .D(\CU/cw[18] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw1[18] ) );
  DFFR_X1 \CU/cw1_reg[20]  ( .D(\CU/cw[20] ), .CK(CLK), .RN(RST), .Q(
        \CU/cw1[20] ) );
  DFFR_X1 \CU/cw1_reg[22]  ( .D(1'b1), .CK(CLK), .RN(RST), .Q(IRAM_EN), .QN(
        n3018) );
  REGISTER_FILE_WIDTH32_LENGTH5 \DP/RegFILE  ( .CLK(CLK), .RST(RST), .EN(
        \CU/cw2[11] ), .RD1(w_RF_RD1), .RD2(w_RF_RD2), .WR(w_RF_WE), .DATAIN({
        n3056, n3054, n3039, n3057, n3041, n3055, n3040, n3038, n3044, n3045, 
        n3046, n3042, n3047, n3048, n3043, n3049, n3051, n3053, n3052, n3050, 
        n3032, n3028, n3029, n3033, n3034, n51623, n3036, n43969, n43968, 
        n51619, n3026, n3027}), .OUT1({\DP/RegA_IN[31] , \DP/RegA_IN[30] , 
        \DP/RegA_IN[29] , \DP/RegA_IN[28] , \DP/RegA_IN[27] , \DP/RegA_IN[26] , 
        \DP/RegA_IN[25] , \DP/RegA_IN[24] , \DP/RegA_IN[23] , \DP/RegA_IN[22] , 
        \DP/RegA_IN[21] , \DP/RegA_IN[20] , \DP/RegA_IN[19] , \DP/RegA_IN[18] , 
        \DP/RegA_IN[17] , \DP/RegA_IN[16] , \DP/RegA_IN[15] , \DP/RegA_IN[14] , 
        \DP/RegA_IN[13] , \DP/RegA_IN[12] , \DP/RegA_IN[11] , \DP/RegA_IN[10] , 
        \DP/RegA_IN[9] , \DP/RegA_IN[8] , \DP/RegA_IN[7] , \DP/RegA_IN[6] , 
        \DP/RegA_IN[5] , \DP/RegA_IN[4] , \DP/RegA_IN[3] , \DP/RegA_IN[2] , 
        \DP/RegA_IN[1] , \DP/RegA_IN[0] }), .OUT2({\DP/RegB_IN[31] , 
        \DP/RegB_IN[30] , \DP/RegB_IN[29] , \DP/RegB_IN[28] , \DP/RegB_IN[27] , 
        \DP/RegB_IN[26] , \DP/RegB_IN[25] , \DP/RegB_IN[24] , \DP/RegB_IN[23] , 
        \DP/RegB_IN[22] , \DP/RegB_IN[21] , \DP/RegB_IN[20] , \DP/RegB_IN[19] , 
        \DP/RegB_IN[18] , \DP/RegB_IN[17] , \DP/RegB_IN[16] , \DP/RegB_IN[15] , 
        \DP/RegB_IN[14] , \DP/RegB_IN[13] , \DP/RegB_IN[12] , \DP/RegB_IN[11] , 
        \DP/RegB_IN[10] , \DP/RegB_IN[9] , \DP/RegB_IN[8] , \DP/RegB_IN[7] , 
        \DP/RegB_IN[6] , \DP/RegB_IN[5] , \DP/RegB_IN[4] , \DP/RegB_IN[3] , 
        \DP/RegB_IN[2] , \DP/RegB_IN[1] , \DP/RegB_IN[0] }), .ADD_WR({
        \DP/RD4[4] , \DP/RD4[3] , \DP/RD4[2] , \DP/RD4[1] , \DP/RD4[0] }), 
        .ADD_RD1({\DP/IMMS26[25] , \DP/IMMS26[24] , \DP/IMMS26[23] , 
        \DP/IMMS26[22] , \DP/IMMS26[21] }), .ADD_RD2(w_RS2) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[0]  ( .D(n5154), .CK(n5185), .Q(n53562) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[1]  ( .D(n5155), .CK(n5185), .Q(n53563) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[2]  ( .D(n5156), .CK(n5185), .Q(n53564) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[3]  ( .D(n7489), .CK(n5185), .Q(n53565) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[4]  ( .D(n5158), .CK(n5185), .Q(n53566) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[5]  ( .D(n7478), .CK(n5185), .Q(n53567) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[6]  ( .D(n47727), .CK(n5185), .Q(n53568) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[7]  ( .D(n51537), .CK(n5185), .Q(n53569) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[8]  ( .D(n47726), .CK(n5185), .Q(n53570) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[9]  ( .D(n51536), .CK(n5185), .Q(n53571) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[10]  ( .D(n43886), .CK(n5185), .Q(n53572) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[11]  ( .D(n51535), .CK(n5185), .Q(n53573) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[12]  ( .D(n40065), .CK(n5185), .Q(n53574) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[13]  ( .D(n53610), .CK(n5185), .Q(n53575) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[14]  ( .D(n51533), .CK(n5185), .Q(n53576) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[15]  ( .D(n53609), .CK(n5185), .Q(n53577) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[16]  ( .D(n51532), .CK(n5185), .Q(n53578) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[17]  ( .D(n53608), .CK(n5185), .Q(n53579) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[18]  ( .D(n51531), .CK(n5185), .Q(n53580) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[19]  ( .D(n53607), .CK(n5185), .Q(n53581) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[20]  ( .D(n40060), .CK(n5185), .Q(n53582) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[21]  ( .D(n51529), .CK(n5185), .Q(n53583) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[22]  ( .D(n40059), .CK(n5185), .Q(n53584) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[23]  ( .D(n53606), .CK(n5185), .Q(n53585) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[24]  ( .D(n51527), .CK(n5185), .Q(n53586) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[25]  ( .D(n53605), .CK(n5185), .Q(n53587) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[26]  ( .D(n51524), .CK(n5185), .Q(n53588) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[27]  ( .D(n53604), .CK(n5185), .Q(n53589) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[28]  ( .D(n51525), .CK(n5185), .Q(n53590) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[29]  ( .D(n53603), .CK(n5185), .Q(n53591) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[30]  ( .D(n5184), .CK(n5185), .Q(n53592) );
  DFF_X1 \DP/RegA/DOUT_reg[0]  ( .D(n5186), .CK(n5307), .QN(n53499) );
  DFF_X1 \DP/RegA/DOUT_reg[1]  ( .D(n5187), .CK(n5307), .QN(n53506) );
  DFF_X1 \DP/RegA/DOUT_reg[2]  ( .D(n5188), .CK(n5307), .QN(n53505) );
  DFF_X1 \DP/RegA/DOUT_reg[3]  ( .D(n5189), .CK(n5307), .QN(n53504) );
  DFF_X1 \DP/RegA/DOUT_reg[4]  ( .D(n5190), .CK(n5307), .QN(n53503) );
  DFF_X1 \DP/RegA/DOUT_reg[5]  ( .D(n5191), .CK(n5307), .QN(n53510) );
  DFF_X1 \DP/RegA/DOUT_reg[6]  ( .D(n5192), .CK(n5307), .QN(n53509) );
  DFF_X1 \DP/RegA/DOUT_reg[7]  ( .D(n5193), .CK(n5307), .QN(n53508) );
  DFF_X1 \DP/RegA/DOUT_reg[8]  ( .D(n5194), .CK(n5307), .QN(n53507) );
  DFF_X1 \DP/RegA/DOUT_reg[9]  ( .D(n5195), .CK(n5307), .QN(n53514) );
  DFF_X1 \DP/RegA/DOUT_reg[10]  ( .D(n5196), .CK(n5307), .QN(n53512) );
  DFF_X1 \DP/RegA/DOUT_reg[11]  ( .D(n5197), .CK(n5307), .QN(n53511) );
  DFF_X1 \DP/RegA/DOUT_reg[12]  ( .D(n5198), .CK(n5307), .QN(n53483) );
  DFF_X1 \DP/RegA/DOUT_reg[13]  ( .D(n5199), .CK(n5307), .QN(n53490) );
  DFF_X1 \DP/RegA/DOUT_reg[14]  ( .D(n5200), .CK(n5307), .QN(n53489) );
  DFF_X1 \DP/RegA/DOUT_reg[15]  ( .D(n5201), .CK(n5307), .QN(n53488) );
  DFF_X1 \DP/RegA/DOUT_reg[16]  ( .D(n5202), .CK(n5307), .QN(n53487) );
  DFF_X1 \DP/RegA/DOUT_reg[17]  ( .D(n5203), .CK(n5307), .QN(n53494) );
  DFF_X1 \DP/RegA/DOUT_reg[18]  ( .D(n5204), .CK(n5307), .QN(n53493) );
  DFF_X1 \DP/RegA/DOUT_reg[19]  ( .D(n5205), .CK(n5307), .QN(n53492) );
  DFF_X1 \DP/RegA/DOUT_reg[20]  ( .D(n5206), .CK(n5307), .QN(n53491) );
  DFF_X1 \DP/RegA/DOUT_reg[21]  ( .D(n5207), .CK(n5307), .QN(n53498) );
  DFF_X1 \DP/RegA/DOUT_reg[22]  ( .D(n5208), .CK(n5307), .QN(n53497) );
  DFF_X1 \DP/RegA/DOUT_reg[23]  ( .D(n5209), .CK(n5307), .QN(n53496) );
  DFF_X1 \DP/RegA/DOUT_reg[24]  ( .D(n5210), .CK(n5307), .QN(n53495) );
  DFF_X1 \DP/RegA/DOUT_reg[25]  ( .D(n5211), .CK(n5307), .QN(n53485) );
  DFF_X1 \DP/RegA/DOUT_reg[26]  ( .D(n5212), .CK(n5307), .QN(n53502) );
  DFF_X1 \DP/RegA/DOUT_reg[27]  ( .D(n5213), .CK(n5307), .QN(n53501) );
  DFF_X1 \DP/RegA/DOUT_reg[28]  ( .D(n5214), .CK(n5307), .QN(n53500) );
  DFF_X1 \DP/RegA/DOUT_reg[29]  ( .D(n5215), .CK(n5307), .QN(n53484) );
  DFF_X1 \DP/RegA/DOUT_reg[30]  ( .D(n5216), .CK(n5307), .QN(n53486) );
  DFF_X1 \DP/RegA/DOUT_reg[31]  ( .D(n5217), .CK(n5307), .QN(n53513) );
  DFF_X1 \DP/RegB/DOUT_reg[0]  ( .D(n5218), .CK(n5307), .QN(n53419) );
  DFF_X1 \DP/RegB/DOUT_reg[1]  ( .D(n5219), .CK(n5307), .QN(n53420) );
  DFF_X1 \DP/RegB/DOUT_reg[2]  ( .D(n5220), .CK(n5307), .QN(n53421) );
  DFF_X1 \DP/RegB/DOUT_reg[3]  ( .D(n5221), .CK(n5307), .QN(n53422) );
  DFF_X1 \DP/RegB/DOUT_reg[4]  ( .D(n5222), .CK(n5307), .QN(n53423) );
  DFF_X1 \DP/RegB/DOUT_reg[5]  ( .D(n5223), .CK(n5307), .QN(n53424) );
  DFF_X1 \DP/RegB/DOUT_reg[6]  ( .D(n5224), .CK(n5307), .QN(n53425) );
  DFF_X1 \DP/RegB/DOUT_reg[7]  ( .D(n5225), .CK(n5307), .QN(n53426) );
  DFF_X1 \DP/RegB/DOUT_reg[8]  ( .D(n5226), .CK(n5307), .QN(n53427) );
  DFF_X1 \DP/RegB/DOUT_reg[9]  ( .D(n5227), .CK(n5307), .QN(n53428) );
  DFF_X1 \DP/RegB/DOUT_reg[10]  ( .D(n5228), .CK(n5307), .QN(n53429) );
  DFF_X1 \DP/RegB/DOUT_reg[11]  ( .D(n5229), .CK(n5307), .QN(n53430) );
  DFF_X1 \DP/RegB/DOUT_reg[12]  ( .D(n5230), .CK(n5307), .QN(n53431) );
  DFF_X1 \DP/RegB/DOUT_reg[13]  ( .D(n5231), .CK(n5307), .QN(n53432) );
  DFF_X1 \DP/RegB/DOUT_reg[14]  ( .D(n5232), .CK(n5307), .QN(n53433) );
  DFF_X1 \DP/RegB/DOUT_reg[15]  ( .D(n5233), .CK(n5307), .QN(n53434) );
  DFF_X1 \DP/RegB/DOUT_reg[16]  ( .D(n5234), .CK(n5307), .QN(n53435) );
  DFF_X1 \DP/RegB/DOUT_reg[17]  ( .D(n5235), .CK(n5307), .QN(n53436) );
  DFF_X1 \DP/RegB/DOUT_reg[18]  ( .D(n5236), .CK(n5307), .QN(n53437) );
  DFF_X1 \DP/RegB/DOUT_reg[19]  ( .D(n5237), .CK(n5307), .QN(n53438) );
  DFF_X1 \DP/RegB/DOUT_reg[20]  ( .D(n5238), .CK(n5307), .QN(n53439) );
  DFF_X1 \DP/RegB/DOUT_reg[21]  ( .D(n5239), .CK(n5307), .QN(n53440) );
  DFF_X1 \DP/RegB/DOUT_reg[22]  ( .D(n5240), .CK(n5307), .QN(n53441) );
  DFF_X1 \DP/RegB/DOUT_reg[23]  ( .D(n5241), .CK(n5307), .QN(n53442) );
  DFF_X1 \DP/RegB/DOUT_reg[24]  ( .D(n5242), .CK(n5307), .QN(n53443) );
  DFF_X1 \DP/RegB/DOUT_reg[25]  ( .D(n5243), .CK(n5307), .QN(n53444) );
  DFF_X1 \DP/RegB/DOUT_reg[26]  ( .D(n5244), .CK(n5307), .QN(n53445) );
  DFF_X1 \DP/RegB/DOUT_reg[27]  ( .D(n5245), .CK(n5307), .QN(n53446) );
  DFF_X1 \DP/RegB/DOUT_reg[28]  ( .D(n5246), .CK(n5307), .QN(n53447) );
  DFF_X1 \DP/RegB/DOUT_reg[29]  ( .D(n5247), .CK(n5307), .QN(n53448) );
  DFF_X1 \DP/RegB/DOUT_reg[30]  ( .D(n5248), .CK(n5307), .QN(n53449) );
  DFF_X1 \DP/RegB/DOUT_reg[31]  ( .D(n5249), .CK(n5307), .QN(n53450) );
  DFF_X1 \DP/RegIMM/DOUT_reg[0]  ( .D(n5250), .CK(n5307), .QN(n53400) );
  DFF_X1 \DP/RegIMM/DOUT_reg[1]  ( .D(n5251), .CK(n5307), .QN(n53399) );
  DFF_X1 \DP/RegIMM/DOUT_reg[2]  ( .D(n5252), .CK(n5307), .QN(n53398) );
  DFF_X1 \DP/RegIMM/DOUT_reg[3]  ( .D(n5253), .CK(n5307), .QN(n53397) );
  DFF_X1 \DP/RegIMM/DOUT_reg[4]  ( .D(n5254), .CK(n5307), .QN(n53396) );
  DFF_X1 \DP/RegIMM/DOUT_reg[5]  ( .D(n5255), .CK(n5307), .QN(n53395) );
  DFF_X1 \DP/RegIMM/DOUT_reg[6]  ( .D(n5256), .CK(n5307), .QN(n53394) );
  DFF_X1 \DP/RegIMM/DOUT_reg[7]  ( .D(n5257), .CK(n5307), .QN(n53393) );
  DFF_X1 \DP/RegIMM/DOUT_reg[8]  ( .D(n5258), .CK(n5307), .QN(n53392) );
  DFF_X1 \DP/RegIMM/DOUT_reg[9]  ( .D(n5259), .CK(n5307), .QN(n53391) );
  DFF_X1 \DP/RegIMM/DOUT_reg[10]  ( .D(n5260), .CK(n5307), .QN(n53390) );
  DFF_X1 \DP/RegIMM/DOUT_reg[11]  ( .D(n5261), .CK(n5307), .QN(n53389) );
  DFF_X1 \DP/RegIMM/DOUT_reg[12]  ( .D(n5262), .CK(n5307), .QN(n53413) );
  DFF_X1 \DP/RegIMM/DOUT_reg[13]  ( .D(n5263), .CK(n5307), .QN(n53412) );
  DFF_X1 \DP/RegIMM/DOUT_reg[14]  ( .D(n5264), .CK(n5307), .QN(n53411) );
  DFF_X1 \DP/RegIMM/DOUT_reg[15]  ( .D(n5265), .CK(n5307), .QN(n53410) );
  DFF_X1 \DP/RegIMM/DOUT_reg[16]  ( .D(n5266), .CK(n5307), .QN(n53409) );
  DFF_X1 \DP/RegIMM/DOUT_reg[17]  ( .D(n5267), .CK(n5307), .QN(n53408) );
  DFF_X1 \DP/RegIMM/DOUT_reg[18]  ( .D(n5268), .CK(n5307), .QN(n53407) );
  DFF_X1 \DP/RegIMM/DOUT_reg[19]  ( .D(n5269), .CK(n5307), .QN(n53406) );
  DFF_X1 \DP/RegIMM/DOUT_reg[20]  ( .D(n5270), .CK(n5307), .QN(n53405) );
  DFF_X1 \DP/RegIMM/DOUT_reg[21]  ( .D(n5271), .CK(n5307), .QN(n53404) );
  DFF_X1 \DP/RegIMM/DOUT_reg[22]  ( .D(n5272), .CK(n5307), .QN(n53403) );
  DFF_X1 \DP/RegIMM/DOUT_reg[23]  ( .D(n5273), .CK(n5307), .QN(n53402) );
  DFF_X1 \DP/RegIMM/DOUT_reg[24]  ( .D(n5274), .CK(n5307), .QN(n53401) );
  DFF_X1 \DP/RegIMM/DOUT_reg[25]  ( .D(n1176), .CK(n5307), .QN(n53262) );
  DFF_X1 \DP/RegRD2/DOUT_reg[0]  ( .D(\DP/RegRD2/n14 ), .CK(n5307), .Q(n53270)
         );
  DFF_X1 \DP/RegRD2/DOUT_reg[1]  ( .D(\DP/RegRD2/n13 ), .CK(n5307), .Q(n53269)
         );
  DFF_X1 \DP/RegRD2/DOUT_reg[2]  ( .D(\DP/RegRD2/n12 ), .CK(n5307), .Q(n53268)
         );
  DFF_X1 \DP/RegRD2/DOUT_reg[3]  ( .D(\DP/RegRD2/n11 ), .CK(n5307), .Q(n53267)
         );
  DFF_X1 \DP/RegRD2/DOUT_reg[4]  ( .D(\DP/RegRD2/n10 ), .CK(n5307), .Q(n53266)
         );
  DFF_X1 \DP/RegNPC2/DOUT_reg[0]  ( .D(n5275), .CK(n5307), .Q(n53451) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[1]  ( .D(n5276), .CK(n5307), .Q(n53452) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[2]  ( .D(n5277), .CK(n5307), .Q(n53453) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[3]  ( .D(n5278), .CK(n5307), .Q(n53454) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[4]  ( .D(n5279), .CK(n5307), .Q(n53455) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[5]  ( .D(n5280), .CK(n5307), .Q(n53456) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[6]  ( .D(n5281), .CK(n5307), .Q(n53457) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[7]  ( .D(n5282), .CK(n5307), .Q(n53458) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[8]  ( .D(n5283), .CK(n5307), .Q(n53459) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[9]  ( .D(n5284), .CK(n5307), .Q(n53460) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[10]  ( .D(n5285), .CK(n5307), .Q(n53461) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[11]  ( .D(n5286), .CK(n5307), .Q(n53462) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[12]  ( .D(n5287), .CK(n5307), .Q(n53463) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[13]  ( .D(n5288), .CK(n5307), .Q(n53464) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[14]  ( .D(n5289), .CK(n5307), .Q(n53465) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[15]  ( .D(n5290), .CK(n5307), .Q(n53466) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[16]  ( .D(n5291), .CK(n5307), .Q(n53467) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[17]  ( .D(n5292), .CK(n5307), .Q(n53468) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[18]  ( .D(n5293), .CK(n5307), .Q(n53469) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[19]  ( .D(n5294), .CK(n5307), .Q(n53470) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[20]  ( .D(n5295), .CK(n5307), .Q(n53471) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[21]  ( .D(n5296), .CK(n5307), .Q(n53472) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[22]  ( .D(n5297), .CK(n5307), .Q(n53473) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[23]  ( .D(n5298), .CK(n5307), .Q(n53474) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[24]  ( .D(n5299), .CK(n5307), .Q(n53475) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[25]  ( .D(n5300), .CK(n5307), .Q(n53476) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[26]  ( .D(n5301), .CK(n5307), .Q(n53477) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[27]  ( .D(n5302), .CK(n5307), .Q(n53478) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[28]  ( .D(n5303), .CK(n5307), .Q(n53479) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[29]  ( .D(n5304), .CK(n5307), .Q(n53480) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[30]  ( .D(n5305), .CK(n5307), .Q(n53481) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[31]  ( .D(n5306), .CK(n5307), .Q(n53482) );
  DLH_X1 \DP/ALU0/s_LOGIC_reg[2]  ( .G(n53611), .D(n53759), .Q(
        \DP/ALU0/s_LOGIC[2] ) );
  DLH_X1 \DP/ALU0/s_LOGIC_reg[3]  ( .G(n53611), .D(n20899), .Q(
        \DP/ALU0/s_LOGIC[3] ) );
  DLH_X1 \DP/ALU0/s_ADD_SUB_reg  ( .G(\DP/ALU0/N20 ), .D(n53612), .Q(
        \DP/ALU0/s_ADD_SUB ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[0]  ( .G(\DP/ALU0/n112 ), .D(n3092), .Q(
        \DP/ALU0/S_B_LHI[0] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[1]  ( .G(\DP/ALU0/n112 ), .D(n3089), .Q(
        \DP/ALU0/S_B_LHI[1] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[2]  ( .G(\DP/ALU0/n112 ), .D(n3086), .Q(
        \DP/ALU0/S_B_LHI[2] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[3]  ( .G(\DP/ALU0/n112 ), .D(n3083), .Q(
        \DP/ALU0/S_B_LHI[3] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[4]  ( .G(\DP/ALU0/n112 ), .D(n3080), .Q(
        \DP/ALU0/S_B_LHI[4] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[5]  ( .G(\DP/ALU0/n112 ), .D(n3077), .Q(
        \DP/ALU0/S_B_LHI[5] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[6]  ( .G(\DP/ALU0/n112 ), .D(n3074), .Q(
        \DP/ALU0/S_B_LHI[6] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[7]  ( .G(\DP/ALU0/n112 ), .D(n3071), .Q(
        \DP/ALU0/S_B_LHI[7] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[8]  ( .G(\DP/ALU0/n112 ), .D(n3068), .Q(
        \DP/ALU0/S_B_LHI[8] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[9]  ( .G(\DP/ALU0/n112 ), .D(n3065), .Q(
        \DP/ALU0/S_B_LHI[9] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[10]  ( .G(\DP/ALU0/n112 ), .D(n3062), .Q(
        \DP/ALU0/S_B_LHI[10] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[11]  ( .G(\DP/ALU0/n112 ), .D(n3059), .Q(
        \DP/ALU0/S_B_LHI[11] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[12]  ( .G(\DP/ALU0/n112 ), .D(n3147), .Q(
        \DP/ALU0/S_B_LHI[12] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[13]  ( .G(\DP/ALU0/n112 ), .D(n3145), .Q(
        \DP/ALU0/S_B_LHI[13] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[14]  ( .G(\DP/ALU0/n112 ), .D(n3143), .Q(
        \DP/ALU0/S_B_LHI[14] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[15]  ( .G(\DP/ALU0/n112 ), .D(n3141), .Q(
        \DP/ALU0/S_B_LHI[15] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[0]  ( .G(n53818), .D(n3092), .Q(
        \DP/ALU0/S_B_MULT[0] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[2]  ( .G(n53818), .D(n3086), .Q(
        \DP/ALU0/S_B_MULT[2] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[4]  ( .G(n53818), .D(n3080), .Q(
        \DP/ALU0/S_B_MULT[4] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[6]  ( .G(n53818), .D(n3074), .Q(
        \DP/ALU0/S_B_MULT[6] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[8]  ( .G(n53818), .D(n3068), .Q(
        \DP/ALU0/S_B_MULT[8] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[10]  ( .G(n53818), .D(n3062), .Q(
        \DP/ALU0/S_B_MULT[10] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[12]  ( .G(n53818), .D(n3147), .Q(
        \DP/ALU0/S_B_MULT[12] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[14]  ( .G(n53818), .D(n3143), .Q(
        \DP/ALU0/S_B_MULT[14] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[15]  ( .G(n53818), .D(n3141), .Q(
        \DP/ALU0/S_B_MULT[15] ) );
  DLH_X1 \DP/ALU0/s_SHIFT_reg[0]  ( .G(n53816), .D(\DP/ALU0/n114 ), .Q(
        \DP/ALU0/s_SHIFT[0] ) );
  DLH_X1 \DP/ALU0/s_SHIFT_reg[1]  ( .G(n53613), .D(n5402), .Q(
        \DP/ALU0/s_SHIFT[1] ) );
  DLH_X1 \DP/ALU0/S_B_SHIFT_reg[0]  ( .G(n53613), .D(n3092), .Q(
        \DP/ALU0/S_B_SHIFT[0] ) );
  DLH_X1 \DP/ALU0/S_B_SHIFT_reg[1]  ( .G(n53816), .D(n3089), .Q(
        \DP/ALU0/S_B_SHIFT[1] ) );
  DLH_X1 \DP/ALU0/S_B_SHIFT_reg[2]  ( .G(n53613), .D(n3086), .Q(
        \DP/ALU0/S_B_SHIFT[2] ) );
  DLH_X1 \DP/ALU0/S_B_SHIFT_reg[3]  ( .G(n53613), .D(n3083), .Q(
        \DP/ALU0/S_B_SHIFT[3] ) );
  DLH_X1 \DP/ALU0/S_B_SHIFT_reg[4]  ( .G(n53613), .D(n3080), .Q(
        \DP/ALU0/S_B_SHIFT[4] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[0]  ( .G(n53816), .D(n3091), .Q(
        \DP/ALU0/s_A_SHIFT[0] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[1]  ( .G(n53816), .D(n3088), .Q(
        \DP/ALU0/s_A_SHIFT[1] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[2]  ( .G(n53816), .D(n3085), .Q(
        \DP/ALU0/s_A_SHIFT[2] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[3]  ( .G(n53816), .D(n3082), .Q(
        \DP/ALU0/s_A_SHIFT[3] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[4]  ( .G(n53816), .D(n3079), .Q(
        \DP/ALU0/s_A_SHIFT[4] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[5]  ( .G(n53613), .D(n3076), .Q(
        \DP/ALU0/s_A_SHIFT[5] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[6]  ( .G(n53613), .D(n3073), .Q(
        \DP/ALU0/s_A_SHIFT[6] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[7]  ( .G(n53816), .D(n3070), .Q(
        \DP/ALU0/s_A_SHIFT[7] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[8]  ( .G(n53816), .D(n3067), .Q(
        \DP/ALU0/s_A_SHIFT[8] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[9]  ( .G(n53816), .D(n3064), .Q(
        \DP/ALU0/s_A_SHIFT[9] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[10]  ( .G(n53816), .D(n3061), .Q(
        \DP/ALU0/s_A_SHIFT[10] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[11]  ( .G(n53816), .D(n3058), .Q(
        \DP/ALU0/s_A_SHIFT[11] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[12]  ( .G(n53816), .D(n3146), .Q(
        \DP/ALU0/s_A_SHIFT[12] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[13]  ( .G(n53816), .D(n3144), .Q(
        \DP/ALU0/s_A_SHIFT[13] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[14]  ( .G(n53816), .D(n3142), .Q(
        \DP/ALU0/s_A_SHIFT[14] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[15]  ( .G(n53816), .D(n3140), .Q(
        \DP/ALU0/s_A_SHIFT[15] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[16]  ( .G(n53816), .D(n3138), .Q(
        \DP/ALU0/s_A_SHIFT[16] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[17]  ( .G(n53816), .D(n3136), .Q(
        \DP/ALU0/s_A_SHIFT[17] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[18]  ( .G(n53613), .D(n3134), .Q(
        \DP/ALU0/s_A_SHIFT[18] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[19]  ( .G(n53613), .D(n3132), .Q(
        \DP/ALU0/s_A_SHIFT[19] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[20]  ( .G(n53816), .D(n3130), .Q(
        \DP/ALU0/s_A_SHIFT[20] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[21]  ( .G(n53613), .D(n3128), .Q(
        \DP/ALU0/s_A_SHIFT[21] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[22]  ( .G(n53816), .D(n3126), .Q(
        \DP/ALU0/s_A_SHIFT[22] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[23]  ( .G(n53816), .D(n3124), .Q(
        \DP/ALU0/s_A_SHIFT[23] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[24]  ( .G(n53816), .D(n3104), .Q(
        \DP/ALU0/s_A_SHIFT[24] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[25]  ( .G(n53613), .D(n3152), .Q(
        \DP/ALU0/s_A_SHIFT[25] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[26]  ( .G(n53613), .D(n3101), .Q(
        \DP/ALU0/s_A_SHIFT[26] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[27]  ( .G(n53613), .D(n3098), .Q(
        \DP/ALU0/s_A_SHIFT[27] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[28]  ( .G(n53816), .D(n3094), .Q(
        \DP/ALU0/s_A_SHIFT[28] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[29]  ( .G(n53816), .D(n3150), .Q(
        \DP/ALU0/s_A_SHIFT[29] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[30]  ( .G(n53816), .D(n3148), .Q(
        \DP/ALU0/s_A_SHIFT[30] ) );
  DLH_X1 \DP/ALU0/s_A_SHIFT_reg[31]  ( .G(n53816), .D(n3107), .Q(
        \DP/ALU0/s_A_SHIFT[31] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[0]  ( .G(n53611), .D(n3092), .Q(
        \DP/ALU0/S_B_LOGIC[0] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[1]  ( .G(n53611), .D(n3089), .Q(
        \DP/ALU0/S_B_LOGIC[1] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[2]  ( .G(n53611), .D(n3086), .Q(
        \DP/ALU0/S_B_LOGIC[2] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[3]  ( .G(n53611), .D(n3083), .Q(
        \DP/ALU0/S_B_LOGIC[3] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[4]  ( .G(n53611), .D(n3080), .Q(
        \DP/ALU0/S_B_LOGIC[4] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[5]  ( .G(n53611), .D(n3077), .Q(
        \DP/ALU0/S_B_LOGIC[5] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[6]  ( .G(n53611), .D(n3074), .Q(
        \DP/ALU0/S_B_LOGIC[6] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[7]  ( .G(n53611), .D(n3071), .Q(
        \DP/ALU0/S_B_LOGIC[7] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[8]  ( .G(n53611), .D(n3068), .Q(
        \DP/ALU0/S_B_LOGIC[8] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[9]  ( .G(n53611), .D(n3065), .Q(
        \DP/ALU0/S_B_LOGIC[9] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[10]  ( .G(n53611), .D(n3062), .Q(
        \DP/ALU0/S_B_LOGIC[10] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[11]  ( .G(n53611), .D(n3059), .Q(
        \DP/ALU0/S_B_LOGIC[11] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[12]  ( .G(n53611), .D(n3147), .Q(
        \DP/ALU0/S_B_LOGIC[12] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[13]  ( .G(n53611), .D(n3145), .Q(
        \DP/ALU0/S_B_LOGIC[13] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[14]  ( .G(n53611), .D(n3143), .Q(
        \DP/ALU0/S_B_LOGIC[14] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[15]  ( .G(n53611), .D(n3141), .Q(
        \DP/ALU0/S_B_LOGIC[15] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[16]  ( .G(n53611), .D(n3139), .Q(
        \DP/ALU0/S_B_LOGIC[16] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[17]  ( .G(n53611), .D(n3137), .Q(
        \DP/ALU0/S_B_LOGIC[17] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[18]  ( .G(n53611), .D(n3135), .Q(
        \DP/ALU0/S_B_LOGIC[18] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[19]  ( .G(n53611), .D(n3133), .Q(
        \DP/ALU0/S_B_LOGIC[19] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[20]  ( .G(n53611), .D(n3131), .Q(
        \DP/ALU0/S_B_LOGIC[20] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[21]  ( .G(n53611), .D(n3129), .Q(
        \DP/ALU0/S_B_LOGIC[21] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[22]  ( .G(n53611), .D(n3127), .Q(
        \DP/ALU0/S_B_LOGIC[22] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[23]  ( .G(n53611), .D(n3125), .Q(
        \DP/ALU0/S_B_LOGIC[23] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[24]  ( .G(n53611), .D(n3105), .Q(
        \DP/ALU0/S_B_LOGIC[24] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[25]  ( .G(n53611), .D(n3153), .Q(
        \DP/ALU0/S_B_LOGIC[25] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[26]  ( .G(n53611), .D(n3102), .Q(
        \DP/ALU0/S_B_LOGIC[26] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[27]  ( .G(n53611), .D(n3099), .Q(
        \DP/ALU0/S_B_LOGIC[27] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[28]  ( .G(n53611), .D(n3095), .Q(
        \DP/ALU0/S_B_LOGIC[28] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[29]  ( .G(n53611), .D(n3151), .Q(
        \DP/ALU0/S_B_LOGIC[29] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[30]  ( .G(n53611), .D(n3149), .Q(
        \DP/ALU0/S_B_LOGIC[30] ) );
  DLH_X1 \DP/ALU0/S_B_LOGIC_reg[31]  ( .G(n53611), .D(n3108), .Q(
        \DP/ALU0/S_B_LOGIC[31] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[0]  ( .G(n53611), .D(n3091), .Q(
        \DP/ALU0/s_A_LOGIC[0] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[1]  ( .G(n53611), .D(n3088), .Q(
        \DP/ALU0/s_A_LOGIC[1] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[2]  ( .G(n53611), .D(n3085), .Q(
        \DP/ALU0/s_A_LOGIC[2] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[3]  ( .G(n53611), .D(n3082), .Q(
        \DP/ALU0/s_A_LOGIC[3] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[4]  ( .G(n53611), .D(n3079), .Q(
        \DP/ALU0/s_A_LOGIC[4] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[5]  ( .G(n53611), .D(n3076), .Q(
        \DP/ALU0/s_A_LOGIC[5] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[6]  ( .G(n53611), .D(n3073), .Q(
        \DP/ALU0/s_A_LOGIC[6] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[7]  ( .G(n53611), .D(n3070), .Q(
        \DP/ALU0/s_A_LOGIC[7] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[8]  ( .G(n53611), .D(n3067), .Q(
        \DP/ALU0/s_A_LOGIC[8] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[9]  ( .G(n53611), .D(n3064), .Q(
        \DP/ALU0/s_A_LOGIC[9] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[10]  ( .G(n53611), .D(n3061), .Q(
        \DP/ALU0/s_A_LOGIC[10] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[11]  ( .G(n53611), .D(n3058), .Q(
        \DP/ALU0/s_A_LOGIC[11] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[12]  ( .G(n53611), .D(n3146), .Q(
        \DP/ALU0/s_A_LOGIC[12] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[13]  ( .G(n53611), .D(n3144), .Q(
        \DP/ALU0/s_A_LOGIC[13] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[14]  ( .G(n53611), .D(n3142), .Q(
        \DP/ALU0/s_A_LOGIC[14] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[15]  ( .G(n53611), .D(n3140), .Q(
        \DP/ALU0/s_A_LOGIC[15] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[16]  ( .G(n53611), .D(n3138), .Q(
        \DP/ALU0/s_A_LOGIC[16] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[17]  ( .G(n53611), .D(n3136), .Q(
        \DP/ALU0/s_A_LOGIC[17] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[18]  ( .G(n53611), .D(n3134), .Q(
        \DP/ALU0/s_A_LOGIC[18] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[19]  ( .G(n53611), .D(n3132), .Q(
        \DP/ALU0/s_A_LOGIC[19] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[20]  ( .G(n53611), .D(n3130), .Q(
        \DP/ALU0/s_A_LOGIC[20] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[21]  ( .G(n53611), .D(n3128), .Q(
        \DP/ALU0/s_A_LOGIC[21] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[22]  ( .G(n53611), .D(n3126), .Q(
        \DP/ALU0/s_A_LOGIC[22] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[23]  ( .G(n53611), .D(n3124), .Q(
        \DP/ALU0/s_A_LOGIC[23] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[24]  ( .G(n53611), .D(n3104), .Q(
        \DP/ALU0/s_A_LOGIC[24] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[25]  ( .G(n53611), .D(n3152), .Q(
        \DP/ALU0/s_A_LOGIC[25] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[26]  ( .G(n53611), .D(n3101), .Q(
        \DP/ALU0/s_A_LOGIC[26] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[27]  ( .G(n53611), .D(n3098), .Q(
        \DP/ALU0/s_A_LOGIC[27] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[28]  ( .G(n53611), .D(n3094), .Q(
        \DP/ALU0/s_A_LOGIC[28] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[29]  ( .G(n53611), .D(n3150), .Q(
        \DP/ALU0/s_A_LOGIC[29] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[30]  ( .G(n53611), .D(n3148), .Q(
        \DP/ALU0/s_A_LOGIC[30] ) );
  DLH_X1 \DP/ALU0/s_A_LOGIC_reg[31]  ( .G(n53611), .D(n3107), .Q(
        \DP/ALU0/s_A_LOGIC[31] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[0]  ( .G(\DP/ALU0/N20 ), .D(n3092), .Q(
        \DP/ALU0/S_B_ADDER[0] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[1]  ( .G(\DP/ALU0/N20 ), .D(n3089), .Q(
        \DP/ALU0/S_B_ADDER[1] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[2]  ( .G(\DP/ALU0/N20 ), .D(n3086), .Q(
        \DP/ALU0/S_B_ADDER[2] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[3]  ( .G(\DP/ALU0/N20 ), .D(n3083), .Q(
        \DP/ALU0/S_B_ADDER[3] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[4]  ( .G(\DP/ALU0/N20 ), .D(n3080), .Q(
        \DP/ALU0/S_B_ADDER[4] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[5]  ( .G(\DP/ALU0/N20 ), .D(n3077), .Q(
        \DP/ALU0/S_B_ADDER[5] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[6]  ( .G(\DP/ALU0/N20 ), .D(n3074), .Q(
        \DP/ALU0/S_B_ADDER[6] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[7]  ( .G(\DP/ALU0/N20 ), .D(n3071), .Q(
        \DP/ALU0/S_B_ADDER[7] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[8]  ( .G(\DP/ALU0/N20 ), .D(n3068), .Q(
        \DP/ALU0/S_B_ADDER[8] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[9]  ( .G(\DP/ALU0/N20 ), .D(n3065), .Q(
        \DP/ALU0/S_B_ADDER[9] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[10]  ( .G(\DP/ALU0/N20 ), .D(n3062), .Q(
        \DP/ALU0/S_B_ADDER[10] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[11]  ( .G(\DP/ALU0/N20 ), .D(n3059), .Q(
        \DP/ALU0/S_B_ADDER[11] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[12]  ( .G(\DP/ALU0/N20 ), .D(n3147), .Q(
        \DP/ALU0/S_B_ADDER[12] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[13]  ( .G(\DP/ALU0/N20 ), .D(n3145), .Q(
        \DP/ALU0/S_B_ADDER[13] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[14]  ( .G(\DP/ALU0/N20 ), .D(n3143), .Q(
        \DP/ALU0/S_B_ADDER[14] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[15]  ( .G(\DP/ALU0/N20 ), .D(n3141), .Q(
        \DP/ALU0/S_B_ADDER[15] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[16]  ( .G(\DP/ALU0/N20 ), .D(n3139), .Q(
        \DP/ALU0/S_B_ADDER[16] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[17]  ( .G(\DP/ALU0/N20 ), .D(n3137), .Q(
        \DP/ALU0/S_B_ADDER[17] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[18]  ( .G(\DP/ALU0/N20 ), .D(n3135), .Q(
        \DP/ALU0/S_B_ADDER[18] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[19]  ( .G(\DP/ALU0/N20 ), .D(n3133), .Q(
        \DP/ALU0/S_B_ADDER[19] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[20]  ( .G(\DP/ALU0/N20 ), .D(n3131), .Q(
        \DP/ALU0/S_B_ADDER[20] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[21]  ( .G(\DP/ALU0/N20 ), .D(n3129), .Q(
        \DP/ALU0/S_B_ADDER[21] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[22]  ( .G(\DP/ALU0/N20 ), .D(n3127), .Q(
        \DP/ALU0/S_B_ADDER[22] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[23]  ( .G(\DP/ALU0/N20 ), .D(n3125), .Q(
        \DP/ALU0/S_B_ADDER[23] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[24]  ( .G(\DP/ALU0/N20 ), .D(n3105), .Q(
        \DP/ALU0/S_B_ADDER[24] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[25]  ( .G(\DP/ALU0/N20 ), .D(n3153), .Q(
        \DP/ALU0/S_B_ADDER[25] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[26]  ( .G(\DP/ALU0/N20 ), .D(n3102), .Q(
        \DP/ALU0/S_B_ADDER[26] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[27]  ( .G(\DP/ALU0/N20 ), .D(n3099), .Q(
        \DP/ALU0/S_B_ADDER[27] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[28]  ( .G(\DP/ALU0/N20 ), .D(n3095), .Q(
        \DP/ALU0/S_B_ADDER[28] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[29]  ( .G(\DP/ALU0/N20 ), .D(n3151), .Q(
        \DP/ALU0/S_B_ADDER[29] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[30]  ( .G(\DP/ALU0/N20 ), .D(n3149), .Q(
        \DP/ALU0/S_B_ADDER[30] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[31]  ( .G(\DP/ALU0/N20 ), .D(n3108), .Q(
        \DP/ALU0/S_B_ADDER[31] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[0]  ( .G(\DP/ALU0/N20 ), .D(n3091), .Q(
        \DP/ALU0/s_A_ADDER[0] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[1]  ( .G(\DP/ALU0/N20 ), .D(n3088), .Q(
        \DP/ALU0/s_A_ADDER[1] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[2]  ( .G(\DP/ALU0/N20 ), .D(n3085), .Q(
        \DP/ALU0/s_A_ADDER[2] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[3]  ( .G(\DP/ALU0/N20 ), .D(n3082), .Q(
        \DP/ALU0/s_A_ADDER[3] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[4]  ( .G(\DP/ALU0/N20 ), .D(n3079), .Q(
        \DP/ALU0/s_A_ADDER[4] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[5]  ( .G(\DP/ALU0/N20 ), .D(n3076), .Q(
        \DP/ALU0/s_A_ADDER[5] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[6]  ( .G(\DP/ALU0/N20 ), .D(n3073), .Q(
        \DP/ALU0/s_A_ADDER[6] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[7]  ( .G(\DP/ALU0/N20 ), .D(n3070), .Q(
        \DP/ALU0/s_A_ADDER[7] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[8]  ( .G(\DP/ALU0/N20 ), .D(n3067), .Q(
        \DP/ALU0/s_A_ADDER[8] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[9]  ( .G(\DP/ALU0/N20 ), .D(n3064), .Q(
        \DP/ALU0/s_A_ADDER[9] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[10]  ( .G(\DP/ALU0/N20 ), .D(n3061), .Q(
        \DP/ALU0/s_A_ADDER[10] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[11]  ( .G(\DP/ALU0/N20 ), .D(n3058), .Q(
        \DP/ALU0/s_A_ADDER[11] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[12]  ( .G(\DP/ALU0/N20 ), .D(n3146), .Q(
        \DP/ALU0/s_A_ADDER[12] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[13]  ( .G(\DP/ALU0/N20 ), .D(n3144), .Q(
        \DP/ALU0/s_A_ADDER[13] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[14]  ( .G(\DP/ALU0/N20 ), .D(n3142), .Q(
        \DP/ALU0/s_A_ADDER[14] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[15]  ( .G(\DP/ALU0/N20 ), .D(n3140), .Q(
        \DP/ALU0/s_A_ADDER[15] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[16]  ( .G(\DP/ALU0/N20 ), .D(n3138), .Q(
        \DP/ALU0/s_A_ADDER[16] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[17]  ( .G(\DP/ALU0/N20 ), .D(n3136), .Q(
        \DP/ALU0/s_A_ADDER[17] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[18]  ( .G(\DP/ALU0/N20 ), .D(n3134), .Q(
        \DP/ALU0/s_A_ADDER[18] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[19]  ( .G(\DP/ALU0/N20 ), .D(n3132), .Q(
        \DP/ALU0/s_A_ADDER[19] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[20]  ( .G(\DP/ALU0/N20 ), .D(n3130), .Q(
        \DP/ALU0/s_A_ADDER[20] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[21]  ( .G(\DP/ALU0/N20 ), .D(n3128), .Q(
        \DP/ALU0/s_A_ADDER[21] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[22]  ( .G(\DP/ALU0/N20 ), .D(n3126), .Q(
        \DP/ALU0/s_A_ADDER[22] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[23]  ( .G(\DP/ALU0/N20 ), .D(n3124), .Q(
        \DP/ALU0/s_A_ADDER[23] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[24]  ( .G(\DP/ALU0/N20 ), .D(n3104), .Q(
        \DP/ALU0/s_A_ADDER[24] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[25]  ( .G(\DP/ALU0/N20 ), .D(n3152), .Q(
        \DP/ALU0/s_A_ADDER[25] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[26]  ( .G(\DP/ALU0/N20 ), .D(n3101), .Q(
        \DP/ALU0/s_A_ADDER[26] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[27]  ( .G(\DP/ALU0/N20 ), .D(n3098), .Q(
        \DP/ALU0/s_A_ADDER[27] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[28]  ( .G(\DP/ALU0/N20 ), .D(n3094), .Q(
        \DP/ALU0/s_A_ADDER[28] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[29]  ( .G(\DP/ALU0/N20 ), .D(n3150), .Q(
        \DP/ALU0/s_A_ADDER[29] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[30]  ( .G(\DP/ALU0/N20 ), .D(n3148), .Q(
        \DP/ALU0/s_A_ADDER[30] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[31]  ( .G(\DP/ALU0/N20 ), .D(n3107), .Q(
        \DP/ALU0/s_A_ADDER[31] ) );
  DLH_X1 \DP/ALU0/s_SIGN_reg  ( .G(n51572), .D(\DP/ALU0/N27 ), .Q(
        \DP/ALU0/s_SIGN ) );
  DFF_X1 \DP/RegALU3/DOUT_reg[10]  ( .D(\DP/RegALU3/n89 ), .CK(n4991), .Q(
        n53756), .QN(n49808) );
  DFF_X1 \DP/RegALU3/DOUT_reg[11]  ( .D(\DP/RegALU3/n88 ), .CK(n4991), .QN(
        n49843) );
  DFF_X1 \DP/RegALU3/DOUT_reg[13]  ( .D(\DP/RegALU3/n86 ), .CK(n4991), .QN(
        n49810) );
  DFF_X1 \DP/RegALU3/DOUT_reg[17]  ( .D(\DP/RegALU3/n82 ), .CK(n4991), .Q(
        n53707), .QN(n49844) );
  DFF_X1 \DP/RegALU3/DOUT_reg[19]  ( .D(\DP/RegALU3/n80 ), .CK(n4991), .Q(
        n53708), .QN(n49815) );
  DFF_X1 \DP/RegALU3/DOUT_reg[27]  ( .D(\DP/RegALU3/n72 ), .CK(n4991), .Q(
        n7623), .QN(n53672) );
  DFF_X1 \DP/RegME/DOUT_reg[0]  ( .D(n4927), .CK(n4991), .QN(n53279) );
  DFF_X1 \DP/RegME/DOUT_reg[1]  ( .D(n4928), .CK(n4991), .QN(n53329) );
  DFF_X1 \DP/RegME/DOUT_reg[2]  ( .D(n4929), .CK(n4991), .QN(n53343) );
  DFF_X1 \DP/RegME/DOUT_reg[3]  ( .D(n4930), .CK(n4991), .QN(n53345) );
  DFF_X1 \DP/RegME/DOUT_reg[4]  ( .D(n4931), .CK(n4991), .QN(n53349) );
  DFF_X1 \DP/RegME/DOUT_reg[5]  ( .D(n4932), .CK(n4991), .QN(n53353) );
  DFF_X1 \DP/RegME/DOUT_reg[6]  ( .D(n4933), .CK(n4991), .QN(n53357) );
  DFF_X1 \DP/RegME/DOUT_reg[7]  ( .D(n4934), .CK(n4991), .QN(n53596) );
  DFF_X1 \DP/RegME/DOUT_reg[8]  ( .D(n4935), .CK(n4991), .QN(n53362) );
  DFF_X1 \DP/RegME/DOUT_reg[9]  ( .D(n4936), .CK(n4991), .QN(n53365) );
  DFF_X1 \DP/RegME/DOUT_reg[10]  ( .D(n4937), .CK(n4991), .QN(n53289) );
  DFF_X1 \DP/RegME/DOUT_reg[11]  ( .D(n4938), .CK(n4991), .QN(n53296) );
  DFF_X1 \DP/RegME/DOUT_reg[12]  ( .D(n4939), .CK(n4991), .QN(n53302) );
  DFF_X1 \DP/RegME/DOUT_reg[13]  ( .D(n4940), .CK(n4991), .QN(n53308) );
  DFF_X1 \DP/RegME/DOUT_reg[14]  ( .D(n4941), .CK(n4991), .QN(n53314) );
  DFF_X1 \DP/RegME/DOUT_reg[15]  ( .D(n4942), .CK(n4991), .QN(n53317) );
  DFF_X1 \DP/RegME/DOUT_reg[16]  ( .D(n4943), .CK(n4991), .QN(n53318) );
  DFF_X1 \DP/RegME/DOUT_reg[17]  ( .D(n4944), .CK(n4991), .QN(n53328) );
  DFF_X1 \DP/RegME/DOUT_reg[18]  ( .D(n4945), .CK(n4991), .QN(n53342) );
  DFF_X1 \DP/RegME/DOUT_reg[19]  ( .D(n4946), .CK(n4991), .QN(n53344) );
  DFF_X1 \DP/RegME/DOUT_reg[20]  ( .D(n4947), .CK(n4991), .QN(n53348) );
  DFF_X1 \DP/RegME/DOUT_reg[21]  ( .D(n4948), .CK(n4991), .QN(n53352) );
  DFF_X1 \DP/RegME/DOUT_reg[22]  ( .D(n4949), .CK(n4991), .QN(n53356) );
  DFF_X1 \DP/RegME/DOUT_reg[23]  ( .D(n4950), .CK(n4991), .QN(n53595) );
  DFF_X1 \DP/RegME/DOUT_reg[24]  ( .D(n4951), .CK(n4991), .QN(n53278) );
  DFF_X1 \DP/RegME/DOUT_reg[25]  ( .D(n4952), .CK(n4991), .QN(n53327) );
  DFF_X1 \DP/RegME/DOUT_reg[26]  ( .D(n4953), .CK(n4991), .QN(n53288) );
  DFF_X1 \DP/RegME/DOUT_reg[27]  ( .D(n4954), .CK(n4991), .QN(n53293) );
  DFF_X1 \DP/RegME/DOUT_reg[28]  ( .D(n4955), .CK(n4991), .QN(n53299) );
  DFF_X1 \DP/RegME/DOUT_reg[29]  ( .D(n4956), .CK(n4991), .QN(n53305) );
  DFF_X1 \DP/RegME/DOUT_reg[30]  ( .D(n4957), .CK(n4991), .QN(n53311) );
  DFF_X1 \DP/RegME/DOUT_reg[31]  ( .D(n4958), .CK(n4991), .QN(n53290) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[0]  ( .D(n4959), .CK(n4991), .QN(n53725) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[1]  ( .D(n4960), .CK(n4991), .QN(n53718) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[2]  ( .D(n4961), .CK(n4991), .QN(n53719) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[3]  ( .D(n4962), .CK(n4991), .QN(n53728) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[4]  ( .D(n4963), .CK(n4991), .QN(n53711) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[5]  ( .D(n4964), .CK(n4991), .QN(n53715) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[6]  ( .D(n4965), .CK(n4991), .QN(n53729) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[7]  ( .D(n4966), .CK(n4991), .QN(n53742) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[8]  ( .D(n4967), .CK(n4991), .QN(n53740) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[9]  ( .D(n4968), .CK(n4991), .QN(n53714) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[10]  ( .D(n4969), .CK(n4991), .QN(n53712) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[11]  ( .D(n4970), .CK(n4991), .QN(n53726) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[12]  ( .D(n4971), .CK(n4991), .QN(n53721) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[13]  ( .D(n4972), .CK(n4991), .QN(n53723) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[14]  ( .D(n4973), .CK(n4991), .QN(n53732) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[15]  ( .D(n4974), .CK(n4991), .QN(n53722) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[16]  ( .D(n4975), .CK(n4991), .QN(n53730) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[17]  ( .D(n4976), .CK(n4991), .QN(n53720) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[18]  ( .D(n4977), .CK(n4991), .QN(n53739) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[19]  ( .D(n4978), .CK(n4991), .QN(n53716) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[20]  ( .D(n4979), .CK(n4991), .QN(n53738) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[21]  ( .D(n4980), .CK(n4991), .QN(n53731) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[22]  ( .D(n4981), .CK(n4991), .QN(n53733) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[23]  ( .D(n4982), .CK(n4991), .QN(n53735) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[24]  ( .D(n4983), .CK(n4991), .QN(n53724) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[25]  ( .D(n4984), .CK(n4991), .QN(n53727) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[26]  ( .D(n4985), .CK(n4991), .QN(n53713) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[27]  ( .D(n4986), .CK(n4991), .QN(n53737) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[28]  ( .D(n4987), .CK(n4991), .QN(n53734) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[29]  ( .D(n4988), .CK(n4991), .QN(n53736) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[30]  ( .D(n4989), .CK(n4991), .QN(n53717) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[31]  ( .D(n4990), .CK(n4991), .QN(n53741) );
  DFF_X1 \DP/RegLMD/DOUT_reg[0]  ( .D(n4992), .CK(n5088), .QN(n53282) );
  DFF_X1 \DP/RegLMD/DOUT_reg[1]  ( .D(n4993), .CK(n5088), .QN(n53330) );
  DFF_X1 \DP/RegLMD/DOUT_reg[2]  ( .D(n4994), .CK(n5088), .QN(n53340) );
  DFF_X1 \DP/RegLMD/DOUT_reg[3]  ( .D(n4995), .CK(n5088), .QN(n53346) );
  DFF_X1 \DP/RegLMD/DOUT_reg[4]  ( .D(n4996), .CK(n5088), .QN(n53350) );
  DFF_X1 \DP/RegLMD/DOUT_reg[5]  ( .D(n4997), .CK(n5088), .QN(n53354) );
  DFF_X1 \DP/RegLMD/DOUT_reg[6]  ( .D(n4998), .CK(n5088), .QN(n53358) );
  DFF_X1 \DP/RegLMD/DOUT_reg[8]  ( .D(n5000), .CK(n5088), .Q(n53360) );
  DFF_X1 \DP/RegLMD/DOUT_reg[9]  ( .D(n5001), .CK(n5088), .Q(n53363) );
  DFF_X1 \DP/RegLMD/DOUT_reg[10]  ( .D(n5002), .CK(n5088), .Q(n53284) );
  DFF_X1 \DP/RegLMD/DOUT_reg[11]  ( .D(n5003), .CK(n5088), .Q(n53295) );
  DFF_X1 \DP/RegLMD/DOUT_reg[12]  ( .D(n5004), .CK(n5088), .Q(n53301) );
  DFF_X1 \DP/RegLMD/DOUT_reg[13]  ( .D(n5005), .CK(n5088), .Q(n53306) );
  DFF_X1 \DP/RegLMD/DOUT_reg[14]  ( .D(n5006), .CK(n5088), .Q(n53312) );
  DFF_X1 \DP/RegLMD/DOUT_reg[15]  ( .D(n5007), .CK(n5088), .Q(n53315) );
  DFF_X1 \DP/RegLMD/DOUT_reg[16]  ( .D(n5008), .CK(n5088), .QN(n53280) );
  DFF_X1 \DP/RegLMD/DOUT_reg[17]  ( .D(n5009), .CK(n5088), .QN(n53319) );
  DFF_X1 \DP/RegLMD/DOUT_reg[18]  ( .D(n5010), .CK(n5088), .QN(n53321) );
  DFF_X1 \DP/RegLMD/DOUT_reg[19]  ( .D(n5011), .CK(n5088), .QN(n53324) );
  DFF_X1 \DP/RegLMD/DOUT_reg[20]  ( .D(n5012), .CK(n5088), .QN(n53333) );
  DFF_X1 \DP/RegLMD/DOUT_reg[21]  ( .D(n5013), .CK(n5088), .QN(n53335) );
  DFF_X1 \DP/RegLMD/DOUT_reg[22]  ( .D(n5014), .CK(n5088), .QN(n53337) );
  DFF_X1 \DP/RegLMD/DOUT_reg[23]  ( .D(n5015), .CK(n5088), .QN(n53339) );
  DFF_X1 \DP/RegLMD/DOUT_reg[24]  ( .D(n5016), .CK(n5088), .QN(n53277) );
  DFF_X1 \DP/RegLMD/DOUT_reg[25]  ( .D(n5017), .CK(n5088), .QN(n53326) );
  DFF_X1 \DP/RegLMD/DOUT_reg[26]  ( .D(n5018), .CK(n5088), .QN(n53287) );
  DFF_X1 \DP/RegLMD/DOUT_reg[27]  ( .D(n5019), .CK(n5088), .QN(n53292) );
  DFF_X1 \DP/RegLMD/DOUT_reg[28]  ( .D(n5020), .CK(n5088), .QN(n53298) );
  DFF_X1 \DP/RegLMD/DOUT_reg[29]  ( .D(n5021), .CK(n5088), .QN(n53304) );
  DFF_X1 \DP/RegLMD/DOUT_reg[30]  ( .D(n5022), .CK(n5088), .QN(n53310) );
  DFF_X1 \DP/RegLMD/DOUT_reg[31]  ( .D(n5023), .CK(n5088), .QN(n53260) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[0]  ( .D(n5024), .CK(n5088), .QN(n53367) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[1]  ( .D(n5025), .CK(n5088), .QN(n53366) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[3]  ( .D(n5027), .CK(n5088), .QN(n49939) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[5]  ( .D(n5029), .CK(n5088), .Q(n53372) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[6]  ( .D(n5030), .CK(n5088), .QN(n53414) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[7]  ( .D(n5031), .CK(n5088), .Q(n49955) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[13]  ( .D(n5037), .CK(n5088), .Q(n49952) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[19]  ( .D(n5043), .CK(n5088), .Q(n53381) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[20]  ( .D(n5044), .CK(n5088), .QN(n53376) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[21]  ( .D(n5045), .CK(n5088), .Q(n53380) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[23]  ( .D(n5047), .CK(n5088), .Q(n53378), .QN(
        n53789) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[25]  ( .D(n5049), .CK(n5088), .Q(n53374) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[31]  ( .D(n5055), .CK(n5088), .Q(n53388) );
  DFF_X1 \DP/RegALU4/DOUT_reg[0]  ( .D(n5056), .CK(n5088), .QN(n53283) );
  DFF_X1 \DP/RegALU4/DOUT_reg[1]  ( .D(n5057), .CK(n5088), .QN(n53331) );
  DFF_X1 \DP/RegALU4/DOUT_reg[2]  ( .D(n5058), .CK(n5088), .QN(n53341) );
  DFF_X1 \DP/RegALU4/DOUT_reg[3]  ( .D(n5059), .CK(n5088), .QN(n53347) );
  DFF_X1 \DP/RegALU4/DOUT_reg[4]  ( .D(n5060), .CK(n5088), .QN(n53351) );
  DFF_X1 \DP/RegALU4/DOUT_reg[5]  ( .D(n5061), .CK(n5088), .QN(n53355) );
  DFF_X1 \DP/RegALU4/DOUT_reg[6]  ( .D(n5062), .CK(n5088), .QN(n53359) );
  DFF_X1 \DP/RegALU4/DOUT_reg[7]  ( .D(n5063), .CK(n5088), .QN(n53371) );
  DFF_X1 \DP/RegALU4/DOUT_reg[8]  ( .D(n5064), .CK(n5088), .QN(n53361) );
  DFF_X1 \DP/RegALU4/DOUT_reg[9]  ( .D(n5065), .CK(n5088), .QN(n53364) );
  DFF_X1 \DP/RegALU4/DOUT_reg[10]  ( .D(n5066), .CK(n5088), .QN(n53285) );
  DFF_X1 \DP/RegALU4/DOUT_reg[11]  ( .D(n5067), .CK(n5088), .QN(n53294) );
  DFF_X1 \DP/RegALU4/DOUT_reg[12]  ( .D(n5068), .CK(n5088), .QN(n53300) );
  DFF_X1 \DP/RegALU4/DOUT_reg[13]  ( .D(n5069), .CK(n5088), .QN(n53307) );
  DFF_X1 \DP/RegALU4/DOUT_reg[14]  ( .D(n5070), .CK(n5088), .QN(n53313) );
  DFF_X1 \DP/RegALU4/DOUT_reg[15]  ( .D(n5071), .CK(n5088), .QN(n53316) );
  DFF_X1 \DP/RegALU4/DOUT_reg[16]  ( .D(n5072), .CK(n5088), .Q(n53281) );
  DFF_X1 \DP/RegALU4/DOUT_reg[17]  ( .D(n5073), .CK(n5088), .Q(n53320) );
  DFF_X1 \DP/RegALU4/DOUT_reg[18]  ( .D(n5074), .CK(n5088), .Q(n53322) );
  DFF_X1 \DP/RegALU4/DOUT_reg[19]  ( .D(n5075), .CK(n5088), .Q(n53323) );
  DFF_X1 \DP/RegALU4/DOUT_reg[20]  ( .D(n5076), .CK(n5088), .Q(n53332) );
  DFF_X1 \DP/RegALU4/DOUT_reg[21]  ( .D(n5077), .CK(n5088), .Q(n53334) );
  DFF_X1 \DP/RegALU4/DOUT_reg[22]  ( .D(n5078), .CK(n5088), .Q(n53336) );
  DFF_X1 \DP/RegALU4/DOUT_reg[23]  ( .D(n5079), .CK(n5088), .Q(n53338) );
  DFF_X1 \DP/RegALU4/DOUT_reg[24]  ( .D(n5080), .CK(n5088), .Q(n53276) );
  DFF_X1 \DP/RegALU4/DOUT_reg[25]  ( .D(n5081), .CK(n5088), .Q(n53325) );
  DFF_X1 \DP/RegALU4/DOUT_reg[26]  ( .D(n5082), .CK(n5088), .Q(n53286) );
  DFF_X1 \DP/RegALU4/DOUT_reg[27]  ( .D(n5083), .CK(n5088), .Q(n53291) );
  DFF_X1 \DP/RegALU4/DOUT_reg[28]  ( .D(n5084), .CK(n5088), .Q(n53297) );
  DFF_X1 \DP/RegALU4/DOUT_reg[29]  ( .D(n5085), .CK(n5088), .Q(n53303) );
  DFF_X1 \DP/RegALU4/DOUT_reg[30]  ( .D(n5086), .CK(n5088), .Q(n53309) );
  DFF_X1 \DP/RegALU4/DOUT_reg[31]  ( .D(n5087), .CK(n5088), .Q(n53259) );
  DFF_X1 \DP/FU/RS2_EX_reg[0]  ( .D(n3253), .CK(n4923), .QN(n53273) );
  DFFR_X1 \DP/FU/RS2_ID_reg[0]  ( .D(w_RS2[0]), .CK(CLK), .RN(RST), .Q(n3253), 
        .QN(n7679) );
  DFFR_X1 \DP/FU/RS2_ID_reg[1]  ( .D(w_RS2[1]), .CK(CLK), .RN(RST), .Q(n18754), 
        .QN(n22592) );
  DFF_X1 \DP/FU/RS2_EX_reg[2]  ( .D(n3214), .CK(n4923), .Q(n53275) );
  DFFR_X1 \DP/FU/RS2_ID_reg[2]  ( .D(w_RS2[2]), .CK(CLK), .RN(RST), .Q(n3214), 
        .QN(n37948) );
  DFFR_X1 \DP/FU/RS2_ID_reg[3]  ( .D(w_RS2[3]), .CK(CLK), .RN(RST), .QN(n7286)
         );
  DFFR_X1 \DP/FU/RS2_ID_reg[4]  ( .D(w_RS2[4]), .CK(CLK), .RN(RST), .QN(n53261) );
  DFFR_X1 \DP/FU/RS1_ID_reg[0]  ( .D(\DP/IMMS26[21] ), .CK(CLK), .RN(RST), .Q(
        n53758), .QN(n53264) );
  DFFR_X1 \DP/FU/RS1_ID_reg[1]  ( .D(\DP/IMMS26[22] ), .CK(CLK), .RN(RST), 
        .QN(n49913) );
  DFFR_X1 \DP/FU/RS1_ID_reg[2]  ( .D(\DP/IMMS26[23] ), .CK(CLK), .RN(RST), 
        .QN(n53265) );
  DFFR_X1 \DP/FU/RS1_ID_reg[3]  ( .D(\DP/IMMS26[24] ), .CK(CLK), .RN(RST), .Q(
        n53754), .QN(n53263) );
  DFFR_X1 \DP/FU/RS1_ID_reg[4]  ( .D(\DP/IMMS26[25] ), .CK(CLK), .RN(RST), 
        .QN(n49917) );
  SNPS_CLOCK_GATE_HIGH_DLX_WIDTH32_0 \clk_gate_DP/RegNPC2/DOUT_reg  ( .CLK(CLK), .EN(\DP/RegRD2/n7 ), .ENCLK(n5307), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_DLX_WIDTH32_1 \clk_gate_DP/RegNPC1/DOUT_reg  ( .CLK(CLK), .EN(n897), .ENCLK(n5185), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_DLX_WIDTH32_2 \clk_gate_DP/RegALU4/DOUT_reg  ( .CLK(CLK), .EN(\DP/RegRD4/n7 ), .ENCLK(n5088), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_DLX_WIDTH32_3 \clk_gate_DP/RegNPC3/DOUT_reg  ( .CLK(CLK), .EN(n5463), .ENCLK(n4991), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_DLX_WIDTH32_4 \clk_gate_DP/FU/RS2_EX_reg  ( .CLK(CLK), 
        .EN(RST), .ENCLK(n4923), .TE(1'b0) );
  FA_X1 \intadd_0/U28  ( .A(n51773), .B(\intadd_0/B[0] ), .CI(\intadd_0/CI ), 
        .CO(\intadd_0/n27 ), .S(\intadd_0/SUM[0] ) );
  FA_X1 \intadd_0/U27  ( .A(n51774), .B(\intadd_0/B[1] ), .CI(\intadd_0/n27 ), 
        .CO(\intadd_0/n26 ), .S(\intadd_0/SUM[1] ) );
  FA_X1 \intadd_0/U26  ( .A(n51775), .B(\intadd_0/B[2] ), .CI(\intadd_0/n26 ), 
        .CO(\intadd_0/n25 ), .S(\intadd_0/SUM[2] ) );
  FA_X1 \intadd_0/U25  ( .A(n51776), .B(\intadd_0/B[3] ), .CI(\intadd_0/n25 ), 
        .CO(\intadd_0/n24 ), .S(\intadd_0/SUM[3] ) );
  FA_X1 \intadd_0/U24  ( .A(n51777), .B(\intadd_0/B[4] ), .CI(\intadd_0/n24 ), 
        .CO(\intadd_0/n23 ), .S(\intadd_0/SUM[4] ) );
  FA_X1 \intadd_0/U23  ( .A(n51778), .B(\intadd_0/B[5] ), .CI(\intadd_0/n23 ), 
        .CO(\intadd_0/n22 ), .S(\intadd_0/SUM[5] ) );
  FA_X1 \intadd_0/U22  ( .A(n51779), .B(\intadd_0/B[6] ), .CI(\intadd_0/n22 ), 
        .CO(\intadd_0/n21 ), .S(\intadd_0/SUM[6] ) );
  FA_X1 \intadd_0/U21  ( .A(n51780), .B(\intadd_0/B[7] ), .CI(\intadd_0/n21 ), 
        .CO(\intadd_0/n20 ), .S(\intadd_0/SUM[7] ) );
  FA_X1 \intadd_0/U20  ( .A(n51781), .B(\intadd_0/B[8] ), .CI(\intadd_0/n20 ), 
        .CO(\intadd_0/n19 ), .S(\intadd_0/SUM[8] ) );
  FA_X1 \intadd_0/U19  ( .A(n51782), .B(\intadd_0/B[9] ), .CI(\intadd_0/n19 ), 
        .CO(\intadd_0/n18 ), .S(\intadd_0/SUM[9] ) );
  FA_X1 \intadd_0/U18  ( .A(n51783), .B(\intadd_0/B[10] ), .CI(\intadd_0/n18 ), 
        .CO(\intadd_0/n17 ), .S(\intadd_0/SUM[10] ) );
  FA_X1 \intadd_0/U17  ( .A(n51784), .B(\intadd_0/B[11] ), .CI(\intadd_0/n17 ), 
        .CO(\intadd_0/n16 ), .S(\intadd_0/SUM[11] ) );
  FA_X1 \intadd_0/U16  ( .A(n51785), .B(\intadd_0/B[12] ), .CI(\intadd_0/n16 ), 
        .CO(\intadd_0/n15 ), .S(\intadd_0/SUM[12] ) );
  FA_X1 \intadd_0/U15  ( .A(n51786), .B(\intadd_0/B[13] ), .CI(\intadd_0/n15 ), 
        .CO(\intadd_0/n14 ), .S(\intadd_0/SUM[13] ) );
  FA_X1 \intadd_0/U14  ( .A(n51787), .B(\intadd_0/B[14] ), .CI(\intadd_0/n14 ), 
        .CO(\intadd_0/n13 ), .S(\intadd_0/SUM[14] ) );
  FA_X1 \intadd_0/U13  ( .A(n51788), .B(\intadd_0/B[15] ), .CI(\intadd_0/n13 ), 
        .CO(\intadd_0/n12 ), .S(\intadd_0/SUM[15] ) );
  FA_X1 \intadd_0/U12  ( .A(n51789), .B(\intadd_0/B[16] ), .CI(\intadd_0/n12 ), 
        .CO(\intadd_0/n11 ), .S(\intadd_0/SUM[16] ) );
  FA_X1 \intadd_0/U11  ( .A(n51790), .B(\intadd_0/B[17] ), .CI(\intadd_0/n11 ), 
        .CO(\intadd_0/n10 ), .S(\intadd_0/SUM[17] ) );
  FA_X1 \intadd_0/U10  ( .A(n51791), .B(\intadd_0/B[18] ), .CI(\intadd_0/n10 ), 
        .CO(\intadd_0/n9 ), .S(\intadd_0/SUM[18] ) );
  FA_X1 \intadd_0/U9  ( .A(n51792), .B(\intadd_0/B[19] ), .CI(\intadd_0/n9 ), 
        .CO(\intadd_0/n8 ), .S(\intadd_0/SUM[19] ) );
  FA_X1 \intadd_0/U8  ( .A(n51793), .B(\intadd_0/B[20] ), .CI(\intadd_0/n8 ), 
        .CO(\intadd_0/n7 ), .S(\intadd_0/SUM[20] ) );
  FA_X1 \intadd_0/U7  ( .A(n51794), .B(\intadd_0/B[21] ), .CI(\intadd_0/n7 ), 
        .CO(\intadd_0/n6 ), .S(\intadd_0/SUM[21] ) );
  FA_X1 \intadd_0/U6  ( .A(n51795), .B(\intadd_0/B[22] ), .CI(\intadd_0/n6 ), 
        .CO(\intadd_0/n5 ), .S(\intadd_0/SUM[22] ) );
  FA_X1 \intadd_0/U5  ( .A(n51796), .B(\intadd_0/B[23] ), .CI(\intadd_0/n5 ), 
        .CO(\intadd_0/n4 ), .S(\intadd_0/SUM[23] ) );
  FA_X1 \intadd_0/U4  ( .A(n51797), .B(\intadd_0/B[24] ), .CI(\intadd_0/n4 ), 
        .CO(\intadd_0/n3 ), .S(\intadd_0/SUM[24] ) );
  FA_X1 \intadd_0/U3  ( .A(n51798), .B(\intadd_0/B[25] ), .CI(\intadd_0/n3 ), 
        .CO(\intadd_0/n2 ), .S(\intadd_0/SUM[25] ) );
  FA_X1 \intadd_0/U2  ( .A(n51799), .B(\intadd_0/B[26] ), .CI(\intadd_0/n2 ), 
        .CO(\intadd_0/n1 ), .S(\intadd_0/SUM[26] ) );
  FA_X1 \intadd_1/U14  ( .A(\intadd_1/A[0] ), .B(n51666), .CI(\intadd_1/CI ), 
        .CO(\intadd_1/n13 ), .S(\intadd_1/SUM[0] ) );
  FA_X1 \intadd_1/U13  ( .A(n51662), .B(\intadd_1/B[1] ), .CI(\intadd_1/n13 ), 
        .CO(\intadd_1/n12 ), .S(\intadd_1/SUM[1] ) );
  FA_X1 \intadd_1/U12  ( .A(n51658), .B(\intadd_1/B[2] ), .CI(\intadd_1/n12 ), 
        .CO(\intadd_1/n11 ), .S(\intadd_1/SUM[2] ) );
  FA_X1 \intadd_1/U11  ( .A(n51654), .B(\intadd_1/B[3] ), .CI(\intadd_1/n11 ), 
        .CO(\intadd_1/n10 ), .S(\intadd_1/SUM[3] ) );
  FA_X1 \intadd_1/U10  ( .A(n51651), .B(\intadd_1/B[4] ), .CI(\intadd_1/n10 ), 
        .CO(\intadd_1/n9 ), .S(\intadd_1/SUM[4] ) );
  FA_X1 \intadd_1/U9  ( .A(n51648), .B(\intadd_1/B[5] ), .CI(\intadd_1/n9 ), 
        .CO(\intadd_1/n8 ), .S(\intadd_1/SUM[5] ) );
  FA_X1 \intadd_1/U8  ( .A(n51646), .B(\intadd_1/B[6] ), .CI(\intadd_1/n8 ), 
        .CO(\intadd_1/n7 ), .S(\intadd_1/SUM[6] ) );
  FA_X1 \intadd_1/U7  ( .A(n51644), .B(\intadd_1/B[7] ), .CI(\intadd_1/n7 ), 
        .CO(\intadd_1/n6 ), .S(\intadd_1/SUM[7] ) );
  FA_X1 \intadd_1/U6  ( .A(n51643), .B(\intadd_1/B[8] ), .CI(\intadd_1/n6 ), 
        .CO(\intadd_1/n5 ), .S(\intadd_1/SUM[8] ) );
  FA_X1 \intadd_1/U5  ( .A(n51642), .B(\intadd_1/B[9] ), .CI(\intadd_1/n5 ), 
        .CO(\intadd_1/n4 ), .S(\intadd_1/SUM[9] ) );
  FA_X1 \intadd_1/U4  ( .A(n51641), .B(\intadd_1/B[10] ), .CI(\intadd_1/n4 ), 
        .CO(\intadd_1/n3 ), .S(\intadd_1/SUM[10] ) );
  FA_X1 \intadd_1/U3  ( .A(\intadd_1/A[11] ), .B(\intadd_1/B[11] ), .CI(
        \intadd_1/n3 ), .CO(\intadd_1/n2 ), .S(\intadd_1/SUM[11] ) );
  FA_X1 \intadd_1/U2  ( .A(\intadd_1/A[12] ), .B(\intadd_1/B[12] ), .CI(
        \intadd_1/n2 ), .CO(\intadd_1/n1 ), .S(\intadd_1/SUM[12] ) );
  FA_X1 \intadd_2/U14  ( .A(\intadd_2/A[0] ), .B(\intadd_2/B[0] ), .CI(
        \intadd_2/CI ), .CO(\intadd_2/n13 ), .S(\intadd_2/SUM[0] ) );
  FA_X1 \intadd_2/U13  ( .A(\intadd_2/A[1] ), .B(\intadd_2/B[1] ), .CI(
        \intadd_2/n13 ), .CO(\intadd_2/n12 ), .S(\intadd_2/SUM[1] ) );
  FA_X1 \intadd_2/U12  ( .A(\intadd_2/A[2] ), .B(\intadd_2/B[2] ), .CI(
        \intadd_2/n12 ), .CO(\intadd_2/n11 ), .S(\intadd_2/SUM[2] ) );
  FA_X1 \intadd_2/U11  ( .A(\intadd_2/A[3] ), .B(\intadd_2/B[3] ), .CI(
        \intadd_2/n11 ), .CO(\intadd_2/n10 ), .S(\intadd_2/SUM[3] ) );
  FA_X1 \intadd_2/U10  ( .A(\intadd_2/A[4] ), .B(\intadd_2/B[4] ), .CI(
        \intadd_2/n10 ), .CO(\intadd_2/n9 ), .S(\intadd_2/SUM[4] ) );
  FA_X1 \intadd_2/U9  ( .A(\intadd_2/A[5] ), .B(\intadd_2/B[5] ), .CI(
        \intadd_2/n9 ), .CO(\intadd_2/n8 ), .S(\intadd_2/SUM[5] ) );
  FA_X1 \intadd_2/U8  ( .A(\intadd_2/A[6] ), .B(\intadd_2/B[6] ), .CI(
        \intadd_2/n8 ), .CO(\intadd_2/n7 ), .S(\intadd_2/SUM[6] ) );
  FA_X1 \intadd_2/U7  ( .A(\intadd_2/A[7] ), .B(\intadd_2/B[7] ), .CI(
        \intadd_2/n7 ), .CO(\intadd_2/n6 ), .S(\intadd_2/SUM[7] ) );
  FA_X1 \intadd_2/U6  ( .A(\intadd_2/A[8] ), .B(\intadd_2/B[8] ), .CI(
        \intadd_2/n6 ), .CO(\intadd_2/n5 ), .S(\intadd_2/SUM[8] ) );
  FA_X1 \intadd_2/U5  ( .A(\intadd_2/A[9] ), .B(\intadd_2/B[9] ), .CI(
        \intadd_2/n5 ), .CO(\intadd_2/n4 ), .S(\intadd_2/SUM[9] ) );
  FA_X1 \intadd_2/U4  ( .A(\intadd_2/A[10] ), .B(\intadd_2/B[10] ), .CI(
        \intadd_2/n4 ), .CO(\intadd_2/n3 ), .S(\intadd_2/SUM[10] ) );
  FA_X1 \intadd_2/U3  ( .A(\intadd_2/A[11] ), .B(\intadd_2/B[11] ), .CI(
        \intadd_2/n3 ), .CO(\intadd_2/n2 ), .S(\intadd_2/SUM[11] ) );
  FA_X1 \intadd_2/U2  ( .A(\intadd_2/A[12] ), .B(\intadd_2/B[12] ), .CI(
        \intadd_2/n2 ), .CO(\intadd_2/n1 ), .S(\intadd_2/SUM[12] ) );
  FA_X1 \intadd_3/U14  ( .A(\intadd_3/A[0] ), .B(\intadd_3/B[0] ), .CI(n51684), 
        .CO(\intadd_3/n13 ), .S(\intadd_3/SUM[0] ) );
  FA_X1 \intadd_3/U13  ( .A(\intadd_3/A[1] ), .B(n51680), .CI(\intadd_3/n13 ), 
        .CO(\intadd_3/n12 ), .S(\intadd_3/SUM[1] ) );
  FA_X1 \intadd_3/U12  ( .A(\intadd_3/A[2] ), .B(n51675), .CI(\intadd_3/n12 ), 
        .CO(\intadd_3/n11 ), .S(\intadd_2/CI ) );
  FA_X1 \intadd_3/U11  ( .A(\intadd_3/A[3] ), .B(n51671), .CI(\intadd_3/n11 ), 
        .CO(\intadd_3/n10 ), .S(\intadd_2/B[1] ) );
  FA_X1 \intadd_3/U10  ( .A(\intadd_3/A[4] ), .B(n51667), .CI(\intadd_3/n10 ), 
        .CO(\intadd_3/n9 ), .S(\intadd_2/B[2] ) );
  FA_X1 \intadd_3/U9  ( .A(\intadd_3/A[5] ), .B(n51663), .CI(\intadd_3/n9 ), 
        .CO(\intadd_3/n8 ), .S(\intadd_2/B[3] ) );
  FA_X1 \intadd_3/U8  ( .A(\intadd_3/A[6] ), .B(n51659), .CI(\intadd_3/n8 ), 
        .CO(\intadd_3/n7 ), .S(\intadd_2/B[4] ) );
  FA_X1 \intadd_3/U7  ( .A(\intadd_3/A[7] ), .B(n51655), .CI(\intadd_3/n7 ), 
        .CO(\intadd_3/n6 ), .S(\intadd_2/B[5] ) );
  FA_X1 \intadd_3/U6  ( .A(\intadd_3/A[8] ), .B(n51652), .CI(\intadd_3/n6 ), 
        .CO(\intadd_3/n5 ), .S(\intadd_2/B[6] ) );
  FA_X1 \intadd_3/U5  ( .A(\intadd_3/A[9] ), .B(n51649), .CI(\intadd_3/n5 ), 
        .CO(\intadd_3/n4 ), .S(\intadd_2/B[7] ) );
  FA_X1 \intadd_3/U4  ( .A(\intadd_3/A[10] ), .B(n51647), .CI(\intadd_3/n4 ), 
        .CO(\intadd_3/n3 ), .S(\intadd_2/B[8] ) );
  FA_X1 \intadd_3/U3  ( .A(\intadd_3/A[11] ), .B(\intadd_3/B[11] ), .CI(
        \intadd_3/n3 ), .CO(\intadd_3/n2 ), .S(\intadd_2/B[9] ) );
  FA_X1 \intadd_3/U2  ( .A(\intadd_3/A[12] ), .B(\intadd_3/B[12] ), .CI(
        \intadd_3/n2 ), .CO(\intadd_3/n1 ), .S(\intadd_2/B[10] ) );
  FA_X1 \intadd_4/U14  ( .A(\intadd_4/A[0] ), .B(n51691), .CI(\intadd_4/CI ), 
        .CO(\intadd_4/n13 ), .S(\intadd_4/SUM[0] ) );
  FA_X1 \intadd_4/U13  ( .A(n51688), .B(\intadd_4/B[1] ), .CI(\intadd_4/n13 ), 
        .CO(\intadd_4/n12 ), .S(\intadd_4/SUM[1] ) );
  FA_X1 \intadd_4/U12  ( .A(n51685), .B(\intadd_4/B[2] ), .CI(\intadd_4/n12 ), 
        .CO(\intadd_4/n11 ), .S(\intadd_4/SUM[2] ) );
  FA_X1 \intadd_4/U11  ( .A(n51681), .B(\intadd_4/B[3] ), .CI(\intadd_4/n11 ), 
        .CO(\intadd_4/n10 ), .S(\intadd_4/SUM[3] ) );
  FA_X1 \intadd_4/U10  ( .A(n51676), .B(\intadd_4/B[4] ), .CI(\intadd_4/n10 ), 
        .CO(\intadd_4/n9 ), .S(\intadd_4/SUM[4] ) );
  FA_X1 \intadd_4/U9  ( .A(n51672), .B(\intadd_4/B[5] ), .CI(\intadd_4/n9 ), 
        .CO(\intadd_4/n8 ), .S(\intadd_4/SUM[5] ) );
  FA_X1 \intadd_4/U8  ( .A(n51668), .B(\intadd_4/B[6] ), .CI(\intadd_4/n8 ), 
        .CO(\intadd_4/n7 ), .S(\intadd_4/SUM[6] ) );
  FA_X1 \intadd_4/U7  ( .A(n51664), .B(\intadd_4/B[7] ), .CI(\intadd_4/n7 ), 
        .CO(\intadd_4/n6 ), .S(\intadd_4/SUM[7] ) );
  FA_X1 \intadd_4/U6  ( .A(n51660), .B(\intadd_4/B[8] ), .CI(\intadd_4/n6 ), 
        .CO(\intadd_4/n5 ), .S(\intadd_4/SUM[8] ) );
  FA_X1 \intadd_4/U5  ( .A(n51656), .B(\intadd_4/B[9] ), .CI(\intadd_4/n5 ), 
        .CO(\intadd_4/n4 ), .S(\intadd_4/SUM[9] ) );
  FA_X1 \intadd_4/U4  ( .A(n51653), .B(\intadd_4/B[10] ), .CI(\intadd_4/n4 ), 
        .CO(\intadd_4/n3 ), .S(\intadd_4/SUM[10] ) );
  FA_X1 \intadd_4/U3  ( .A(\intadd_4/A[11] ), .B(\intadd_4/B[11] ), .CI(
        \intadd_4/n3 ), .CO(\intadd_4/n2 ), .S(\intadd_4/SUM[11] ) );
  FA_X1 \intadd_4/U2  ( .A(\intadd_4/A[12] ), .B(\intadd_4/B[12] ), .CI(
        \intadd_4/n2 ), .CO(\intadd_4/n1 ), .S(\intadd_4/SUM[12] ) );
  FA_X1 \intadd_5/U14  ( .A(\intadd_5/A[0] ), .B(\intadd_5/B[0] ), .CI(n51696), 
        .CO(\intadd_5/n13 ), .S(\intadd_5/SUM[0] ) );
  FA_X1 \intadd_5/U13  ( .A(\intadd_5/A[1] ), .B(n51694), .CI(\intadd_5/n13 ), 
        .CO(\intadd_5/n12 ), .S(\intadd_5/SUM[1] ) );
  FA_X1 \intadd_5/U12  ( .A(\intadd_5/A[2] ), .B(n51692), .CI(\intadd_5/n12 ), 
        .CO(\intadd_5/n11 ), .S(\intadd_5/SUM[2] ) );
  FA_X1 \intadd_5/U11  ( .A(\intadd_5/A[3] ), .B(n51689), .CI(\intadd_5/n11 ), 
        .CO(\intadd_5/n10 ), .S(\intadd_5/SUM[3] ) );
  FA_X1 \intadd_5/U10  ( .A(\intadd_5/A[4] ), .B(n51686), .CI(\intadd_5/n10 ), 
        .CO(\intadd_5/n9 ), .S(\intadd_5/SUM[4] ) );
  FA_X1 \intadd_5/U9  ( .A(\intadd_5/A[5] ), .B(n51682), .CI(\intadd_5/n9 ), 
        .CO(\intadd_5/n8 ), .S(\intadd_5/SUM[5] ) );
  FA_X1 \intadd_5/U8  ( .A(\intadd_5/A[6] ), .B(n51677), .CI(\intadd_5/n8 ), 
        .CO(\intadd_5/n7 ), .S(\intadd_5/SUM[6] ) );
  FA_X1 \intadd_5/U7  ( .A(\intadd_5/A[7] ), .B(n51673), .CI(\intadd_5/n7 ), 
        .CO(\intadd_5/n6 ), .S(\intadd_5/SUM[7] ) );
  FA_X1 \intadd_5/U6  ( .A(\intadd_5/A[8] ), .B(n51669), .CI(\intadd_5/n6 ), 
        .CO(\intadd_5/n5 ), .S(\intadd_5/SUM[8] ) );
  FA_X1 \intadd_5/U5  ( .A(\intadd_5/A[9] ), .B(n51665), .CI(\intadd_5/n5 ), 
        .CO(\intadd_5/n4 ), .S(\intadd_5/SUM[9] ) );
  FA_X1 \intadd_5/U4  ( .A(\intadd_5/A[10] ), .B(n51661), .CI(\intadd_5/n4 ), 
        .CO(\intadd_5/n3 ), .S(\intadd_5/SUM[10] ) );
  FA_X1 \intadd_5/U3  ( .A(\intadd_5/A[11] ), .B(n19108), .CI(\intadd_5/n3 ), 
        .CO(\intadd_5/n2 ), .S(\intadd_5/SUM[11] ) );
  FA_X1 \intadd_5/U2  ( .A(\intadd_5/A[12] ), .B(\intadd_5/B[12] ), .CI(
        \intadd_5/n2 ), .CO(\intadd_5/n1 ), .S(\intadd_5/SUM[12] ) );
  FA_X1 \intadd_6/U14  ( .A(\intadd_6/A[0] ), .B(n51699), .CI(\intadd_6/CI ), 
        .CO(\intadd_6/n13 ), .S(\intadd_6/SUM[0] ) );
  FA_X1 \intadd_6/U13  ( .A(n51698), .B(\intadd_6/B[1] ), .CI(\intadd_6/n13 ), 
        .CO(\intadd_6/n12 ), .S(\intadd_6/SUM[1] ) );
  FA_X1 \intadd_6/U12  ( .A(n51697), .B(\intadd_6/B[2] ), .CI(\intadd_6/n12 ), 
        .CO(\intadd_6/n11 ), .S(\intadd_6/SUM[2] ) );
  FA_X1 \intadd_6/U11  ( .A(n51695), .B(\intadd_6/B[3] ), .CI(\intadd_6/n11 ), 
        .CO(\intadd_6/n10 ), .S(\intadd_6/SUM[3] ) );
  FA_X1 \intadd_6/U10  ( .A(n51693), .B(\intadd_6/B[4] ), .CI(\intadd_6/n10 ), 
        .CO(\intadd_6/n9 ), .S(\intadd_6/SUM[4] ) );
  FA_X1 \intadd_6/U9  ( .A(n51690), .B(\intadd_6/B[5] ), .CI(\intadd_6/n9 ), 
        .CO(\intadd_6/n8 ), .S(\intadd_6/SUM[5] ) );
  FA_X1 \intadd_6/U8  ( .A(n51687), .B(\intadd_6/B[6] ), .CI(\intadd_6/n8 ), 
        .CO(\intadd_6/n7 ), .S(\intadd_6/SUM[6] ) );
  FA_X1 \intadd_6/U7  ( .A(n51683), .B(\intadd_6/B[7] ), .CI(\intadd_6/n7 ), 
        .CO(\intadd_6/n6 ), .S(\intadd_6/SUM[7] ) );
  FA_X1 \intadd_6/U6  ( .A(n51678), .B(\intadd_6/B[8] ), .CI(\intadd_6/n6 ), 
        .CO(\intadd_6/n5 ), .S(\intadd_6/SUM[8] ) );
  FA_X1 \intadd_6/U5  ( .A(n51674), .B(\intadd_6/B[9] ), .CI(\intadd_6/n5 ), 
        .CO(\intadd_6/n4 ), .S(\intadd_6/SUM[9] ) );
  FA_X1 \intadd_6/U4  ( .A(n51670), .B(\intadd_6/B[10] ), .CI(\intadd_6/n4 ), 
        .CO(\intadd_6/n3 ), .S(\intadd_6/SUM[10] ) );
  FA_X1 \intadd_6/U3  ( .A(\intadd_6/A[11] ), .B(\intadd_6/B[11] ), .CI(
        \intadd_6/n3 ), .CO(\intadd_6/n2 ), .S(\intadd_6/SUM[11] ) );
  FA_X1 \intadd_6/U2  ( .A(\intadd_6/A[12] ), .B(\intadd_6/B[12] ), .CI(
        \intadd_6/n2 ), .CO(\intadd_6/n1 ), .S(\intadd_6/SUM[12] ) );
  FA_X1 \intadd_7/U14  ( .A(\intadd_7/A[0] ), .B(\intadd_7/B[0] ), .CI(
        \intadd_7/CI ), .CO(\intadd_7/n13 ), .S(\intadd_7/SUM[0] ) );
  FA_X1 \intadd_7/U13  ( .A(\intadd_7/A[1] ), .B(\intadd_7/B[1] ), .CI(
        \intadd_7/n13 ), .CO(\intadd_7/n12 ), .S(\intadd_7/SUM[1] ) );
  FA_X1 \intadd_7/U12  ( .A(\intadd_7/A[2] ), .B(\intadd_7/B[2] ), .CI(
        \intadd_7/n12 ), .CO(\intadd_7/n11 ), .S(\intadd_7/SUM[2] ) );
  FA_X1 \intadd_7/U11  ( .A(\intadd_7/A[3] ), .B(\intadd_7/B[3] ), .CI(
        \intadd_7/n11 ), .CO(\intadd_7/n10 ), .S(\intadd_7/SUM[3] ) );
  FA_X1 \intadd_7/U10  ( .A(\intadd_7/A[4] ), .B(\intadd_7/B[4] ), .CI(
        \intadd_7/n10 ), .CO(\intadd_7/n9 ), .S(\intadd_7/SUM[4] ) );
  FA_X1 \intadd_7/U9  ( .A(\intadd_7/A[5] ), .B(\intadd_7/B[5] ), .CI(
        \intadd_7/n9 ), .CO(\intadd_7/n8 ), .S(\intadd_7/SUM[5] ) );
  FA_X1 \intadd_7/U8  ( .A(\intadd_7/A[6] ), .B(\intadd_7/B[6] ), .CI(
        \intadd_7/n8 ), .CO(\intadd_7/n7 ), .S(\intadd_7/SUM[6] ) );
  FA_X1 \intadd_7/U7  ( .A(\intadd_7/A[7] ), .B(\intadd_7/B[7] ), .CI(
        \intadd_7/n7 ), .CO(\intadd_7/n6 ), .S(\intadd_7/SUM[7] ) );
  FA_X1 \intadd_7/U6  ( .A(\intadd_7/A[8] ), .B(\intadd_7/B[8] ), .CI(
        \intadd_7/n6 ), .CO(\intadd_7/n5 ), .S(\intadd_7/SUM[8] ) );
  FA_X1 \intadd_7/U5  ( .A(\intadd_7/A[9] ), .B(\intadd_7/B[9] ), .CI(
        \intadd_7/n5 ), .CO(\intadd_7/n4 ), .S(\intadd_7/SUM[9] ) );
  FA_X1 \intadd_7/U4  ( .A(\intadd_7/A[10] ), .B(\intadd_7/B[10] ), .CI(
        \intadd_7/n4 ), .CO(\intadd_7/n3 ), .S(\intadd_7/SUM[10] ) );
  FA_X1 \intadd_7/U3  ( .A(\intadd_7/A[11] ), .B(\intadd_7/B[11] ), .CI(
        \intadd_7/n3 ), .CO(\intadd_7/n2 ), .S(\intadd_7/SUM[11] ) );
  FA_X1 \intadd_7/U2  ( .A(\intadd_7/A[12] ), .B(\intadd_7/B[12] ), .CI(
        \intadd_7/n2 ), .CO(\intadd_7/n1 ), .S(\intadd_7/SUM[12] ) );
  DFFR_X1 \CU/cw1_reg[9]  ( .D(n3191), .CK(CLK), .RN(RST), .Q(\CU/cw1[9] ) );
  DFFR_X1 \CU/cw1_reg[15]  ( .D(n3190), .CK(CLK), .RN(RST), .Q(\CU/cw1[15] )
         );
  DFFR_X1 \CU/cw1_reg[19]  ( .D(n9315), .CK(CLK), .RN(RST), .Q(\CU/cw1[19] )
         );
  FA_X1 \intadd_8/U5  ( .A(\intadd_0/n1 ), .B(n51800), .CI(\intadd_8/CI ), 
        .CO(\intadd_8/n4 ), .S(\intadd_8/SUM[0] ) );
  FA_X1 \intadd_8/U4  ( .A(n51801), .B(\intadd_8/B[1] ), .CI(\intadd_8/n4 ), 
        .CO(\intadd_8/n3 ), .S(\intadd_8/SUM[1] ) );
  FA_X1 \intadd_8/U3  ( .A(n51802), .B(\intadd_8/B[2] ), .CI(\intadd_8/n3 ), 
        .CO(\intadd_8/n2 ), .S(\intadd_8/SUM[2] ) );
  FA_X1 \intadd_8/U2  ( .A(n51803), .B(\intadd_8/B[3] ), .CI(\intadd_8/n2 ), 
        .CO(\intadd_8/n1 ), .S(\intadd_8/SUM[3] ) );
  DFF_X1 \DP/RegRD3/DOUT_reg[4]  ( .D(\DP/RegRD3/n10 ), .CK(n4991), .Q(n53515), 
        .QN(n53693) );
  DFF_X1 \DP/RegRD3/DOUT_reg[3]  ( .D(\DP/RegRD3/n11 ), .CK(n4991), .Q(n49866)
         );
  DFF_X1 \DP/RegNPC4/DOUT_reg[30]  ( .D(n5054), .CK(n5088), .QN(n53386) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[28]  ( .D(n5052), .CK(n5088), .QN(n49937) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[26]  ( .D(n5050), .CK(n5088), .Q(n53702), .QN(
        n53387) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[22]  ( .D(n5046), .CK(n5088), .QN(n53379) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[12]  ( .D(n5036), .CK(n5088), .QN(n53383) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[10]  ( .D(n5034), .CK(n5088), .QN(n53368) );
  DFF_X1 \IR/DOUT_reg[10]  ( .D(n5139), .CK(n5185), .Q(n53552), .QN(n53745) );
  DFF_X1 \IR/DOUT_reg[9]  ( .D(n5138), .CK(n5185), .Q(n53551), .QN(n53747) );
  DFF_X1 \IR/DOUT_reg[8]  ( .D(n5137), .CK(n5185), .QN(n49909) );
  DFF_X1 \DP/RegALU3/DOUT_reg[28]  ( .D(\DP/RegALU3/n71 ), .CK(n4991), .Q(
        n49872), .QN(n53665) );
  DFF_X1 \DP/RegALU3/DOUT_reg[15]  ( .D(\DP/RegALU3/n84 ), .CK(n4991), .QN(
        n49809) );
  DFF_X1 \DP/RegALU3/DOUT_reg[9]  ( .D(\DP/RegALU3/n90 ), .CK(n4991), .QN(
        n49832) );
  DFF_X1 \DP/RegALU3/DOUT_reg[6]  ( .D(\DP/RegALU3/n93 ), .CK(n4991), .Q(
        n53757), .QN(n49811) );
  DFF_X1 \DP/RegALU3/DOUT_reg[25]  ( .D(\DP/RegALU3/n74 ), .CK(n4991), .Q(
        n53709), .QN(n49842) );
  DFF_X1 \DP/RegALU3/DOUT_reg[21]  ( .D(\DP/RegALU3/n78 ), .CK(n4991), .Q(
        n7660), .QN(n53668) );
  DFF_X1 \DP/RegALU3/DOUT_reg[0]  ( .D(n4925), .CK(n4991), .Q(DRAM_ADDR[0]), 
        .QN(n3260) );
  DFF_X1 \DP/RegALU3/DOUT_reg[23]  ( .D(\DP/RegALU3/n76 ), .CK(n4991), .Q(
        n7661), .QN(n53669) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[17]  ( .D(n5041), .CK(n5088), .Q(n53377) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[9]  ( .D(n5033), .CK(n5088), .Q(n49958) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[3]  ( .G(n53818), .D(n3083), .Q(
        \DP/ALU0/S_B_MULT[3] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[13]  ( .G(n53818), .D(n3145), .Q(
        \DP/ALU0/S_B_MULT[13] ) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[15]  ( .D(n5039), .CK(n5088), .Q(n53384) );
  DFF_X1 \DP/FU/RS2_EX_reg[1]  ( .D(n18754), .CK(n4923), .QN(n53272) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[7]  ( .G(n53818), .D(n3071), .Q(
        \DP/ALU0/S_B_MULT[7] ) );
  DFF_X1 \PC/DOUT_reg[6]  ( .D(n5119), .CK(n5185), .Q(n53794), .QN(n49907) );
  DFF_X1 \DP/RegRD4/DOUT_reg[0]  ( .D(\DP/RegRD4/n12 ), .CK(n5088), .Q(
        \DP/RD4[0] ), .QN(n26670) );
  DFF_X1 \DP/RegRD4/DOUT_reg[2]  ( .D(\DP/RegRD4/n13 ), .CK(n5088), .Q(
        \DP/RD4[2] ), .QN(n3015) );
  DFF_X1 \DP/RegRD3/DOUT_reg[2]  ( .D(\DP/RegRD3/n12 ), .CK(n4991), .Q(n53753), 
        .QN(n7617) );
  DFF_X1 \DP/RegRD3/DOUT_reg[1]  ( .D(\DP/RegRD3/n13 ), .CK(n4991), .Q(n49819)
         );
  DFF_X1 \DP/RegRD3/DOUT_reg[0]  ( .D(\DP/RegRD3/n14 ), .CK(n4991), .Q(n49857), 
        .QN(n53673) );
  DFF_X1 \DP/RegRD4/DOUT_reg[4]  ( .D(\DP/RegRD4/n14 ), .CK(n5088), .Q(
        \DP/RD4[4] ) );
  DFF_X1 \DP/RegRD4/DOUT_reg[3]  ( .D(\DP/RegRD4/n10 ), .CK(n5088), .Q(
        \DP/RD4[3] ), .QN(n49659) );
  DFF_X1 \DP/RegLMD/DOUT_reg[7]  ( .D(n4999), .CK(n5088), .Q(n49869) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[2]  ( .D(n5026), .CK(n5088), .QN(n49938) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[29]  ( .D(n5053), .CK(n5088), .Q(n53373), .QN(
        n53787) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[24]  ( .D(n5048), .CK(n5088), .QN(n49942) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[18]  ( .D(n5042), .CK(n5088), .Q(n53781), .QN(
        n53382) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[16]  ( .D(n5040), .CK(n5088), .Q(n53797), .QN(
        n49951) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[14]  ( .D(n5038), .CK(n5088), .QN(n53385) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[11]  ( .D(n5035), .CK(n5088), .Q(n53369), .QN(
        n53801) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[8]  ( .D(n5032), .CK(n5088), .Q(n53798), .QN(
        n53370) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[4]  ( .D(n5028), .CK(n5088), .Q(n53743), .QN(
        n49940) );
  DFF_X1 \IR/DOUT_reg[29]  ( .D(n5121), .CK(n5185), .Q(w_IR_OUT[29]), .QN(
        n53681) );
  DFF_X1 \IR/DOUT_reg[28]  ( .D(n5125), .CK(n5185), .Q(w_IR_OUT[28]), .QN(
        n53651) );
  DFF_X1 \IR/DOUT_reg[27]  ( .D(n5151), .CK(n5185), .Q(w_IR_OUT[27]), .QN(
        n53682) );
  DFF_X1 \IR/DOUT_reg[26]  ( .D(n5150), .CK(n5185), .Q(w_IR_OUT[26]), .QN(
        n53678) );
  DFF_X1 \IR/DOUT_reg[25]  ( .D(n5122), .CK(n5185), .Q(\DP/IMMS26[25] ), .QN(
        \IR/n61 ) );
  DFF_X1 \IR/DOUT_reg[24]  ( .D(n5127), .CK(n5185), .Q(\DP/IMMS26[24] ), .QN(
        \IR/n60 ) );
  DFF_X1 \IR/DOUT_reg[23]  ( .D(n5124), .CK(n5185), .Q(\DP/IMMS26[23] ), .QN(
        \IR/n59 ) );
  DFF_X1 \IR/DOUT_reg[22]  ( .D(n5126), .CK(n5185), .Q(\DP/IMMS26[22] ), .QN(
        \IR/n58 ) );
  DFF_X1 \IR/DOUT_reg[21]  ( .D(n5128), .CK(n5185), .Q(\DP/IMMS26[21] ), .QN(
        \IR/n57 ) );
  DFF_X1 \IR/DOUT_reg[20]  ( .D(n5149), .CK(n5185), .Q(n53561), .QN(n53699) );
  DFF_X1 \IR/DOUT_reg[19]  ( .D(n5148), .CK(n5185), .Q(n53560), .QN(n53698) );
  DFF_X1 \IR/DOUT_reg[18]  ( .D(n5147), .CK(n5185), .Q(n53559), .QN(n53697) );
  DFF_X1 \IR/DOUT_reg[17]  ( .D(n5146), .CK(n5185), .Q(n53558), .QN(n53696) );
  DFF_X1 \IR/DOUT_reg[16]  ( .D(n5145), .CK(n5185), .Q(n53557), .QN(n53695) );
  DFF_X1 \IR/DOUT_reg[15]  ( .D(n5144), .CK(n5185), .Q(n53704), .QN(n7667) );
  DFF_X1 \IR/DOUT_reg[14]  ( .D(n5143), .CK(n5185), .Q(n53556), .QN(n53751) );
  DFF_X1 \IR/DOUT_reg[13]  ( .D(n5142), .CK(n5185), .Q(n53555), .QN(n53750) );
  DFF_X1 \IR/DOUT_reg[12]  ( .D(n5141), .CK(n5185), .Q(n53554), .QN(n53749) );
  DFF_X1 \IR/DOUT_reg[11]  ( .D(n5140), .CK(n5185), .Q(n53553), .QN(n53748) );
  DFF_X1 \IR/DOUT_reg[7]  ( .D(n5136), .CK(n5185), .QN(n49908) );
  DFF_X1 \IR/DOUT_reg[6]  ( .D(n5135), .CK(n5185), .Q(n53550), .QN(n53746) );
  DFF_X1 \IR/DOUT_reg[5]  ( .D(n5134), .CK(n5185), .Q(n49853), .QN(n53687) );
  DFF_X1 \IR/DOUT_reg[4]  ( .D(n5133), .CK(n5185), .Q(n53688), .QN(n7616) );
  DFF_X1 \IR/DOUT_reg[3]  ( .D(n5132), .CK(n5185), .Q(n53549), .QN(n53649) );
  DFF_X1 \IR/DOUT_reg[2]  ( .D(n5131), .CK(n5185), .Q(n53689), .QN(n7564) );
  DFF_X1 \IR/DOUT_reg[1]  ( .D(n5130), .CK(n5185), .Q(n53548), .QN(n53686) );
  DFF_X1 \IR/DOUT_reg[0]  ( .D(n5129), .CK(n5185), .Q(n53652), .QN(n49849) );
  DFF_X1 \DP/RegALU3/DOUT_reg[30]  ( .D(\DP/RegALU3/n69 ), .CK(n4991), .Q(
        n53710), .QN(n49834) );
  DFF_X1 \DP/RegALU3/DOUT_reg[3]  ( .D(\DP/RegALU3/n96 ), .CK(n4991), .Q(
        DRAM_ADDR[3]), .QN(n3254) );
  DFF_X1 \DP/RegALU3/DOUT_reg[12]  ( .D(\DP/RegALU3/n87 ), .CK(n4991), .Q(
        n53755), .QN(n49814) );
  DFF_X1 \DP/RegALU3/DOUT_reg[4]  ( .D(n9277), .CK(n4991), .Q(DRAM_ADDR[4]), 
        .QN(n3248) );
  DFF_X1 \DP/RegALU3/DOUT_reg[1]  ( .D(n4926), .CK(n4991), .Q(DRAM_ADDR[1]), 
        .QN(n3273) );
  DFF_X1 \DP/RegALU3/DOUT_reg[7]  ( .D(\DP/RegALU3/n92 ), .CK(n4991), .Q(n7620), .QN(n53662) );
  DFF_X1 \DP/RegALU3/DOUT_reg[29]  ( .D(\DP/RegALU3/n70 ), .CK(n4991), .Q(
        n7625), .QN(n53663) );
  DFF_X1 \DP/RegALU3/DOUT_reg[14]  ( .D(\DP/RegALU3/n85 ), .CK(n4991), .Q(
        n7624), .QN(n53660) );
  DFF_X1 \DP/RegALU3/DOUT_reg[8]  ( .D(\DP/RegALU3/n91 ), .CK(n4991), .Q(n7676), .QN(n53661) );
  DFF_X1 \DP/RegALU3/DOUT_reg[5]  ( .D(\DP/RegALU3/n94 ), .CK(n4991), .Q(
        DRAM_ADDR[5]), .QN(n3249) );
  DFF_X1 \DP/RegALU3/DOUT_reg[2]  ( .D(\DP/RegALU3/n97 ), .CK(n4991), .Q(
        DRAM_ADDR[2]), .QN(n3247) );
  DFF_X1 \DP/RegALU3/DOUT_reg[31]  ( .D(\DP/RegALU3/n68 ), .CK(n4991), .Q(
        n7626), .QN(n53664) );
  DFF_X1 \DP/RegALU3/DOUT_reg[26]  ( .D(\DP/RegALU3/n73 ), .CK(n4991), .Q(
        n53648), .QN(n49838) );
  DFF_X1 \DP/RegALU3/DOUT_reg[24]  ( .D(\DP/RegALU3/n75 ), .CK(n4991), .Q(
        n53706), .QN(n49839) );
  DFF_X1 \DP/RegALU3/DOUT_reg[22]  ( .D(\DP/RegALU3/n77 ), .CK(n4991), .Q(
        n7622), .QN(n53670) );
  DFF_X1 \DP/RegALU3/DOUT_reg[20]  ( .D(\DP/RegALU3/n79 ), .CK(n4991), .Q(
        n7621), .QN(n53667) );
  DFF_X1 \DP/RegALU3/DOUT_reg[18]  ( .D(\DP/RegALU3/n81 ), .CK(n4991), .Q(
        n7663), .QN(n53666) );
  DFF_X1 \DP/RegALU3/DOUT_reg[16]  ( .D(\DP/RegALU3/n83 ), .CK(n4991), .Q(
        n7662), .QN(n53671) );
  DFF_X1 \DP/RegNPC4/DOUT_reg[27]  ( .D(n5051), .CK(n5088), .Q(n53375) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[9]  ( .G(n53818), .D(n3065), .Q(
        \DP/ALU0/S_B_MULT[9] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[1]  ( .G(n53818), .D(n3089), .Q(
        \DP/ALU0/S_B_MULT[1] ) );
  DFF_X1 \IR/DOUT_reg[30]  ( .D(n5152), .CK(n5185), .Q(w_IR_OUT[30]), .QN(
        n53683) );
  DFF_X1 \DP/FU/RS2_EX_reg[3]  ( .D(n7286), .CK(n4923), .Q(n53271) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[5]  ( .G(n53818), .D(n3077), .Q(
        \DP/ALU0/S_B_MULT[5] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[31]  ( .D(n5153), .CK(n5185), .Q(n53593) );
  DFF_X1 \PC/DOUT_reg[9]  ( .D(n5096), .CK(n5185), .Q(w_PC_OUT[9]), .QN(n53779) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[15]  ( .G(\DP/ALU0/n109 ), .D(n3140), .Q(
        \DP/ALU0/s_A_MULT[15] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[1]  ( .G(n53818), .D(n3088), .Q(
        \DP/ALU0/s_A_MULT[1] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[11]  ( .G(n53818), .D(n3059), .Q(
        \DP/ALU0/S_B_MULT[11] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[12]  ( .G(n53818), .D(n3146), .Q(
        \DP/ALU0/s_A_MULT[12] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[3]  ( .G(\DP/ALU0/n109 ), .D(n3082), .Q(
        \DP/ALU0/s_A_MULT[3] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[9]  ( .G(\DP/ALU0/n109 ), .D(n3064), .Q(
        \DP/ALU0/s_A_MULT[9] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[2]  ( .G(\DP/ALU0/n109 ), .D(n3085), .Q(
        \DP/ALU0/s_A_MULT[2] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[10]  ( .G(\DP/ALU0/n109 ), .D(n3061), .Q(
        \DP/ALU0/s_A_MULT[10] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[7]  ( .G(\DP/ALU0/n109 ), .D(n3070), .Q(
        \DP/ALU0/s_A_MULT[7] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[5]  ( .G(\DP/ALU0/n109 ), .D(n3076), .Q(
        \DP/ALU0/s_A_MULT[5] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[11]  ( .G(\DP/ALU0/n109 ), .D(n3058), .Q(
        \DP/ALU0/s_A_MULT[11] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[4]  ( .G(\DP/ALU0/n109 ), .D(n3079), .Q(
        \DP/ALU0/s_A_MULT[4] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[6]  ( .G(\DP/ALU0/n109 ), .D(n3073), .Q(
        \DP/ALU0/s_A_MULT[6] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[8]  ( .G(\DP/ALU0/n109 ), .D(n3067), .Q(
        \DP/ALU0/s_A_MULT[8] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[13]  ( .G(\DP/ALU0/n109 ), .D(n3144), .Q(
        \DP/ALU0/s_A_MULT[13] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[14]  ( .G(\DP/ALU0/n109 ), .D(n3142), .Q(
        \DP/ALU0/s_A_MULT[14] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[0]  ( .G(\DP/ALU0/n109 ), .D(n3091), .Q(
        \DP/ALU0/s_A_MULT[0] ) );
  DFF_X1 \DP/RegRD4/DOUT_reg[1]  ( .D(\DP/RegRD4/n11 ), .CK(n5088), .Q(
        \DP/RD4[1] ) );
  DFFR_X2 \CU/cw5_reg[0]  ( .D(\CU/cw4[0] ), .CK(CLK), .RN(RST), .Q(n53705), 
        .QN(n53650) );
  DFFR_X2 \CU/cw5_reg[2]  ( .D(\CU/cw4[2] ), .CK(CLK), .RN(RST), .Q(n53647), 
        .QN(n53684) );
  DFF_X1 \DP/FU/RS2_EX_reg[4]  ( .D(n53261), .CK(n4923), .Q(n53274) );
  OAI33_X1 U35941 ( .A1(1'b0), .A2(n53854), .A3(n53635), .B1(n49849), .B2(
        n53862), .B3(n7564), .ZN(n53637) );
  OAI33_X1 U35942 ( .A1(1'b0), .A2(n53627), .A3(n53628), .B1(
        \DP/ALU0/S_B_MULT[13] ), .B2(n54858), .B3(n54056), .ZN(n53630) );
  NOR4_X1 U35943 ( .A1(n55330), .A2(n53552), .A3(n53550), .A4(n53551), .ZN(
        n53614) );
  NAND3_X1 U35944 ( .A1(n53614), .A2(n49908), .A3(n49909), .ZN(n53826) );
  INV_X1 U35945 ( .A(n54858), .ZN(n53615) );
  OAI21_X1 U35946 ( .B1(\DP/ALU0/S_B_MULT[7] ), .B2(\DP/ALU0/S_B_MULT[8] ), 
        .A(n53615), .ZN(n53616) );
  NAND3_X1 U35947 ( .A1(\DP/ALU0/S_B_MULT[9] ), .A2(n54037), .A3(n54055), .ZN(
        n53617) );
  OAI21_X1 U35948 ( .B1(\DP/ALU0/S_B_MULT[9] ), .B2(n53616), .A(n53617), .ZN(
        n53618) );
  INV_X1 U35949 ( .A(n54741), .ZN(n53619) );
  INV_X1 U35950 ( .A(\intadd_4/n1 ), .ZN(n53620) );
  OAI221_X1 U35951 ( .B1(n54741), .B2(n54740), .C1(n53619), .C2(n53620), .A(
        n54738), .ZN(n53621) );
  XOR2_X1 U35952 ( .A(n53618), .B(n53621), .Z(n54697) );
  AOI21_X1 U35953 ( .B1(n53678), .B2(n53871), .A(n53870), .ZN(n53622) );
  NAND4_X1 U35954 ( .A1(n53872), .A2(n53867), .A3(n53868), .A4(n53622), .ZN(
        \CU/cw[17] ) );
  NAND2_X1 U35955 ( .A1(n49955), .A2(n53798), .ZN(n53623) );
  NOR3_X1 U35956 ( .A1(n55333), .A2(n53414), .A3(n53623), .ZN(n54932) );
  INV_X1 U35957 ( .A(n54613), .ZN(n53624) );
  INV_X1 U35958 ( .A(n54611), .ZN(n53625) );
  AOI221_X1 U35959 ( .B1(n54608), .B2(n53624), .C1(\intadd_2/n1 ), .C2(n54613), 
        .A(n53625), .ZN(n53626) );
  NAND2_X1 U35960 ( .A1(n54055), .A2(n54054), .ZN(n53627) );
  INV_X1 U35961 ( .A(\DP/ALU0/S_B_MULT[13] ), .ZN(n53628) );
  XOR2_X1 U35963 ( .A(n53626), .B(n53630), .Z(n54111) );
  AND3_X1 U35964 ( .A1(w_PC_OUT[13]), .A2(n53594), .A3(n55317), .ZN(n55347) );
  AOI21_X1 U35965 ( .B1(n53891), .B2(n53863), .A(w_IR_OUT[26]), .ZN(n53631) );
  NAND2_X1 U35966 ( .A1(n53678), .A2(n53853), .ZN(n53632) );
  AOI21_X1 U35967 ( .B1(n53632), .B2(n53870), .A(n53631), .ZN(n53633) );
  INV_X1 U35968 ( .A(n53879), .ZN(n53634) );
  INV_X1 U35969 ( .A(n49849), .ZN(n53635) );
  AOI211_X1 U35971 ( .C1(n53852), .C2(n53634), .A(n53859), .B(n53637), .ZN(
        n53638) );
  OAI211_X1 U35972 ( .C1(n53853), .C2(n53883), .A(n53633), .B(n53638), .ZN(
        \CU/aluOpcodei[2] ) );
  INV_X4 U35973 ( .A(n53774), .ZN(n53611) );
  AND2_X1 U35974 ( .A1(n54530), .A2(n54548), .ZN(n54547) );
  AND2_X1 U35975 ( .A1(n55359), .A2(n53777), .ZN(n55288) );
  OR2_X1 U35976 ( .A1(n55353), .A2(n53791), .ZN(n55358) );
  OR2_X1 U35977 ( .A1(n54974), .A2(n53768), .ZN(n53694) );
  OR3_X1 U35978 ( .A1(n54974), .A2(n53768), .A3(n53786), .ZN(n53685) );
  NAND2_X1 U35979 ( .A1(n54941), .A2(n53374), .ZN(n54974) );
  INV_X1 U35980 ( .A(n55312), .ZN(n55181) );
  INV_X2 U35981 ( .A(n54411), .ZN(n55175) );
  INV_X1 U35982 ( .A(n55186), .ZN(n55306) );
  INV_X2 U35983 ( .A(n55177), .ZN(n55137) );
  NAND2_X2 U35984 ( .A1(n53814), .A2(n55282), .ZN(n55284) );
  OR2_X2 U35985 ( .A1(n53815), .A2(n55282), .ZN(n55283) );
  OR2_X1 U35986 ( .A1(n54952), .A2(n53788), .ZN(n54947) );
  OR3_X1 U35987 ( .A1(\DP/ALU0/S_B_MULT[7] ), .A2(\DP/ALU0/S_B_MULT[8] ), .A3(
        n54038), .ZN(n54776) );
  OR3_X1 U35988 ( .A1(\DP/ALU0/S_B_MULT[5] ), .A2(\DP/ALU0/S_B_MULT[6] ), .A3(
        n54034), .ZN(n54810) );
  OR3_X1 U35989 ( .A1(\DP/ALU0/S_B_MULT[1] ), .A2(\DP/ALU0/S_B_MULT[2] ), .A3(
        n54020), .ZN(n54921) );
  OR3_X1 U35990 ( .A1(\DP/ALU0/S_B_MULT[3] ), .A2(\DP/ALU0/S_B_MULT[4] ), .A3(
        n54005), .ZN(n54846) );
  OR3_X1 U35991 ( .A1(\DP/ALU0/S_B_MULT[13] ), .A2(\DP/ALU0/S_B_MULT[14] ), 
        .A3(n53986), .ZN(n54660) );
  OR3_X1 U35992 ( .A1(\DP/ALU0/S_B_MULT[11] ), .A2(\DP/ALU0/S_B_MULT[12] ), 
        .A3(n54057), .ZN(n54694) );
  AOI21_X1 U35993 ( .B1(w_EQ_COND), .B2(n55281), .A(n55280), .ZN(n55282) );
  NAND2_X1 U35994 ( .A1(n54953), .A2(n53380), .ZN(n54952) );
  OR2_X1 U35995 ( .A1(n54970), .A2(n53775), .ZN(n54955) );
  NAND2_X1 U35996 ( .A1(n54967), .A2(n49952), .ZN(n54970) );
  OR2_X1 U35997 ( .A1(n53783), .A2(n53784), .ZN(n55344) );
  OR2_X1 U35998 ( .A1(n55338), .A2(n53778), .ZN(n53783) );
  OR2_X1 U35999 ( .A1(n53799), .A2(n53800), .ZN(n54963) );
  NAND2_X2 U36000 ( .A1(n53937), .A2(n53763), .ZN(n55120) );
  AND2_X2 U36001 ( .A1(w_MuxA_SEL), .A2(n53937), .ZN(n55118) );
  NAND2_X2 U36002 ( .A1(n53923), .A2(n53762), .ZN(n55106) );
  NAND2_X2 U36003 ( .A1(w_MuxB_SEL), .A2(n53923), .ZN(n55126) );
  AND2_X1 U36004 ( .A1(n55330), .A2(n55329), .ZN(n55331) );
  AND2_X1 U36005 ( .A1(n53794), .A2(n55295), .ZN(n55339) );
  NOR2_X2 U36006 ( .A1(n53920), .A2(n54598), .ZN(n54548) );
  NAND2_X1 U36007 ( .A1(n55134), .A2(n53372), .ZN(n55333) );
  NAND2_X1 U36008 ( .A1(n53919), .A2(n53647), .ZN(n54598) );
  NOR2_X1 U36009 ( .A1(w_IR_OUT[27]), .A2(w_IR_OUT[30]), .ZN(n53853) );
  OR2_X2 U36010 ( .A1(n53974), .A2(n51572), .ZN(\DP/ALU0/N20 ) );
  BUF_X1 U36011 ( .A(n53613), .Z(n53816) );
  NAND2_X2 U36012 ( .A1(n53810), .A2(n53974), .ZN(n55303) );
  BUF_X1 U36013 ( .A(n55198), .Z(n53810) );
  AOI21_X2 U36014 ( .B1(\DP/ALU0/s_A_MULT[13] ), .B2(n54620), .A(n53989), .ZN(
        n54856) );
  AOI21_X2 U36015 ( .B1(\DP/ALU0/s_A_MULT[11] ), .B2(n54615), .A(n54622), .ZN(
        n54870) );
  AOI21_X2 U36016 ( .B1(\DP/ALU0/s_A_MULT[4] ), .B2(n54634), .A(n54633), .ZN(
        n54890) );
  AOI21_X2 U36017 ( .B1(\DP/ALU0/s_A_MULT[5] ), .B2(n54638), .A(n54637), .ZN(
        n54894) );
  AOI21_X2 U36018 ( .B1(\DP/ALU0/s_A_MULT[6] ), .B2(n54642), .A(n54641), .ZN(
        n54898) );
  AOI21_X2 U36019 ( .B1(\DP/ALU0/s_A_MULT[7] ), .B2(n54646), .A(n54645), .ZN(
        n54902) );
  AOI21_X2 U36020 ( .B1(\DP/ALU0/s_A_MULT[8] ), .B2(n54650), .A(n54649), .ZN(
        n54906) );
  AOI21_X2 U36021 ( .B1(\DP/ALU0/s_A_MULT[9] ), .B2(n54654), .A(n54653), .ZN(
        n54914) );
  AOI21_X2 U36022 ( .B1(\DP/ALU0/s_A_MULT[10] ), .B2(n54617), .A(n54616), .ZN(
        n54869) );
  AOI21_X2 U36023 ( .B1(n54470), .B2(\DP/ALU0/s_A_MULT[2] ), .A(n54630), .ZN(
        n54885) );
  NOR3_X2 U36024 ( .A1(w_IR_OUT[28]), .A2(n53886), .A3(n53890), .ZN(n45959) );
  INV_X1 U36025 ( .A(n54846), .ZN(n53639) );
  INV_X1 U36026 ( .A(n54776), .ZN(n53640) );
  INV_X1 U36027 ( .A(n54810), .ZN(n53641) );
  INV_X1 U36028 ( .A(n54660), .ZN(n53642) );
  INV_X1 U36029 ( .A(n54921), .ZN(n53643) );
  INV_X1 U36030 ( .A(n54694), .ZN(n53644) );
  NOR3_X2 U36031 ( .A1(w_MuxSW_SEL[0]), .A2(w_MuxSW_SEL[1]), .A3(n53677), .ZN(
        n54582) );
  NOR2_X2 U36032 ( .A1(n3021), .A2(n53822), .ZN(n55199) );
  AOI211_X2 U36033 ( .C1(n26670), .C2(n54499), .A(n54498), .B(n54497), .ZN(
        n54537) );
  NOR2_X2 U36034 ( .A1(\DP/ALU0/S_B_MULT[5] ), .A2(n55298), .ZN(n54851) );
  NOR2_X2 U36035 ( .A1(n54005), .A2(n55298), .ZN(n54850) );
  NOR2_X2 U36036 ( .A1(n54039), .A2(n54040), .ZN(n54733) );
  NOR2_X2 U36037 ( .A1(\DP/ALU0/S_B_MULT[9] ), .A2(n54037), .ZN(n54775) );
  NOR2_X2 U36038 ( .A1(\DP/ALU0/S_B_MULT[11] ), .A2(n54041), .ZN(n54732) );
  NOR2_X2 U36039 ( .A1(\DP/ALU0/S_B_MULT[15] ), .A2(n53985), .ZN(n54659) );
  INV_X1 U36040 ( .A(n55103), .ZN(n53645) );
  NOR4_X1 U36041 ( .A1(n53918), .A2(n53912), .A3(n53911), .A4(n53910), .ZN(
        n55121) );
  NOR2_X2 U36042 ( .A1(\DP/ALU0/S_B_MULT[0] ), .A2(n54854), .ZN(n54864) );
  NOR3_X2 U36043 ( .A1(w_MuxSW_SEL[0]), .A2(w_MuxSW_SEL[2]), .A3(n53752), .ZN(
        n54602) );
  NOR4_X4 U36044 ( .A1(n53936), .A2(n53930), .A3(n53929), .A4(n53928), .ZN(
        n55099) );
  NOR2_X2 U36045 ( .A1(n54299), .A2(n54298), .ZN(n55176) );
  NOR2_X2 U36046 ( .A1(\DP/ALU0/S_B_MULT[5] ), .A2(n54025), .ZN(n54849) );
  NOR2_X2 U36047 ( .A1(\DP/ALU0/S_B_MULT[13] ), .A2(n54054), .ZN(n54693) );
  NOR2_X2 U36048 ( .A1(\DP/ALU0/S_B_MULT[3] ), .A2(n54018), .ZN(n54920) );
  NOR2_X2 U36049 ( .A1(\DP/ALU0/S_B_MULT[7] ), .A2(n54032), .ZN(n54809) );
  NOR2_X2 U36050 ( .A1(\DP/ALU0/S_B_MULT[15] ), .A2(n54312), .ZN(n54661) );
  NOR2_X2 U36051 ( .A1(\DP/ALU0/S_B_MULT[11] ), .A2(n54380), .ZN(n54728) );
  NOR2_X2 U36052 ( .A1(\DP/ALU0/S_B_MULT[9] ), .A2(n54403), .ZN(n54777) );
  INV_X1 U36053 ( .A(n55300), .ZN(n55166) );
  BUF_X1 U36054 ( .A(\DP/ALU0/n109 ), .Z(n53818) );
  OR2_X1 U36055 ( .A1(n53900), .A2(n53890), .ZN(n55329) );
  NAND4_X1 U36056 ( .A1(n53825), .A2(n53853), .A3(n53651), .A4(n53678), .ZN(
        n55330) );
  NOR2_X1 U36057 ( .A1(n55350), .A2(n53690), .ZN(n55349) );
  OR2_X1 U36058 ( .A1(n53688), .A2(n53826), .ZN(n53881) );
  NOR2_X1 U36059 ( .A1(n55331), .A2(n53699), .ZN(w_RS2[4]) );
  NOR2_X1 U36060 ( .A1(n55331), .A2(n53698), .ZN(w_RS2[3]) );
  NOR2_X1 U36061 ( .A1(n55331), .A2(n53695), .ZN(w_RS2[0]) );
  INV_X1 U36062 ( .A(n53886), .ZN(n53825) );
  INV_X1 U36063 ( .A(n55354), .ZN(n53815) );
  NOR2_X1 U36064 ( .A1(n55321), .A2(n53658), .ZN(n55355) );
  NOR2_X1 U36065 ( .A1(n55352), .A2(n53691), .ZN(n55351) );
  NOR3_X1 U36066 ( .A1(n3270), .A2(n7228), .A3(n7229), .ZN(n55286) );
  INV_X2 U36067 ( .A(n55187), .ZN(n53809) );
  OAI21_X1 U36068 ( .B1(n55316), .B2(n53680), .A(n53947), .ZN(n53613) );
  INV_X1 U36069 ( .A(n53815), .ZN(n53814) );
  NOR2_X1 U36070 ( .A1(n55331), .A2(n53697), .ZN(w_RS2[2]) );
  AND2_X1 U36071 ( .A1(n53781), .A2(n53782), .ZN(n53780) );
  AND2_X1 U36072 ( .A1(n53377), .A2(n53796), .ZN(n53782) );
  AND2_X1 U36073 ( .A1(n53797), .A2(n53384), .ZN(n53796) );
  AND3_X1 U36074 ( .A1(n54506), .A2(w_SIGN_LD_EN), .A3(n53315), .ZN(n53920) );
  INV_X1 U36075 ( .A(n53815), .ZN(n53813) );
  INV_X1 U36076 ( .A(n53812), .ZN(n53811) );
  AND2_X1 U36077 ( .A1(n53810), .A2(\DP/ALU0/n112 ), .ZN(n54288) );
  NOR2_X1 U36078 ( .A1(n53946), .A2(n53945), .ZN(\DP/ALU0/n109 ) );
  NOR2_X1 U36079 ( .A1(n3020), .A2(n53822), .ZN(n55198) );
  NOR2_X1 U36080 ( .A1(n55331), .A2(n53696), .ZN(w_RS2[1]) );
  OR2_X1 U36081 ( .A1(n53703), .A2(n53385), .ZN(n53775) );
  NOR3_X1 U36082 ( .A1(w_RF_WE4), .A2(w_MuxLD_SEL[0]), .A3(n53701), .ZN(n54506) );
  NAND2_X1 U36083 ( .A1(n55347), .A2(w_PC_OUT[15]), .ZN(n55350) );
  NAND2_X1 U36084 ( .A1(n55339), .A2(w_PC_OUT[7]), .ZN(n55338) );
  INV_X2 U36085 ( .A(n55199), .ZN(n55200) );
  INV_X1 U36086 ( .A(n55289), .ZN(n55293) );
  INV_X1 U36087 ( .A(n55294), .ZN(n53812) );
  NOR2_X1 U36088 ( .A1(n3019), .A2(n53822), .ZN(n55294) );
  INV_X1 U36089 ( .A(n5463), .ZN(n54286) );
  NAND2_X1 U36090 ( .A1(n53810), .A2(n53818), .ZN(n55300) );
  NAND3_X1 U36091 ( .A1(n53810), .A2(n53949), .A3(n53816), .ZN(n55312) );
  NAND3_X1 U36092 ( .A1(n53816), .A2(n53967), .A3(n53810), .ZN(n55186) );
  OR2_X1 U36093 ( .A1(n53801), .A2(n53368), .ZN(n53800) );
  AND2_X1 U36094 ( .A1(n55252), .A2(n55251), .ZN(n55276) );
  NAND2_X1 U36095 ( .A1(w_IR_OUT[27]), .A2(w_IR_OUT[26]), .ZN(n53890) );
  NOR3_X2 U36096 ( .A1(n49940), .A2(n49938), .A3(n49939), .ZN(n55134) );
  NOR2_X1 U36097 ( .A1(n3018), .A2(n53821), .ZN(n55354) );
  AND2_X1 U36098 ( .A1(RST), .A2(DRAM_DATA_IN[31]), .ZN(n5023) );
  AND2_X1 U36099 ( .A1(RST), .A2(DRAM_DATA_IN[30]), .ZN(n5022) );
  AND2_X1 U36100 ( .A1(RST), .A2(DRAM_DATA_IN[29]), .ZN(n5021) );
  AND2_X1 U36101 ( .A1(RST), .A2(DRAM_DATA_IN[28]), .ZN(n5020) );
  AND2_X1 U36102 ( .A1(RST), .A2(DRAM_DATA_IN[27]), .ZN(n5019) );
  AND2_X1 U36103 ( .A1(RST), .A2(DRAM_DATA_IN[26]), .ZN(n5018) );
  AND2_X1 U36104 ( .A1(RST), .A2(DRAM_DATA_IN[25]), .ZN(n5017) );
  AND2_X1 U36105 ( .A1(RST), .A2(DRAM_DATA_IN[24]), .ZN(n5016) );
  AND2_X1 U36106 ( .A1(RST), .A2(DRAM_DATA_IN[23]), .ZN(n5015) );
  AND2_X1 U36107 ( .A1(RST), .A2(IRAM_DATA[31]), .ZN(n5123) );
  AND2_X1 U36108 ( .A1(RST), .A2(DRAM_DATA_IN[22]), .ZN(n5014) );
  AND2_X1 U36109 ( .A1(RST), .A2(DRAM_DATA_IN[21]), .ZN(n5013) );
  AND2_X1 U36110 ( .A1(RST), .A2(DRAM_DATA_IN[20]), .ZN(n5012) );
  AND2_X1 U36111 ( .A1(RST), .A2(DRAM_DATA_IN[19]), .ZN(n5011) );
  AND2_X1 U36112 ( .A1(RST), .A2(DRAM_DATA_IN[18]), .ZN(n5010) );
  AND2_X1 U36113 ( .A1(RST), .A2(DRAM_DATA_IN[17]), .ZN(n5009) );
  AND2_X1 U36114 ( .A1(RST), .A2(DRAM_DATA_IN[16]), .ZN(n5008) );
  OR2_X1 U36115 ( .A1(n53262), .A2(n55106), .ZN(n55124) );
  INV_X1 U36116 ( .A(n55077), .ZN(n55122) );
  INV_X1 U36117 ( .A(n55121), .ZN(n55103) );
  INV_X1 U36118 ( .A(n55115), .ZN(n55100) );
  NAND2_X1 U36119 ( .A1(n53938), .A2(n55116), .ZN(n55115) );
  INV_X1 U36120 ( .A(n55099), .ZN(n55116) );
  OR2_X1 U36121 ( .A1(n54536), .A2(n54566), .ZN(n54606) );
  AND2_X1 U36122 ( .A1(n54536), .A2(n54602), .ZN(n54593) );
  INV_X1 U36123 ( .A(n53806), .ZN(n53805) );
  NOR2_X1 U36124 ( .A1(n54537), .A2(n54566), .ZN(n54603) );
  NAND3_X1 U36125 ( .A1(n53752), .A2(n53677), .A3(w_MuxSW_SEL[0]), .ZN(n54566)
         );
  INV_X1 U36126 ( .A(n54537), .ZN(n54536) );
  INV_X1 U36127 ( .A(RST), .ZN(n53819) );
  INV_X1 U36128 ( .A(RST), .ZN(n53820) );
  INV_X1 U36129 ( .A(RST), .ZN(n53822) );
  BUF_X1 U36130 ( .A(\DP/ALU0/s_ADD_SUB ), .Z(n53817) );
  INV_X1 U36131 ( .A(RST), .ZN(n53821) );
  INV_X1 U36132 ( .A(n55179), .ZN(n55139) );
  INV_X1 U36133 ( .A(n53760), .ZN(n53807) );
  OR2_X1 U36134 ( .A1(n53956), .A2(n53958), .ZN(n53760) );
  INV_X1 U36135 ( .A(n53761), .ZN(n53804) );
  OR2_X1 U36136 ( .A1(n53958), .A2(n53957), .ZN(n53761) );
  BUF_X1 U36137 ( .A(n55174), .Z(n53808) );
  NOR2_X1 U36138 ( .A1(\DP/ALU0/s_SHIFT[1] ), .A2(\DP/ALU0/s_SHIFT[0] ), .ZN(
        n53955) );
  NOR2_X2 U36139 ( .A1(n49942), .A2(n54947), .ZN(n54941) );
  NOR2_X2 U36140 ( .A1(n53376), .A2(n54955), .ZN(n54953) );
  NOR2_X2 U36141 ( .A1(n53383), .A2(n54963), .ZN(n54967) );
  NOR2_X2 U36142 ( .A1(n55358), .A2(n53700), .ZN(n55357) );
  NOR2_X2 U36143 ( .A1(n55344), .A2(n53659), .ZN(n55317) );
  OAI21_X2 U36144 ( .B1(n54582), .B2(n54602), .A(n54563), .ZN(n54564) );
  NOR2_X1 U36145 ( .A1(n53812), .A2(w_MuxIMM_SEL), .ZN(n55289) );
  NOR3_X2 U36146 ( .A1(n53946), .A2(n53679), .A3(n55315), .ZN(\DP/ALU0/n112 )
         );
  INV_X2 U36147 ( .A(n54355), .ZN(n55308) );
  NAND3_X2 U36148 ( .A1(n53810), .A2(\DP/ALU0/s_LOGIC[2] ), .A3(n53611), .ZN(
        n55187) );
  NOR3_X2 U36149 ( .A1(n54507), .A2(n54506), .A3(n54598), .ZN(n54599) );
  AND2_X2 U36150 ( .A1(n55361), .A2(n53790), .ZN(n55359) );
  AND2_X2 U36151 ( .A1(n55357), .A2(n53767), .ZN(n55361) );
  NOR2_X1 U36152 ( .A1(n55341), .A2(n53656), .ZN(n55345) );
  NOR2_X1 U36153 ( .A1(n55338), .A2(n53657), .ZN(n55342) );
  NAND4_X1 U36154 ( .A1(w_MuxIMM_SEL), .A2(n55290), .A3(w_SIGN_EN), .A4(n53704), .ZN(n55292) );
  NOR2_X2 U36155 ( .A1(n55290), .A2(n55289), .ZN(n55291) );
  NOR2_X1 U36156 ( .A1(n53984), .A2(n54858), .ZN(n53771) );
  NOR2_X1 U36157 ( .A1(n54033), .A2(n54858), .ZN(n53769) );
  NOR2_X1 U36158 ( .A1(n54019), .A2(n54858), .ZN(n53770) );
  XOR2_X1 U36159 ( .A(n53983), .B(\DP/ALU0/s_A_MULT[15] ), .Z(n54860) );
  INV_X1 U36160 ( .A(n54691), .ZN(n54687) );
  NOR2_X1 U36161 ( .A1(n53970), .A2(n54299), .ZN(n54182) );
  NOR2_X1 U36162 ( .A1(n55353), .A2(n53655), .ZN(n55323) );
  INV_X1 U36163 ( .A(n54917), .ZN(n54910) );
  INV_X1 U36164 ( .A(n54807), .ZN(n54803) );
  NOR2_X1 U36165 ( .A1(n53970), .A2(n54184), .ZN(n54300) );
  AOI21_X1 U36166 ( .B1(n53772), .B2(n53773), .A(n53759), .ZN(n53774) );
  INV_X1 U36167 ( .A(n55316), .ZN(n53773) );
  NOR2_X1 U36168 ( .A1(w_ALU_OPCODE[2]), .A2(n53646), .ZN(n53772) );
  NAND2_X1 U36169 ( .A1(\DP/ALU0/S_B_MULT[3] ), .A2(n54478), .ZN(n54916) );
  INV_X1 U36170 ( .A(n54859), .ZN(n54863) );
  INV_X1 U36171 ( .A(n54857), .ZN(n54865) );
  NAND2_X1 U36172 ( .A1(n53958), .A2(n53957), .ZN(n55179) );
  NOR2_X1 U36173 ( .A1(n53368), .A2(n53799), .ZN(n54930) );
  NOR2_X1 U36174 ( .A1(n53379), .A2(n54952), .ZN(n54951) );
  NOR2_X1 U36175 ( .A1(n53414), .A2(n55333), .ZN(n55332) );
  NAND2_X1 U36176 ( .A1(n55357), .A2(w_PC_OUT[25]), .ZN(n55362) );
  NOR2_X1 U36177 ( .A1(n54974), .A2(n53387), .ZN(n54977) );
  NOR2_X1 U36178 ( .A1(n49937), .A2(n53694), .ZN(n54982) );
  NAND2_X1 U36179 ( .A1(n53702), .A2(n53375), .ZN(n53768) );
  NOR2_X1 U36180 ( .A1(n53674), .A2(n53744), .ZN(n53767) );
  NAND2_X1 U36181 ( .A1(n53780), .A2(n53381), .ZN(n53703) );
  AND3_X1 U36182 ( .A1(n53679), .A2(w_ALU_OPCODE[2]), .A3(n53948), .ZN(n53759)
         );
  INV_X1 U36183 ( .A(n54603), .ZN(n53806) );
  AND2_X1 U36184 ( .A1(n54055), .A2(n54032), .ZN(n53764) );
  AND2_X1 U36185 ( .A1(n54055), .A2(n54018), .ZN(n53765) );
  AND2_X1 U36186 ( .A1(n54055), .A2(n53985), .ZN(n53766) );
  NOR2_X1 U36187 ( .A1(n53685), .A2(n53386), .ZN(n54978) );
  MUX2_X1 U36188 ( .A(n53769), .B(n53764), .S(\DP/ALU0/S_B_MULT[7] ), .Z(
        n54035) );
  MUX2_X1 U36189 ( .A(n53770), .B(n53765), .S(\DP/ALU0/S_B_MULT[3] ), .Z(
        n54021) );
  MUX2_X1 U36190 ( .A(n53771), .B(n53766), .S(\DP/ALU0/S_B_MULT[15] ), .Z(
        n54062) );
  NOR2_X1 U36191 ( .A1(n49845), .A2(n53776), .ZN(n53777) );
  OR2_X1 U36192 ( .A1(n53779), .A2(n53657), .ZN(n53778) );
  AND2_X1 U36193 ( .A1(n53795), .A2(n53780), .ZN(n54960) );
  NAND2_X1 U36194 ( .A1(n53795), .A2(n53782), .ZN(n54957) );
  OR2_X1 U36195 ( .A1(n53785), .A2(n53656), .ZN(n53784) );
  OR2_X1 U36196 ( .A1(n53787), .A2(n49937), .ZN(n53786) );
  OR2_X1 U36197 ( .A1(n53789), .A2(n53379), .ZN(n53788) );
  AND2_X1 U36198 ( .A1(n53601), .A2(w_PC_OUT[27]), .ZN(n53790) );
  OR2_X1 U36199 ( .A1(n53792), .A2(n53655), .ZN(n53791) );
  INV_X1 U36200 ( .A(n53793), .ZN(n55295) );
  NAND2_X1 U36201 ( .A1(n55286), .A2(IRAM_ADDR[5]), .ZN(n53793) );
  NOR2_X1 U36202 ( .A1(n54970), .A2(n53385), .ZN(n53795) );
  AND2_X1 U36203 ( .A1(n53795), .A2(n53796), .ZN(n54961) );
  NOR2_X1 U36204 ( .A1(n53385), .A2(n54970), .ZN(n54969) );
  NAND2_X1 U36205 ( .A1(n54932), .A2(n49958), .ZN(n53799) );
  NOR3_X1 U36206 ( .A1(\DP/ALU0/S_B_SHIFT[3] ), .A2(\DP/ALU0/S_B_SHIFT[4] ), 
        .A3(n53970), .ZN(n53802) );
  NOR3_X1 U36207 ( .A1(\DP/ALU0/S_B_SHIFT[3] ), .A2(\DP/ALU0/S_B_SHIFT[4] ), 
        .A3(n53970), .ZN(n53803) );
  NAND2_X1 U36208 ( .A1(w_IR_OUT[27]), .A2(n53651), .ZN(n53837) );
  NAND2_X1 U36209 ( .A1(n53681), .A2(n53653), .ZN(n53886) );
  NAND3_X1 U36210 ( .A1(n53825), .A2(w_IR_OUT[28]), .A3(n53853), .ZN(n53898)
         );
  OAI21_X1 U36211 ( .B1(n53837), .B2(n53886), .A(n53898), .ZN(n32429) );
  NOR2_X1 U36212 ( .A1(n53681), .A2(n53653), .ZN(n53847) );
  NAND3_X1 U36213 ( .A1(n53847), .A2(n53651), .A3(n53683), .ZN(n53900) );
  AOI21_X1 U36214 ( .B1(w_IR_OUT[27]), .B2(n53678), .A(n53900), .ZN(n32415) );
  NAND3_X1 U36215 ( .A1(w_IR_OUT[31]), .A2(n53853), .A3(n53681), .ZN(n55128)
         );
  INV_X1 U36216 ( .A(n55128), .ZN(n53824) );
  NAND2_X1 U36217 ( .A1(w_IR_OUT[31]), .A2(n53681), .ZN(n53823) );
  NOR4_X1 U36218 ( .A1(w_IR_OUT[28]), .A2(w_IR_OUT[30]), .A3(n53823), .A4(
        n53890), .ZN(n53894) );
  NOR3_X1 U36219 ( .A1(n32415), .A2(n53824), .A3(n53894), .ZN(n53872) );
  INV_X1 U36220 ( .A(n53872), .ZN(n49781) );
  NOR2_X1 U36221 ( .A1(n7564), .A2(n53881), .ZN(n53828) );
  NAND3_X1 U36222 ( .A1(n53548), .A2(n53828), .A3(n53687), .ZN(n53856) );
  NOR2_X1 U36223 ( .A1(n53837), .A2(n53683), .ZN(n53875) );
  NAND2_X1 U36224 ( .A1(w_IR_OUT[27]), .A2(n53678), .ZN(n53827) );
  NOR3_X1 U36225 ( .A1(n53886), .A2(n53651), .A3(n53683), .ZN(n53893) );
  INV_X1 U36226 ( .A(n53893), .ZN(n53891) );
  NOR2_X1 U36227 ( .A1(n53826), .A2(n53649), .ZN(n53839) );
  NAND4_X1 U36228 ( .A1(n49853), .A2(n53548), .A3(n7564), .A4(n53839), .ZN(
        n53855) );
  NAND2_X1 U36229 ( .A1(w_IR_OUT[29]), .A2(n53653), .ZN(n53846) );
  NOR2_X1 U36230 ( .A1(n53846), .A2(w_IR_OUT[30]), .ZN(n53895) );
  NAND3_X1 U36231 ( .A1(w_IR_OUT[28]), .A2(n53895), .A3(n53678), .ZN(n53883)
         );
  OAI211_X1 U36232 ( .C1(n53827), .C2(n53891), .A(n53855), .B(n53883), .ZN(
        n53832) );
  NAND3_X1 U36233 ( .A1(n49849), .A2(n53828), .A3(n53649), .ZN(n53879) );
  INV_X1 U36234 ( .A(n32429), .ZN(n55127) );
  NOR2_X1 U36235 ( .A1(w_IR_OUT[28]), .A2(n53846), .ZN(n53871) );
  NAND2_X1 U36236 ( .A1(w_IR_OUT[30]), .A2(n53871), .ZN(n53867) );
  NAND3_X1 U36237 ( .A1(n7616), .A2(n49849), .A3(n53839), .ZN(n53829) );
  NAND2_X1 U36238 ( .A1(n49853), .A2(n7564), .ZN(n53882) );
  OAI22_X1 U36239 ( .A1(w_IR_OUT[26]), .A2(n53867), .B1(n53829), .B2(n53882), 
        .ZN(n53859) );
  AOI211_X1 U36240 ( .C1(n53853), .C2(n53871), .A(n49781), .B(n53859), .ZN(
        n53830) );
  OAI211_X1 U36241 ( .C1(n53879), .C2(n53687), .A(n55127), .B(n53830), .ZN(
        n53831) );
  AOI211_X1 U36242 ( .C1(w_IR_OUT[29]), .C2(n53875), .A(n53832), .B(n53831), 
        .ZN(n53834) );
  NAND2_X1 U36243 ( .A1(n49853), .A2(n53686), .ZN(n53852) );
  NOR2_X1 U36244 ( .A1(n53881), .A2(n53852), .ZN(n53878) );
  NAND3_X1 U36245 ( .A1(n53878), .A2(n7564), .A3(n53649), .ZN(n53833) );
  OAI211_X1 U36246 ( .C1(n53856), .C2(n53652), .A(n53834), .B(n53833), .ZN(
        \CU/aluOpcodei[0] ) );
  NOR2_X1 U36247 ( .A1(n53688), .A2(n53652), .ZN(n53835) );
  AOI211_X1 U36248 ( .C1(n53549), .C2(n53835), .A(n53686), .B(n53882), .ZN(
        n53838) );
  INV_X1 U36249 ( .A(n53838), .ZN(n53851) );
  INV_X1 U36250 ( .A(n53852), .ZN(n53836) );
  NAND3_X1 U36251 ( .A1(n53836), .A2(n53839), .A3(n53689), .ZN(n53854) );
  NOR3_X1 U36252 ( .A1(n7616), .A2(n49849), .A3(n53854), .ZN(n53845) );
  INV_X1 U36253 ( .A(n53895), .ZN(n53887) );
  AOI21_X1 U36254 ( .B1(n53887), .B2(n53867), .A(n53890), .ZN(n53844) );
  NAND4_X1 U36255 ( .A1(w_IR_OUT[28]), .A2(w_IR_OUT[30]), .A3(n53847), .A4(
        n53682), .ZN(n53863) );
  OAI22_X1 U36256 ( .A1(n53837), .A2(n53887), .B1(n53678), .B2(n53863), .ZN(
        n53843) );
  NAND2_X1 U36257 ( .A1(n7564), .A2(n53649), .ZN(n53840) );
  AOI22_X1 U36258 ( .A1(n53878), .A2(n53840), .B1(n53839), .B2(n53838), .ZN(
        n53841) );
  OAI22_X1 U36259 ( .A1(n49853), .A2(n53879), .B1(n53841), .B2(n53652), .ZN(
        n53842) );
  NOR4_X1 U36260 ( .A1(n53845), .A2(n53844), .A3(n53843), .A4(n53842), .ZN(
        n53850) );
  NOR3_X1 U36261 ( .A1(w_IR_OUT[27]), .A2(n53651), .A3(n53846), .ZN(n53870) );
  NAND2_X1 U36262 ( .A1(n53847), .A2(n53875), .ZN(n53864) );
  OAI211_X1 U36263 ( .C1(w_IR_OUT[27]), .C2(n53867), .A(n53891), .B(n53864), 
        .ZN(n53848) );
  OAI21_X1 U36264 ( .B1(n53870), .B2(n53848), .A(n53678), .ZN(n53849) );
  OAI211_X1 U36265 ( .C1(n53851), .C2(n53881), .A(n53850), .B(n53849), .ZN(
        \CU/aluOpcodei[1] ) );
  INV_X1 U36267 ( .A(n53878), .ZN(n53862) );
  NAND2_X1 U36268 ( .A1(n53855), .A2(n53854), .ZN(n53876) );
  AOI21_X1 U36269 ( .B1(n53549), .B2(n53652), .A(n53856), .ZN(n53877) );
  NAND2_X1 U36270 ( .A1(n49849), .A2(n53649), .ZN(n53857) );
  AOI22_X1 U36271 ( .A1(n7616), .A2(n53876), .B1(n53877), .B2(n53857), .ZN(
        n53861) );
  OAI21_X1 U36272 ( .B1(w_IR_OUT[27]), .B2(n53678), .A(n53893), .ZN(n53889) );
  NAND2_X1 U36273 ( .A1(n53898), .A2(n53889), .ZN(n53874) );
  AOI21_X1 U36274 ( .B1(w_IR_OUT[28]), .B2(n53895), .A(n53874), .ZN(n53868) );
  OAI22_X1 U36275 ( .A1(n53868), .A2(n53890), .B1(n53682), .B2(n53867), .ZN(
        n53858) );
  AOI211_X1 U36276 ( .C1(w_IR_OUT[30]), .C2(n53870), .A(n53859), .B(n53858), 
        .ZN(n53860) );
  NAND2_X1 U36277 ( .A1(n53861), .A2(n53860), .ZN(\CU/aluOpcodei[3] ) );
  NAND2_X1 U36278 ( .A1(w_IR_OUT[26]), .A2(n53682), .ZN(n53899) );
  NOR4_X1 U36279 ( .A1(n49849), .A2(n53649), .A3(n53862), .A4(n53689), .ZN(
        n53865) );
  NAND2_X1 U36280 ( .A1(n53864), .A2(n53863), .ZN(n53869) );
  AOI211_X1 U36281 ( .C1(n53688), .C2(n53876), .A(n53865), .B(n53869), .ZN(
        n53866) );
  OAI21_X1 U36282 ( .B1(n53899), .B2(n53867), .A(n53866), .ZN(
        \CU/aluOpcodei[4] ) );
  NOR3_X1 U36283 ( .A1(n53871), .A2(n53870), .A3(n53869), .ZN(n53897) );
  NAND2_X1 U36284 ( .A1(n53897), .A2(n53872), .ZN(n53873) );
  AOI211_X1 U36285 ( .C1(n53875), .C2(n53653), .A(n53874), .B(n53873), .ZN(
        n53884) );
  NAND2_X1 U36286 ( .A1(n53884), .A2(n53887), .ZN(\CU/cw[18] ) );
  NOR3_X1 U36287 ( .A1(n53878), .A2(n53877), .A3(n53876), .ZN(n53880) );
  OAI211_X1 U36288 ( .C1(n53882), .C2(n53881), .A(n53880), .B(n53879), .ZN(
        n3025) );
  INV_X1 U36289 ( .A(n3025), .ZN(n53885) );
  NAND3_X1 U36290 ( .A1(n53885), .A2(n53884), .A3(n53883), .ZN(\CU/cw[20] ) );
  NAND3_X1 U36291 ( .A1(n53897), .A2(n55128), .A3(n53887), .ZN(n53888) );
  NOR4_X1 U36292 ( .A1(n53894), .A2(n45959), .A3(n3025), .A4(n53888), .ZN(
        n53892) );
  NAND2_X1 U36293 ( .A1(n53892), .A2(n53889), .ZN(\CU/n142 ) );
  OR3_X1 U36294 ( .A1(n32415), .A2(n32429), .A3(\CU/n142 ), .ZN(\CU/cw[21] )
         );
  NAND4_X1 U36295 ( .A1(n53892), .A2(n55127), .A3(n53891), .A4(n55329), .ZN(
        \CU/cw[3] ) );
  OR2_X1 U36296 ( .A1(n32415), .A2(n3025), .ZN(n9315) );
  NOR4_X1 U36297 ( .A1(n53895), .A2(n53894), .A3(n53893), .A4(n9315), .ZN(
        n53896) );
  NAND3_X1 U36298 ( .A1(n55127), .A2(n53897), .A3(n53896), .ZN(\CU/cw[6] ) );
  NOR2_X1 U36299 ( .A1(w_IR_OUT[26]), .A2(n53898), .ZN(\CU/n138 ) );
  NOR3_X1 U36300 ( .A1(w_IR_OUT[27]), .A2(w_IR_OUT[26]), .A3(n53900), .ZN(
        \CU/n139 ) );
  NOR2_X1 U36301 ( .A1(n53900), .A2(n53899), .ZN(\CU/n140 ) );
  OR2_X1 U36302 ( .A1(n53692), .A2(w_ALU_OPCODE[3]), .ZN(n53902) );
  NAND2_X1 U36303 ( .A1(w_ALU_OPCODE[3]), .A2(n53692), .ZN(n53946) );
  NOR2_X1 U36304 ( .A1(w_ALU_OPCODE[1]), .A2(n53680), .ZN(n53943) );
  INV_X1 U36305 ( .A(n53943), .ZN(n53901) );
  OAI22_X1 U36306 ( .A1(w_ALU_OPCODE[2]), .A2(n53902), .B1(n53946), .B2(n53901), .ZN(n55158) );
  NOR2_X1 U36307 ( .A1(n53946), .A2(n53679), .ZN(n53904) );
  NAND2_X1 U36308 ( .A1(n53646), .A2(n53680), .ZN(n55315) );
  NOR2_X1 U36309 ( .A1(n53646), .A2(n53680), .ZN(n53941) );
  NOR4_X1 U36310 ( .A1(w_ALU_OPCODE[3]), .A2(w_ALU_OPCODE[1]), .A3(n53941), 
        .A4(n53692), .ZN(n53903) );
  AOI21_X1 U36311 ( .B1(n53904), .B2(n55315), .A(n53903), .ZN(n55163) );
  INV_X1 U36312 ( .A(n55163), .ZN(n53905) );
  NOR2_X1 U36313 ( .A1(n55158), .A2(n53905), .ZN(n55314) );
  INV_X1 U36314 ( .A(n55314), .ZN(n51572) );
  NOR2_X1 U36315 ( .A1(w_ALU_OPCODE[2]), .A2(w_ALU_OPCODE[1]), .ZN(n55161) );
  NAND2_X1 U36316 ( .A1(w_ALU_OPCODE[0]), .A2(n55161), .ZN(n53945) );
  NOR2_X1 U36317 ( .A1(w_ALU_OPCODE[3]), .A2(w_ALU_OPCODE[4]), .ZN(n53948) );
  INV_X1 U36318 ( .A(n53948), .ZN(n53906) );
  NAND2_X1 U36319 ( .A1(w_ALU_OPCODE[1]), .A2(n53948), .ZN(n55316) );
  OAI22_X1 U36320 ( .A1(n53945), .A2(n53906), .B1(n55316), .B2(n55315), .ZN(
        n53974) );
  NAND4_X1 U36321 ( .A1(n53261), .A2(n7679), .A3(n7286), .A4(n22592), .ZN(
        n53907) );
  NOR2_X1 U36322 ( .A1(n3214), .A2(n53907), .ZN(n53918) );
  OAI221_X1 U36323 ( .B1(n49857), .B2(n7679), .C1(n53673), .C2(n3253), .A(
        w_RF_WE3), .ZN(n53912) );
  AOI22_X1 U36324 ( .A1(n49819), .A2(n22592), .B1(n53515), .B2(n53261), .ZN(
        n53908) );
  OAI221_X1 U36325 ( .B1(n49819), .B2(n22592), .C1(n53515), .C2(n53261), .A(
        n53908), .ZN(n53911) );
  AOI22_X1 U36326 ( .A1(n49866), .A2(n7286), .B1(n53753), .B2(n37948), .ZN(
        n53909) );
  OAI221_X1 U36327 ( .B1(n49866), .B2(n7286), .C1(n53753), .C2(n37948), .A(
        n53909), .ZN(n53910) );
  OAI221_X1 U36328 ( .B1(n3015), .B2(n3214), .C1(\DP/RD4[2] ), .C2(n37948), 
        .A(w_RF_WE4), .ZN(n53917) );
  AOI22_X1 U36329 ( .A1(\DP/RD4[0] ), .A2(n7679), .B1(\DP/RD4[3] ), .B2(n7286), 
        .ZN(n53913) );
  OAI221_X1 U36330 ( .B1(\DP/RD4[0] ), .B2(n7679), .C1(\DP/RD4[3] ), .C2(n7286), .A(n53913), .ZN(n53916) );
  AOI22_X1 U36331 ( .A1(\DP/RD4[4] ), .A2(n53261), .B1(n22592), .B2(
        \DP/RD4[1] ), .ZN(n53914) );
  OAI221_X1 U36332 ( .B1(\DP/RD4[4] ), .B2(n53261), .C1(\DP/RD4[1] ), .C2(
        n22592), .A(n53914), .ZN(n53915) );
  NOR4_X1 U36333 ( .A1(n53918), .A2(n53917), .A3(n53916), .A4(n53915), .ZN(
        n53922) );
  NOR2_X1 U36334 ( .A1(n55121), .A2(n53922), .ZN(n53923) );
  NOR3_X1 U36335 ( .A1(w_MuxLD_SEL[0]), .A2(w_MuxLD_SEL[1]), .A3(n53654), .ZN(
        n54501) );
  NAND3_X1 U36336 ( .A1(n54501), .A2(n49869), .A3(w_SIGN_LD_EN), .ZN(n53919)
         );
  NAND3_X1 U36337 ( .A1(n53654), .A2(n53701), .A3(w_MuxLD_SEL[0]), .ZN(n54530)
         );
  AOI21_X1 U36338 ( .B1(n53260), .B2(n54548), .A(n54547), .ZN(n53921) );
  OAI21_X1 U36339 ( .B1(n53647), .B2(n53259), .A(n53921), .ZN(n55215) );
  INV_X1 U36340 ( .A(n55215), .ZN(n54510) );
  NAND2_X1 U36341 ( .A1(n55103), .A2(n53922), .ZN(n55077) );
  AOI22_X1 U36342 ( .A1(n7626), .A2(n55121), .B1(n54510), .B2(n55122), .ZN(
        n53924) );
  OAI211_X1 U36343 ( .C1(n53450), .C2(n55126), .A(n53924), .B(n55124), .ZN(
        n3108) );
  NAND4_X1 U36344 ( .A1(n49913), .A2(n53264), .A3(n53265), .A4(n49917), .ZN(
        n53925) );
  NOR2_X1 U36345 ( .A1(n53754), .A2(n53925), .ZN(n53936) );
  OAI221_X1 U36346 ( .B1(n49857), .B2(n53264), .C1(n53673), .C2(n53758), .A(
        w_RF_WE3), .ZN(n53930) );
  AOI22_X1 U36347 ( .A1(n49819), .A2(n49913), .B1(n53515), .B2(n49917), .ZN(
        n53926) );
  OAI221_X1 U36348 ( .B1(n49819), .B2(n49913), .C1(n53515), .C2(n49917), .A(
        n53926), .ZN(n53929) );
  AOI22_X1 U36349 ( .A1(n49866), .A2(n53263), .B1(n53753), .B2(n53265), .ZN(
        n53927) );
  OAI221_X1 U36350 ( .B1(n49866), .B2(n53263), .C1(n53753), .C2(n53265), .A(
        n53927), .ZN(n53928) );
  OAI221_X1 U36351 ( .B1(n49659), .B2(n53754), .C1(\DP/RD4[3] ), .C2(n53263), 
        .A(w_RF_WE4), .ZN(n53935) );
  AOI22_X1 U36352 ( .A1(\DP/RD4[1] ), .A2(n49913), .B1(\DP/RD4[0] ), .B2(
        n53264), .ZN(n53931) );
  OAI221_X1 U36353 ( .B1(\DP/RD4[1] ), .B2(n49913), .C1(\DP/RD4[0] ), .C2(
        n53264), .A(n53931), .ZN(n53934) );
  AOI22_X1 U36354 ( .A1(\DP/RD4[2] ), .A2(n53265), .B1(n49917), .B2(
        \DP/RD4[4] ), .ZN(n53932) );
  OAI221_X1 U36355 ( .B1(\DP/RD4[2] ), .B2(n53265), .C1(\DP/RD4[4] ), .C2(
        n49917), .A(n53932), .ZN(n53933) );
  NOR4_X1 U36356 ( .A1(n53936), .A2(n53935), .A3(n53934), .A4(n53933), .ZN(
        n53938) );
  NOR2_X1 U36357 ( .A1(n55099), .A2(n53938), .ZN(n53937) );
  OAI22_X1 U36358 ( .A1(n53664), .A2(n55116), .B1(n55215), .B2(n55115), .ZN(
        n53939) );
  AOI21_X1 U36359 ( .B1(n53482), .B2(n55118), .A(n53939), .ZN(n53940) );
  OAI21_X1 U36360 ( .B1(n53513), .B2(n55120), .A(n53940), .ZN(n3107) );
  INV_X1 U36361 ( .A(n53941), .ZN(n54926) );
  AND3_X1 U36362 ( .A1(n55315), .A2(n54926), .A3(w_ALU_OPCODE[1]), .ZN(n53942)
         );
  OAI22_X1 U36363 ( .A1(n53943), .A2(n53942), .B1(n3108), .B2(n3107), .ZN(
        n53944) );
  AOI211_X1 U36364 ( .C1(n3107), .C2(n3108), .A(n53946), .B(n53944), .ZN(
        \DP/ALU0/N27 ) );
  NOR2_X1 U36365 ( .A1(n55316), .A2(n54926), .ZN(\DP/ALU0/n114 ) );
  NOR3_X1 U36366 ( .A1(w_ALU_OPCODE[1]), .A2(n53946), .A3(n55315), .ZN(n5402)
         );
  INV_X1 U36367 ( .A(n5402), .ZN(n53947) );
  NAND2_X1 U36368 ( .A1(RST), .A2(n3020), .ZN(n5463) );
  XOR2_X1 U36369 ( .A(n53955), .B(\DP/ALU0/S_B_SHIFT[0] ), .Z(n53967) );
  INV_X1 U36370 ( .A(n53967), .ZN(n53949) );
  INV_X1 U36371 ( .A(\DP/ALU0/s_SHIFT[1] ), .ZN(n53950) );
  INV_X1 U36372 ( .A(\DP/ALU0/s_A_SHIFT[31] ), .ZN(n54303) );
  NOR3_X1 U36373 ( .A1(\DP/ALU0/s_SHIFT[0] ), .A2(n53950), .A3(n54303), .ZN(
        n53968) );
  NOR2_X1 U36374 ( .A1(n53968), .A2(\DP/ALU0/s_A_SHIFT[16] ), .ZN(n53954) );
  INV_X1 U36375 ( .A(\DP/ALU0/S_B_SHIFT[3] ), .ZN(n53951) );
  NOR2_X1 U36376 ( .A1(\DP/ALU0/S_B_SHIFT[4] ), .A2(n53951), .ZN(n53969) );
  OAI21_X1 U36377 ( .B1(n53955), .B2(n53968), .A(n53969), .ZN(n54064) );
  INV_X1 U36378 ( .A(n53955), .ZN(n53970) );
  NOR3_X1 U36379 ( .A1(\DP/ALU0/S_B_SHIFT[3] ), .A2(\DP/ALU0/S_B_SHIFT[4] ), 
        .A3(n53970), .ZN(n54421) );
  INV_X1 U36380 ( .A(n53968), .ZN(n54100) );
  NAND2_X1 U36381 ( .A1(\DP/ALU0/S_B_SHIFT[4] ), .A2(n53951), .ZN(n54299) );
  NOR2_X1 U36382 ( .A1(n54100), .A2(n54299), .ZN(n54255) );
  AOI21_X1 U36383 ( .B1(n53803), .B2(\DP/ALU0/s_A_SHIFT[24] ), .A(n54255), 
        .ZN(n53953) );
  INV_X1 U36384 ( .A(\DP/ALU0/S_B_SHIFT[4] ), .ZN(n53963) );
  AOI21_X1 U36385 ( .B1(\DP/ALU0/s_SHIFT[0] ), .B2(\DP/ALU0/s_SHIFT[1] ), .A(
        n53955), .ZN(n54183) );
  NAND3_X1 U36386 ( .A1(n53951), .A2(n53963), .A3(n54183), .ZN(n54411) );
  AOI22_X1 U36387 ( .A1(\DP/ALU0/s_A_SHIFT[31] ), .A2(n55175), .B1(n54182), 
        .B2(\DP/ALU0/s_A_SHIFT[8] ), .ZN(n53952) );
  OAI211_X1 U36388 ( .C1(n53954), .C2(n54064), .A(n53953), .B(n53952), .ZN(
        n54157) );
  XNOR2_X1 U36389 ( .A(n53955), .B(\DP/ALU0/S_B_SHIFT[1] ), .ZN(n53958) );
  XOR2_X1 U36390 ( .A(n53955), .B(\DP/ALU0/S_B_SHIFT[2] ), .Z(n53956) );
  INV_X1 U36391 ( .A(n53956), .ZN(n53957) );
  NAND2_X1 U36392 ( .A1(n53958), .A2(n53956), .ZN(n55177) );
  INV_X1 U36393 ( .A(\DP/ALU0/s_A_SHIFT[12] ), .ZN(n54241) );
  NAND2_X1 U36394 ( .A1(n54100), .A2(n54241), .ZN(n54122) );
  INV_X1 U36395 ( .A(n54182), .ZN(n54101) );
  AOI22_X1 U36396 ( .A1(\DP/ALU0/S_B_SHIFT[3] ), .A2(\DP/ALU0/S_B_SHIFT[4] ), 
        .B1(n54100), .B2(n54101), .ZN(n53972) );
  INV_X1 U36397 ( .A(n54064), .ZN(n53971) );
  AOI222_X1 U36398 ( .A1(n54122), .A2(n53972), .B1(n53802), .B2(
        \DP/ALU0/s_A_SHIFT[28] ), .C1(\DP/ALU0/s_A_SHIFT[20] ), .C2(n53971), 
        .ZN(n54079) );
  INV_X1 U36399 ( .A(\DP/ALU0/s_A_SHIFT[10] ), .ZN(n54375) );
  NAND2_X1 U36400 ( .A1(n54100), .A2(n54375), .ZN(n54151) );
  AOI222_X1 U36401 ( .A1(n54151), .A2(n53972), .B1(n53803), .B2(
        \DP/ALU0/s_A_SHIFT[26] ), .C1(n53971), .C2(\DP/ALU0/s_A_SHIFT[18] ), 
        .ZN(n54121) );
  AOI22_X1 U36402 ( .A1(n55137), .A2(n54079), .B1(n53807), .B2(n54121), .ZN(
        n53962) );
  NOR2_X1 U36403 ( .A1(n53968), .A2(\DP/ALU0/s_A_SHIFT[14] ), .ZN(n54081) );
  INV_X1 U36404 ( .A(n53972), .ZN(n53960) );
  AOI22_X1 U36405 ( .A1(n53971), .A2(\DP/ALU0/s_A_SHIFT[22] ), .B1(n53802), 
        .B2(\DP/ALU0/s_A_SHIFT[30] ), .ZN(n53959) );
  OAI211_X1 U36406 ( .C1(n54081), .C2(n53960), .A(n53804), .B(n53959), .ZN(
        n53961) );
  OAI211_X1 U36407 ( .C1(n54157), .C2(n55179), .A(n53962), .B(n53961), .ZN(
        n54078) );
  INV_X1 U36408 ( .A(\DP/ALU0/s_A_SHIFT[9] ), .ZN(n54393) );
  NAND2_X1 U36409 ( .A1(n54100), .A2(n54393), .ZN(n54167) );
  AOI222_X1 U36410 ( .A1(n54167), .A2(n53972), .B1(n54421), .B2(
        \DP/ALU0/s_A_SHIFT[25] ), .C1(n53971), .C2(\DP/ALU0/s_A_SHIFT[17] ), 
        .ZN(n54140) );
  AOI221_X1 U36411 ( .B1(\DP/ALU0/s_A_SHIFT[13] ), .B2(\DP/ALU0/S_B_SHIFT[4] ), 
        .C1(\DP/ALU0/s_A_SHIFT[29] ), .C2(n53963), .A(n53968), .ZN(n53964) );
  OAI22_X1 U36412 ( .A1(\DP/ALU0/S_B_SHIFT[4] ), .A2(n54100), .B1(
        \DP/ALU0/S_B_SHIFT[3] ), .B2(n53964), .ZN(n53966) );
  NAND2_X1 U36413 ( .A1(n53970), .A2(n54100), .ZN(n53965) );
  OAI221_X1 U36414 ( .B1(n53966), .B2(n53969), .C1(n53966), .C2(
        \DP/ALU0/s_A_SHIFT[21] ), .A(n53965), .ZN(n54070) );
  OAI22_X1 U36415 ( .A1(n54140), .A2(n55179), .B1(n55177), .B2(n54070), .ZN(
        n53981) );
  OR2_X1 U36416 ( .A1(n53968), .A2(\DP/ALU0/s_A_SHIFT[15] ), .ZN(n54065) );
  INV_X1 U36417 ( .A(n53969), .ZN(n54184) );
  AOI222_X1 U36418 ( .A1(n54065), .A2(n53972), .B1(n54300), .B2(
        \DP/ALU0/s_A_SHIFT[23] ), .C1(\DP/ALU0/s_A_SHIFT[31] ), .C2(n54421), 
        .ZN(n53973) );
  INV_X1 U36419 ( .A(\DP/ALU0/s_A_SHIFT[11] ), .ZN(n54362) );
  NAND2_X1 U36420 ( .A1(n54100), .A2(n54362), .ZN(n54136) );
  AOI222_X1 U36421 ( .A1(n54136), .A2(n53972), .B1(n53803), .B2(
        \DP/ALU0/s_A_SHIFT[27] ), .C1(n53971), .C2(\DP/ALU0/s_A_SHIFT[19] ), 
        .ZN(n54104) );
  OAI22_X1 U36422 ( .A1(n53973), .A2(n53761), .B1(n54104), .B2(n53760), .ZN(
        n53980) );
  AOI22_X1 U36423 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[15] ), .B1(n7626), .B2(
        n54286), .ZN(n53978) );
  NAND2_X1 U36424 ( .A1(\DP/ALU0/S_B_LOGIC[31] ), .A2(\DP/ALU0/s_A_LOGIC[31] ), 
        .ZN(n53976) );
  NAND3_X1 U36425 ( .A1(n53810), .A2(\DP/ALU0/s_LOGIC[3] ), .A3(n53611), .ZN(
        n54355) );
  NAND2_X1 U36426 ( .A1(n55187), .A2(n53976), .ZN(n53975) );
  OAI221_X1 U36427 ( .B1(n53976), .B2(n55308), .C1(\DP/ALU0/S_B_LOGIC[31] ), 
        .C2(\DP/ALU0/s_A_LOGIC[31] ), .A(n53975), .ZN(n53977) );
  OAI211_X1 U36428 ( .C1(\intadd_8/SUM[3] ), .C2(n55303), .A(n53978), .B(
        n53977), .ZN(n53979) );
  AOI221_X1 U36429 ( .B1(n53981), .B2(n55306), .C1(n53980), .C2(n55306), .A(
        n53979), .ZN(n54063) );
  INV_X1 U36430 ( .A(\DP/ALU0/s_A_MULT[12] ), .ZN(n54621) );
  NOR3_X1 U36431 ( .A1(\DP/ALU0/s_A_MULT[2] ), .A2(\DP/ALU0/s_A_MULT[0] ), 
        .A3(\DP/ALU0/s_A_MULT[1] ), .ZN(n54630) );
  INV_X1 U36432 ( .A(\DP/ALU0/s_A_MULT[3] ), .ZN(n54629) );
  NAND2_X1 U36433 ( .A1(n54630), .A2(n54629), .ZN(n54634) );
  NOR2_X1 U36434 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54634), .ZN(n54633) );
  INV_X1 U36435 ( .A(n54633), .ZN(n54638) );
  NOR2_X1 U36436 ( .A1(n54638), .A2(\DP/ALU0/s_A_MULT[5] ), .ZN(n54637) );
  INV_X1 U36437 ( .A(n54637), .ZN(n54642) );
  NOR2_X1 U36438 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54642), .ZN(n54641) );
  INV_X1 U36439 ( .A(n54641), .ZN(n54646) );
  NOR2_X1 U36440 ( .A1(n54646), .A2(\DP/ALU0/s_A_MULT[7] ), .ZN(n54645) );
  INV_X1 U36441 ( .A(n54645), .ZN(n54650) );
  NOR2_X1 U36442 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54650), .ZN(n54649) );
  INV_X1 U36443 ( .A(n54649), .ZN(n54654) );
  NOR2_X1 U36444 ( .A1(n54654), .A2(\DP/ALU0/s_A_MULT[9] ), .ZN(n54653) );
  INV_X1 U36445 ( .A(n54653), .ZN(n54617) );
  NOR2_X1 U36446 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n54617), .ZN(n54616) );
  INV_X1 U36447 ( .A(n54616), .ZN(n54615) );
  NOR2_X1 U36448 ( .A1(n54615), .A2(\DP/ALU0/s_A_MULT[11] ), .ZN(n54622) );
  NAND2_X1 U36449 ( .A1(n54621), .A2(n54622), .ZN(n54620) );
  NOR2_X1 U36450 ( .A1(n54620), .A2(\DP/ALU0/s_A_MULT[13] ), .ZN(n53989) );
  INV_X1 U36451 ( .A(n53989), .ZN(n53982) );
  NOR2_X1 U36452 ( .A1(\DP/ALU0/s_A_MULT[14] ), .A2(n53982), .ZN(n53983) );
  INV_X1 U36453 ( .A(n54860), .ZN(n54055) );
  NAND2_X1 U36454 ( .A1(\DP/ALU0/S_B_MULT[13] ), .A2(\DP/ALU0/S_B_MULT[14] ), 
        .ZN(n53985) );
  INV_X1 U36455 ( .A(\DP/ALU0/S_B_MULT[15] ), .ZN(n53986) );
  NOR2_X1 U36456 ( .A1(\DP/ALU0/S_B_MULT[13] ), .A2(\DP/ALU0/S_B_MULT[14] ), 
        .ZN(n53984) );
  INV_X1 U36457 ( .A(\DP/ALU0/s_A_MULT[15] ), .ZN(n54858) );
  AOI21_X1 U36458 ( .B1(\DP/ALU0/S_B_MULT[14] ), .B2(\DP/ALU0/S_B_MULT[13] ), 
        .A(n53984), .ZN(n54313) );
  NAND2_X1 U36459 ( .A1(\DP/ALU0/S_B_MULT[15] ), .A2(n54313), .ZN(n54664) );
  INV_X1 U36460 ( .A(n54313), .ZN(n54312) );
  AOI22_X1 U36461 ( .A1(\DP/ALU0/s_A_MULT[14] ), .A2(n54659), .B1(
        \DP/ALU0/s_A_MULT[15] ), .B2(n54661), .ZN(n53988) );
  XOR2_X1 U36462 ( .A(n53989), .B(\DP/ALU0/s_A_MULT[14] ), .Z(n54043) );
  INV_X1 U36463 ( .A(n54043), .ZN(n54862) );
  NAND2_X1 U36464 ( .A1(n54862), .A2(n53642), .ZN(n53987) );
  OAI211_X1 U36465 ( .C1(n54860), .C2(n54664), .A(n53988), .B(n53987), .ZN(
        n54090) );
  AOI22_X1 U36466 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54659), .B1(
        \DP/ALU0/s_A_MULT[14] ), .B2(n54661), .ZN(n53991) );
  NAND2_X1 U36467 ( .A1(n54856), .A2(n53642), .ZN(n53990) );
  OAI211_X1 U36468 ( .C1(n54664), .C2(n54043), .A(n53991), .B(n53990), .ZN(
        n54058) );
  NOR2_X1 U36469 ( .A1(\intadd_1/n1 ), .A2(n54058), .ZN(n54108) );
  NOR2_X1 U36470 ( .A1(\DP/ALU0/S_B_MULT[11] ), .A2(\DP/ALU0/S_B_MULT[12] ), 
        .ZN(n54056) );
  AOI21_X1 U36471 ( .B1(\DP/ALU0/S_B_MULT[12] ), .B2(\DP/ALU0/S_B_MULT[11] ), 
        .A(n54056), .ZN(n54342) );
  NAND2_X1 U36472 ( .A1(\DP/ALU0/S_B_MULT[13] ), .A2(n54342), .ZN(n54690) );
  NAND2_X1 U36473 ( .A1(\DP/ALU0/S_B_MULT[11] ), .A2(\DP/ALU0/S_B_MULT[12] ), 
        .ZN(n54054) );
  INV_X1 U36474 ( .A(\DP/ALU0/S_B_MULT[13] ), .ZN(n54057) );
  NAND2_X1 U36475 ( .A1(n54057), .A2(n54342), .ZN(n54691) );
  AOI22_X1 U36476 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54693), .B1(
        \DP/ALU0/s_A_MULT[14] ), .B2(n54687), .ZN(n53993) );
  NAND2_X1 U36477 ( .A1(n54856), .A2(n53644), .ZN(n53992) );
  OAI211_X1 U36478 ( .C1(n54043), .C2(n54690), .A(n53993), .B(n53992), .ZN(
        n54608) );
  AOI22_X1 U36479 ( .A1(\DP/ALU0/s_A_MULT[14] ), .A2(n54693), .B1(
        \DP/ALU0/s_A_MULT[15] ), .B2(n54687), .ZN(n53995) );
  NAND2_X1 U36480 ( .A1(n54862), .A2(n53644), .ZN(n53994) );
  OAI211_X1 U36481 ( .C1(n54860), .C2(n54690), .A(n53995), .B(n53994), .ZN(
        n54613) );
  NOR2_X1 U36482 ( .A1(\DP/ALU0/S_B_MULT[9] ), .A2(\DP/ALU0/S_B_MULT[10] ), 
        .ZN(n54049) );
  NOR2_X1 U36483 ( .A1(\DP/ALU0/S_B_MULT[11] ), .A2(n54049), .ZN(n53996) );
  INV_X1 U36484 ( .A(\DP/ALU0/S_B_MULT[11] ), .ZN(n54039) );
  AOI211_X1 U36485 ( .C1(\DP/ALU0/S_B_MULT[9] ), .C2(\DP/ALU0/S_B_MULT[10] ), 
        .A(n54860), .B(n54039), .ZN(n54046) );
  AOI21_X1 U36486 ( .B1(n53996), .B2(\DP/ALU0/s_A_MULT[15] ), .A(n54046), .ZN(
        n54053) );
  NAND2_X1 U36487 ( .A1(\DP/ALU0/S_B_MULT[7] ), .A2(\DP/ALU0/S_B_MULT[8] ), 
        .ZN(n54037) );
  OAI21_X1 U36488 ( .B1(\DP/ALU0/S_B_MULT[7] ), .B2(\DP/ALU0/S_B_MULT[8] ), 
        .A(n54037), .ZN(n54403) );
  INV_X1 U36489 ( .A(n54403), .ZN(n54404) );
  NAND2_X1 U36490 ( .A1(\DP/ALU0/S_B_MULT[9] ), .A2(n54404), .ZN(n54780) );
  INV_X1 U36491 ( .A(\DP/ALU0/S_B_MULT[9] ), .ZN(n54038) );
  AOI22_X1 U36492 ( .A1(\DP/ALU0/s_A_MULT[14] ), .A2(n54775), .B1(n54862), 
        .B2(n53640), .ZN(n53997) );
  OAI21_X1 U36493 ( .B1(n54860), .B2(n54780), .A(n53997), .ZN(n53998) );
  AOI21_X1 U36494 ( .B1(\DP/ALU0/s_A_MULT[15] ), .B2(n54777), .A(n53998), .ZN(
        n54741) );
  AOI22_X1 U36495 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54775), .B1(
        \DP/ALU0/s_A_MULT[14] ), .B2(n54777), .ZN(n54000) );
  NAND2_X1 U36496 ( .A1(n54856), .A2(n53640), .ZN(n53999) );
  OAI211_X1 U36497 ( .C1(n54780), .C2(n54043), .A(n54000), .B(n53999), .ZN(
        n54740) );
  INV_X1 U36498 ( .A(n54740), .ZN(n54736) );
  NOR2_X1 U36499 ( .A1(\DP/ALU0/S_B_MULT[5] ), .A2(\DP/ALU0/S_B_MULT[6] ), 
        .ZN(n54033) );
  AOI21_X1 U36500 ( .B1(\DP/ALU0/S_B_MULT[6] ), .B2(\DP/ALU0/S_B_MULT[5] ), 
        .A(n54033), .ZN(n54437) );
  NAND2_X1 U36501 ( .A1(\DP/ALU0/S_B_MULT[7] ), .A2(n54437), .ZN(n54806) );
  NAND2_X1 U36502 ( .A1(\DP/ALU0/S_B_MULT[5] ), .A2(\DP/ALU0/S_B_MULT[6] ), 
        .ZN(n54032) );
  INV_X1 U36503 ( .A(\DP/ALU0/S_B_MULT[7] ), .ZN(n54034) );
  NAND2_X1 U36504 ( .A1(n54034), .A2(n54437), .ZN(n54807) );
  AOI22_X1 U36505 ( .A1(\DP/ALU0/s_A_MULT[14] ), .A2(n54809), .B1(
        \DP/ALU0/s_A_MULT[15] ), .B2(n54803), .ZN(n54002) );
  NAND2_X1 U36506 ( .A1(n54862), .A2(n53641), .ZN(n54001) );
  OAI211_X1 U36507 ( .C1(n54860), .C2(n54806), .A(n54002), .B(n54001), .ZN(
        n54749) );
  AOI22_X1 U36508 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54809), .B1(
        \DP/ALU0/s_A_MULT[14] ), .B2(n54803), .ZN(n54003) );
  OAI21_X1 U36509 ( .B1(n54043), .B2(n54806), .A(n54003), .ZN(n54004) );
  AOI21_X1 U36510 ( .B1(n54856), .B2(n53641), .A(n54004), .ZN(n54744) );
  INV_X1 U36511 ( .A(\DP/ALU0/S_B_MULT[5] ), .ZN(n54005) );
  OR2_X1 U36512 ( .A1(\DP/ALU0/S_B_MULT[3] ), .A2(\DP/ALU0/S_B_MULT[4] ), .ZN(
        n54006) );
  NAND2_X1 U36513 ( .A1(\DP/ALU0/S_B_MULT[3] ), .A2(\DP/ALU0/S_B_MULT[4] ), 
        .ZN(n54025) );
  NAND2_X1 U36514 ( .A1(n54006), .A2(n54025), .ZN(n55298) );
  NAND3_X1 U36515 ( .A1(n54006), .A2(n54005), .A3(\DP/ALU0/s_A_MULT[15] ), 
        .ZN(n54026) );
  INV_X1 U36516 ( .A(n54026), .ZN(n54007) );
  AOI22_X1 U36517 ( .A1(\DP/ALU0/s_A_MULT[14] ), .A2(n54849), .B1(n54007), 
        .B2(n54025), .ZN(n54008) );
  OAI21_X1 U36518 ( .B1(n54043), .B2(n54846), .A(n54008), .ZN(n54009) );
  AOI21_X1 U36519 ( .B1(n54850), .B2(n54055), .A(n54009), .ZN(n54815) );
  INV_X1 U36520 ( .A(n54850), .ZN(n54012) );
  AOI22_X1 U36521 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54849), .B1(
        \DP/ALU0/s_A_MULT[14] ), .B2(n54851), .ZN(n54011) );
  NAND2_X1 U36522 ( .A1(n54856), .A2(n53639), .ZN(n54010) );
  OAI211_X1 U36523 ( .C1(n54043), .C2(n54012), .A(n54011), .B(n54010), .ZN(
        n54923) );
  NAND2_X1 U36524 ( .A1(\intadd_6/n1 ), .A2(n54923), .ZN(n54922) );
  NAND2_X1 U36525 ( .A1(\DP/ALU0/S_B_MULT[1] ), .A2(\DP/ALU0/S_B_MULT[2] ), 
        .ZN(n54018) );
  NOR2_X1 U36526 ( .A1(\DP/ALU0/S_B_MULT[1] ), .A2(\DP/ALU0/S_B_MULT[2] ), 
        .ZN(n54019) );
  AOI21_X1 U36527 ( .B1(\DP/ALU0/S_B_MULT[2] ), .B2(\DP/ALU0/S_B_MULT[1] ), 
        .A(n54019), .ZN(n54478) );
  INV_X1 U36528 ( .A(\DP/ALU0/S_B_MULT[3] ), .ZN(n54020) );
  NAND2_X1 U36529 ( .A1(n54020), .A2(n54478), .ZN(n54917) );
  AOI22_X1 U36530 ( .A1(\DP/ALU0/s_A_MULT[14] ), .A2(n54910), .B1(n54856), 
        .B2(n53643), .ZN(n54013) );
  OAI21_X1 U36531 ( .B1(n54043), .B2(n54916), .A(n54013), .ZN(n54014) );
  AOI21_X1 U36532 ( .B1(\DP/ALU0/s_A_MULT[13] ), .B2(n54920), .A(n54014), .ZN(
        n54819) );
  AOI22_X1 U36533 ( .A1(\DP/ALU0/s_A_MULT[14] ), .A2(n54920), .B1(
        \DP/ALU0/s_A_MULT[15] ), .B2(n54910), .ZN(n54016) );
  NAND2_X1 U36534 ( .A1(n54862), .A2(n53643), .ZN(n54015) );
  OAI211_X1 U36535 ( .C1(n54860), .C2(n54916), .A(n54016), .B(n54015), .ZN(
        n54822) );
  INV_X1 U36536 ( .A(\DP/ALU0/S_B_MULT[1] ), .ZN(n54854) );
  NAND2_X1 U36537 ( .A1(\DP/ALU0/S_B_MULT[0] ), .A2(n54854), .ZN(n54857) );
  OAI22_X1 U36538 ( .A1(n54860), .A2(n54854), .B1(n54858), .B2(n54857), .ZN(
        n54817) );
  NOR2_X1 U36539 ( .A1(n54819), .A2(n54817), .ZN(n54816) );
  AOI21_X1 U36540 ( .B1(\intadd_7/n1 ), .B2(n54817), .A(n54816), .ZN(n54820)
         );
  AOI21_X1 U36541 ( .B1(\intadd_7/n1 ), .B2(n54822), .A(n54820), .ZN(n54017)
         );
  OAI21_X1 U36542 ( .B1(n54819), .B2(n54822), .A(n54017), .ZN(n54022) );
  XNOR2_X1 U36543 ( .A(n54022), .B(n54021), .ZN(n54925) );
  NOR2_X1 U36544 ( .A1(n54922), .A2(n54925), .ZN(n54813) );
  NOR2_X1 U36545 ( .A1(\intadd_6/n1 ), .A2(n54923), .ZN(n54023) );
  NAND2_X1 U36546 ( .A1(n54023), .A2(n54925), .ZN(n54811) );
  NAND2_X1 U36547 ( .A1(n54815), .A2(n54811), .ZN(n54024) );
  OAI21_X1 U36548 ( .B1(n54815), .B2(n54813), .A(n54024), .ZN(n54029) );
  NAND3_X1 U36549 ( .A1(n54055), .A2(\DP/ALU0/S_B_MULT[5] ), .A3(n54025), .ZN(
        n54027) );
  NAND2_X1 U36550 ( .A1(n54027), .A2(n54026), .ZN(n54028) );
  XNOR2_X1 U36551 ( .A(n54029), .B(n54028), .ZN(n54745) );
  NAND2_X1 U36552 ( .A1(n54745), .A2(n54744), .ZN(n54030) );
  OAI21_X1 U36553 ( .B1(n54745), .B2(\intadd_5/n1 ), .A(n54030), .ZN(n54747)
         );
  OAI21_X1 U36554 ( .B1(\intadd_5/n1 ), .B2(n54749), .A(n54747), .ZN(n54031)
         );
  AOI21_X1 U36555 ( .B1(n54749), .B2(n54744), .A(n54031), .ZN(n54036) );
  XNOR2_X1 U36556 ( .A(n54036), .B(n54035), .ZN(n54735) );
  MUX2_X1 U36557 ( .A(n54736), .B(\intadd_4/n1 ), .S(n54735), .Z(n54738) );
  INV_X1 U36558 ( .A(n54049), .ZN(n54040) );
  NAND2_X1 U36559 ( .A1(\DP/ALU0/S_B_MULT[9] ), .A2(\DP/ALU0/S_B_MULT[10] ), 
        .ZN(n54041) );
  NAND2_X1 U36560 ( .A1(n54040), .A2(n54041), .ZN(n54380) );
  INV_X1 U36561 ( .A(n54380), .ZN(n54373) );
  NAND2_X1 U36562 ( .A1(\DP/ALU0/S_B_MULT[11] ), .A2(n54373), .ZN(n54729) );
  AOI22_X1 U36563 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54732), .B1(
        \DP/ALU0/s_A_MULT[14] ), .B2(n54728), .ZN(n54042) );
  OAI21_X1 U36564 ( .B1(n54043), .B2(n54729), .A(n54042), .ZN(n54044) );
  AOI21_X1 U36565 ( .B1(n54856), .B2(n54733), .A(n54044), .ZN(n54696) );
  NOR2_X1 U36566 ( .A1(\intadd_3/n1 ), .A2(n54696), .ZN(n54045) );
  NAND2_X1 U36567 ( .A1(n54697), .A2(n54045), .ZN(n54699) );
  INV_X1 U36568 ( .A(n54046), .ZN(n54048) );
  AOI22_X1 U36569 ( .A1(\DP/ALU0/s_A_MULT[14] ), .A2(n54732), .B1(n54862), 
        .B2(n54733), .ZN(n54047) );
  OAI21_X1 U36570 ( .B1(n54049), .B2(n54048), .A(n54047), .ZN(n54050) );
  AOI21_X1 U36571 ( .B1(\DP/ALU0/s_A_MULT[15] ), .B2(n54728), .A(n54050), .ZN(
        n54703) );
  NAND2_X1 U36572 ( .A1(\intadd_3/n1 ), .A2(n54696), .ZN(n54695) );
  NOR2_X1 U36573 ( .A1(n54697), .A2(n54695), .ZN(n54701) );
  NAND2_X1 U36574 ( .A1(n54703), .A2(n54701), .ZN(n54051) );
  OAI21_X1 U36575 ( .B1(n54699), .B2(n54703), .A(n54051), .ZN(n54052) );
  XNOR2_X1 U36576 ( .A(n54053), .B(n54052), .ZN(n54610) );
  MUX2_X1 U36577 ( .A(n54608), .B(\intadd_2/n1 ), .S(n54610), .Z(n54611) );
  NAND2_X1 U36578 ( .A1(n54108), .A2(n54111), .ZN(n54086) );
  NAND2_X1 U36579 ( .A1(\intadd_1/n1 ), .A2(n54058), .ZN(n54107) );
  NOR2_X1 U36580 ( .A1(n54107), .A2(n54111), .ZN(n54085) );
  NAND2_X1 U36581 ( .A1(n54090), .A2(n54085), .ZN(n54059) );
  OAI21_X1 U36582 ( .B1(n54090), .B2(n54086), .A(n54059), .ZN(n54061) );
  AOI21_X1 U36583 ( .B1(n54062), .B2(n54061), .A(n55300), .ZN(n54060) );
  OAI21_X1 U36584 ( .B1(n54062), .B2(n54061), .A(n54060), .ZN(n54076) );
  OAI211_X1 U36585 ( .C1(n55312), .C2(n54078), .A(n54063), .B(n54076), .ZN(
        \DP/RegALU3/n68 ) );
  INV_X1 U36586 ( .A(n54255), .ZN(n54280) );
  NAND2_X1 U36587 ( .A1(n54064), .A2(n54280), .ZN(n54166) );
  AOI22_X1 U36588 ( .A1(n55175), .A2(\DP/ALU0/s_A_SHIFT[30] ), .B1(n54065), 
        .B2(n54166), .ZN(n54067) );
  AOI22_X1 U36589 ( .A1(n54182), .A2(\DP/ALU0/s_A_SHIFT[7] ), .B1(n53803), 
        .B2(\DP/ALU0/s_A_SHIFT[23] ), .ZN(n54066) );
  NAND2_X1 U36590 ( .A1(n54067), .A2(n54066), .ZN(n54171) );
  AOI22_X1 U36591 ( .A1(n55137), .A2(n54104), .B1(n53807), .B2(n54140), .ZN(
        n54068) );
  OAI21_X1 U36592 ( .B1(n55179), .B2(n54171), .A(n54068), .ZN(n54069) );
  AOI21_X1 U36593 ( .B1(n53804), .B2(n54070), .A(n54069), .ZN(n54097) );
  AOI22_X1 U36594 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[14] ), .B1(n54286), .B2(
        n53710), .ZN(n54074) );
  NAND2_X1 U36595 ( .A1(\DP/ALU0/S_B_LOGIC[30] ), .A2(\DP/ALU0/s_A_LOGIC[30] ), 
        .ZN(n54072) );
  NAND2_X1 U36596 ( .A1(n55187), .A2(n54072), .ZN(n54071) );
  OAI221_X1 U36597 ( .B1(n54072), .B2(n55308), .C1(\DP/ALU0/S_B_LOGIC[30] ), 
        .C2(\DP/ALU0/s_A_LOGIC[30] ), .A(n54071), .ZN(n54073) );
  OAI211_X1 U36598 ( .C1(\intadd_8/SUM[2] ), .C2(n55303), .A(n54074), .B(
        n54073), .ZN(n54075) );
  AOI21_X1 U36599 ( .B1(n55181), .B2(n54097), .A(n54075), .ZN(n54077) );
  OAI211_X1 U36600 ( .C1(n54078), .C2(n55186), .A(n54077), .B(n54076), .ZN(
        \DP/RegALU3/n69 ) );
  AOI22_X1 U36601 ( .A1(n55137), .A2(n54121), .B1(n54079), .B2(n53804), .ZN(
        n54084) );
  INV_X1 U36602 ( .A(n54166), .ZN(n54099) );
  AOI22_X1 U36603 ( .A1(n53802), .A2(\DP/ALU0/s_A_SHIFT[22] ), .B1(n55175), 
        .B2(\DP/ALU0/s_A_SHIFT[29] ), .ZN(n54080) );
  OAI21_X1 U36604 ( .B1(n54081), .B2(n54099), .A(n54080), .ZN(n54082) );
  AOI21_X1 U36605 ( .B1(n54182), .B2(\DP/ALU0/s_A_SHIFT[6] ), .A(n54082), .ZN(
        n54181) );
  NAND2_X1 U36606 ( .A1(n55139), .A2(n54181), .ZN(n54083) );
  OAI211_X1 U36607 ( .C1(n54157), .C2(n53760), .A(n54084), .B(n54083), .ZN(
        n54120) );
  INV_X1 U36608 ( .A(n54085), .ZN(n54087) );
  NAND2_X1 U36609 ( .A1(n54087), .A2(n54086), .ZN(n54089) );
  NOR2_X1 U36610 ( .A1(n54090), .A2(n54089), .ZN(n54088) );
  AOI211_X1 U36611 ( .C1(n54090), .C2(n54089), .A(n55300), .B(n54088), .ZN(
        n54096) );
  AOI22_X1 U36612 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[13] ), .B1(n54286), .B2(
        n7625), .ZN(n54094) );
  NAND2_X1 U36613 ( .A1(\DP/ALU0/S_B_LOGIC[29] ), .A2(\DP/ALU0/s_A_LOGIC[29] ), 
        .ZN(n54092) );
  NAND2_X1 U36614 ( .A1(n55187), .A2(n54092), .ZN(n54091) );
  OAI221_X1 U36615 ( .B1(n54092), .B2(n55308), .C1(\DP/ALU0/S_B_LOGIC[29] ), 
        .C2(\DP/ALU0/s_A_LOGIC[29] ), .A(n54091), .ZN(n54093) );
  OAI211_X1 U36616 ( .C1(\intadd_8/SUM[1] ), .C2(n55303), .A(n54094), .B(
        n54093), .ZN(n54095) );
  AOI211_X1 U36617 ( .C1(n54097), .C2(n55306), .A(n54096), .B(n54095), .ZN(
        n54098) );
  OAI21_X1 U36618 ( .B1(n55312), .B2(n54120), .A(n54098), .ZN(\DP/RegALU3/n70 ) );
  INV_X1 U36619 ( .A(\DP/ALU0/s_A_SHIFT[13] ), .ZN(n54330) );
  AOI21_X1 U36620 ( .B1(n54100), .B2(n54330), .A(n54099), .ZN(n54103) );
  INV_X1 U36621 ( .A(\DP/ALU0/s_A_SHIFT[5] ), .ZN(n54348) );
  INV_X1 U36622 ( .A(n54421), .ZN(n54349) );
  INV_X1 U36623 ( .A(\DP/ALU0/s_A_SHIFT[21] ), .ZN(n54214) );
  OAI22_X1 U36624 ( .A1(n54101), .A2(n54348), .B1(n54349), .B2(n54214), .ZN(
        n54102) );
  AOI211_X1 U36625 ( .C1(n55175), .C2(\DP/ALU0/s_A_SHIFT[28] ), .A(n54103), 
        .B(n54102), .ZN(n54201) );
  AOI22_X1 U36626 ( .A1(n55137), .A2(n54140), .B1(n53804), .B2(n54104), .ZN(
        n54105) );
  OAI21_X1 U36627 ( .B1(n53760), .B2(n54171), .A(n54105), .ZN(n54106) );
  AOI21_X1 U36628 ( .B1(n55139), .B2(n54201), .A(n54106), .ZN(n54132) );
  INV_X1 U36629 ( .A(n54107), .ZN(n54109) );
  NOR2_X1 U36630 ( .A1(n54109), .A2(n54108), .ZN(n54112) );
  NOR2_X1 U36631 ( .A1(n54112), .A2(n54111), .ZN(n54110) );
  AOI211_X1 U36632 ( .C1(n54112), .C2(n54111), .A(n55300), .B(n54110), .ZN(
        n54118) );
  AOI22_X1 U36633 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[12] ), .B1(n54286), .B2(
        n49872), .ZN(n54116) );
  NAND2_X1 U36634 ( .A1(\DP/ALU0/S_B_LOGIC[28] ), .A2(\DP/ALU0/s_A_LOGIC[28] ), 
        .ZN(n54114) );
  NAND2_X1 U36635 ( .A1(n55187), .A2(n54114), .ZN(n54113) );
  OAI221_X1 U36636 ( .B1(n54114), .B2(n55308), .C1(\DP/ALU0/S_B_LOGIC[28] ), 
        .C2(\DP/ALU0/s_A_LOGIC[28] ), .A(n54113), .ZN(n54115) );
  OAI211_X1 U36637 ( .C1(\intadd_8/SUM[0] ), .C2(n55303), .A(n54116), .B(
        n54115), .ZN(n54117) );
  AOI211_X1 U36638 ( .C1(n55181), .C2(n54132), .A(n54118), .B(n54117), .ZN(
        n54119) );
  OAI21_X1 U36639 ( .B1(n55186), .B2(n54120), .A(n54119), .ZN(\DP/RegALU3/n71 ) );
  AOI22_X1 U36640 ( .A1(n53807), .A2(n54181), .B1(n54121), .B2(n53804), .ZN(
        n54127) );
  INV_X1 U36641 ( .A(\DP/ALU0/s_A_SHIFT[20] ), .ZN(n54124) );
  AOI22_X1 U36642 ( .A1(\DP/ALU0/s_A_SHIFT[27] ), .A2(n55175), .B1(n54122), 
        .B2(n54166), .ZN(n54123) );
  OAI21_X1 U36643 ( .B1(n54124), .B2(n54349), .A(n54123), .ZN(n54125) );
  AOI21_X1 U36644 ( .B1(n54182), .B2(\DP/ALU0/s_A_SHIFT[4] ), .A(n54125), .ZN(
        n54212) );
  NAND2_X1 U36645 ( .A1(n55139), .A2(n54212), .ZN(n54126) );
  OAI211_X1 U36646 ( .C1(n54157), .C2(n55177), .A(n54127), .B(n54126), .ZN(
        n54150) );
  AOI22_X1 U36647 ( .A1(n55166), .A2(\intadd_1/SUM[12] ), .B1(n54286), .B2(
        n7623), .ZN(n54130) );
  NOR2_X1 U36648 ( .A1(\DP/ALU0/s_A_LOGIC[27] ), .A2(n55187), .ZN(n54128) );
  AOI22_X1 U36649 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[11] ), .B1(
        \DP/ALU0/S_B_LOGIC[27] ), .B2(n54128), .ZN(n54129) );
  OAI211_X1 U36650 ( .C1(\intadd_0/SUM[26] ), .C2(n55303), .A(n54130), .B(
        n54129), .ZN(n54131) );
  AOI21_X1 U36651 ( .B1(n55306), .B2(n54132), .A(n54131), .ZN(n54135) );
  INV_X1 U36652 ( .A(\DP/ALU0/S_B_LOGIC[27] ), .ZN(n54133) );
  OAI221_X1 U36653 ( .B1(\DP/ALU0/S_B_LOGIC[27] ), .B2(n53809), .C1(n54133), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[27] ), .ZN(n54134) );
  OAI211_X1 U36654 ( .C1(n54150), .C2(n55312), .A(n54135), .B(n54134), .ZN(
        \DP/RegALU3/n72 ) );
  INV_X1 U36655 ( .A(\DP/ALU0/s_A_SHIFT[19] ), .ZN(n54138) );
  AOI22_X1 U36656 ( .A1(\DP/ALU0/s_A_SHIFT[26] ), .A2(n55175), .B1(n54136), 
        .B2(n54166), .ZN(n54137) );
  OAI21_X1 U36657 ( .B1(n54349), .B2(n54138), .A(n54137), .ZN(n54139) );
  AOI21_X1 U36658 ( .B1(n54182), .B2(\DP/ALU0/s_A_SHIFT[3] ), .A(n54139), .ZN(
        n54228) );
  AOI22_X1 U36659 ( .A1(n53807), .A2(n54201), .B1(n53804), .B2(n54140), .ZN(
        n54141) );
  OAI21_X1 U36660 ( .B1(n55177), .B2(n54171), .A(n54141), .ZN(n54142) );
  AOI21_X1 U36661 ( .B1(n55139), .B2(n54228), .A(n54142), .ZN(n54162) );
  AOI22_X1 U36662 ( .A1(n55166), .A2(\intadd_1/SUM[11] ), .B1(n54286), .B2(
        n53648), .ZN(n54145) );
  NOR2_X1 U36663 ( .A1(\DP/ALU0/s_A_LOGIC[26] ), .A2(n55187), .ZN(n54143) );
  AOI22_X1 U36664 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[10] ), .B1(
        \DP/ALU0/S_B_LOGIC[26] ), .B2(n54143), .ZN(n54144) );
  OAI211_X1 U36665 ( .C1(\intadd_0/SUM[25] ), .C2(n55303), .A(n54145), .B(
        n54144), .ZN(n54146) );
  AOI21_X1 U36666 ( .B1(n55181), .B2(n54162), .A(n54146), .ZN(n54149) );
  INV_X1 U36667 ( .A(\DP/ALU0/S_B_LOGIC[26] ), .ZN(n54147) );
  OAI221_X1 U36668 ( .B1(\DP/ALU0/S_B_LOGIC[26] ), .B2(n53809), .C1(n54147), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[26] ), .ZN(n54148) );
  OAI211_X1 U36669 ( .C1(n54150), .C2(n55186), .A(n54149), .B(n54148), .ZN(
        \DP/RegALU3/n73 ) );
  AOI22_X1 U36670 ( .A1(n55137), .A2(n54181), .B1(n53807), .B2(n54212), .ZN(
        n54156) );
  INV_X1 U36671 ( .A(\DP/ALU0/s_A_SHIFT[18] ), .ZN(n54153) );
  AOI22_X1 U36672 ( .A1(\DP/ALU0/s_A_SHIFT[25] ), .A2(n55175), .B1(n54151), 
        .B2(n54166), .ZN(n54152) );
  OAI21_X1 U36673 ( .B1(n54349), .B2(n54153), .A(n54152), .ZN(n54154) );
  AOI21_X1 U36674 ( .B1(n54182), .B2(\DP/ALU0/s_A_SHIFT[2] ), .A(n54154), .ZN(
        n54239) );
  NAND2_X1 U36675 ( .A1(n55139), .A2(n54239), .ZN(n54155) );
  OAI211_X1 U36676 ( .C1(n53761), .C2(n54157), .A(n54156), .B(n54155), .ZN(
        n54180) );
  AOI22_X1 U36677 ( .A1(n55166), .A2(\intadd_1/SUM[10] ), .B1(n54286), .B2(
        n53709), .ZN(n54160) );
  NOR2_X1 U36678 ( .A1(\DP/ALU0/S_B_LOGIC[25] ), .A2(n55187), .ZN(n54158) );
  AOI22_X1 U36679 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[9] ), .B1(
        \DP/ALU0/s_A_LOGIC[25] ), .B2(n54158), .ZN(n54159) );
  OAI211_X1 U36680 ( .C1(\intadd_0/SUM[24] ), .C2(n55303), .A(n54160), .B(
        n54159), .ZN(n54161) );
  AOI21_X1 U36681 ( .B1(n55306), .B2(n54162), .A(n54161), .ZN(n54165) );
  INV_X1 U36682 ( .A(\DP/ALU0/s_A_LOGIC[25] ), .ZN(n54163) );
  OAI221_X1 U36683 ( .B1(\DP/ALU0/s_A_LOGIC[25] ), .B2(n53809), .C1(n54163), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[25] ), .ZN(n54164) );
  OAI211_X1 U36684 ( .C1(n54180), .C2(n55312), .A(n54165), .B(n54164), .ZN(
        \DP/RegALU3/n74 ) );
  INV_X1 U36685 ( .A(\DP/ALU0/s_A_SHIFT[17] ), .ZN(n55140) );
  AOI22_X1 U36686 ( .A1(n55175), .A2(\DP/ALU0/s_A_SHIFT[24] ), .B1(n54167), 
        .B2(n54166), .ZN(n54168) );
  OAI21_X1 U36687 ( .B1(n54349), .B2(n55140), .A(n54168), .ZN(n54169) );
  AOI21_X1 U36688 ( .B1(n54182), .B2(\DP/ALU0/s_A_SHIFT[1] ), .A(n54169), .ZN(
        n54256) );
  AOI22_X1 U36689 ( .A1(n55137), .A2(n54201), .B1(n53807), .B2(n54228), .ZN(
        n54170) );
  OAI21_X1 U36690 ( .B1(n53761), .B2(n54171), .A(n54170), .ZN(n54172) );
  AOI21_X1 U36691 ( .B1(n55139), .B2(n54256), .A(n54172), .ZN(n54194) );
  AOI22_X1 U36692 ( .A1(n55166), .A2(\intadd_1/SUM[9] ), .B1(n54286), .B2(
        n53706), .ZN(n54175) );
  NOR2_X1 U36693 ( .A1(\DP/ALU0/S_B_LOGIC[24] ), .A2(n55187), .ZN(n54173) );
  AOI22_X1 U36694 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[8] ), .B1(
        \DP/ALU0/s_A_LOGIC[24] ), .B2(n54173), .ZN(n54174) );
  OAI211_X1 U36695 ( .C1(\intadd_0/SUM[23] ), .C2(n55303), .A(n54175), .B(
        n54174), .ZN(n54176) );
  AOI21_X1 U36696 ( .B1(n55181), .B2(n54194), .A(n54176), .ZN(n54179) );
  INV_X1 U36697 ( .A(\DP/ALU0/s_A_LOGIC[24] ), .ZN(n54177) );
  OAI221_X1 U36698 ( .B1(\DP/ALU0/s_A_LOGIC[24] ), .B2(n53809), .C1(n54177), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[24] ), .ZN(n54178) );
  OAI211_X1 U36699 ( .C1(n54180), .C2(n55186), .A(n54179), .B(n54178), .ZN(
        \DP/RegALU3/n75 ) );
  AOI22_X1 U36700 ( .A1(n55137), .A2(n54212), .B1(n53804), .B2(n54181), .ZN(
        n54189) );
  AOI22_X1 U36701 ( .A1(n54182), .A2(\DP/ALU0/s_A_SHIFT[0] ), .B1(
        \DP/ALU0/s_A_SHIFT[8] ), .B2(n54300), .ZN(n54186) );
  INV_X1 U36702 ( .A(n54183), .ZN(n54298) );
  NOR2_X1 U36703 ( .A1(n54184), .A2(n54298), .ZN(n55174) );
  AOI22_X1 U36704 ( .A1(\DP/ALU0/s_A_SHIFT[31] ), .A2(n55174), .B1(n55175), 
        .B2(\DP/ALU0/s_A_SHIFT[23] ), .ZN(n54185) );
  NAND2_X1 U36705 ( .A1(n54186), .A2(n54185), .ZN(n54187) );
  AOI211_X1 U36706 ( .C1(\DP/ALU0/s_A_SHIFT[16] ), .C2(n53802), .A(n54255), 
        .B(n54187), .ZN(n54267) );
  AOI22_X1 U36707 ( .A1(n53807), .A2(n54239), .B1(n55139), .B2(n54267), .ZN(
        n54188) );
  NAND2_X1 U36708 ( .A1(n54189), .A2(n54188), .ZN(n54211) );
  AOI22_X1 U36709 ( .A1(n55166), .A2(\intadd_1/SUM[8] ), .B1(n54286), .B2(
        n7661), .ZN(n54192) );
  NOR2_X1 U36710 ( .A1(\DP/ALU0/S_B_LOGIC[23] ), .A2(n55187), .ZN(n54190) );
  AOI22_X1 U36711 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[7] ), .B1(
        \DP/ALU0/s_A_LOGIC[23] ), .B2(n54190), .ZN(n54191) );
  OAI211_X1 U36712 ( .C1(\intadd_0/SUM[22] ), .C2(n55303), .A(n54192), .B(
        n54191), .ZN(n54193) );
  AOI21_X1 U36713 ( .B1(n55306), .B2(n54194), .A(n54193), .ZN(n54197) );
  INV_X1 U36714 ( .A(\DP/ALU0/s_A_LOGIC[23] ), .ZN(n54195) );
  OAI221_X1 U36715 ( .B1(\DP/ALU0/s_A_LOGIC[23] ), .B2(n53809), .C1(n54195), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[23] ), .ZN(n54196) );
  OAI211_X1 U36716 ( .C1(n54211), .C2(n55312), .A(n54197), .B(n54196), .ZN(
        \DP/RegALU3/n76 ) );
  INV_X1 U36717 ( .A(\DP/ALU0/s_A_SHIFT[22] ), .ZN(n54200) );
  AOI21_X1 U36718 ( .B1(n53802), .B2(\DP/ALU0/s_A_SHIFT[15] ), .A(n54255), 
        .ZN(n54199) );
  AOI22_X1 U36719 ( .A1(\DP/ALU0/s_A_SHIFT[30] ), .A2(n53808), .B1(n54300), 
        .B2(\DP/ALU0/s_A_SHIFT[7] ), .ZN(n54198) );
  OAI211_X1 U36720 ( .C1(n54411), .C2(n54200), .A(n54199), .B(n54198), .ZN(
        n54284) );
  AOI22_X1 U36721 ( .A1(n55137), .A2(n54228), .B1(n53804), .B2(n54201), .ZN(
        n54202) );
  OAI21_X1 U36722 ( .B1(n55179), .B2(n54284), .A(n54202), .ZN(n54203) );
  AOI21_X1 U36723 ( .B1(n53807), .B2(n54256), .A(n54203), .ZN(n54222) );
  AOI22_X1 U36724 ( .A1(n55166), .A2(\intadd_1/SUM[7] ), .B1(n54286), .B2(
        n7622), .ZN(n54206) );
  NOR2_X1 U36725 ( .A1(\DP/ALU0/S_B_LOGIC[22] ), .A2(n55187), .ZN(n54204) );
  AOI22_X1 U36726 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[6] ), .B1(
        \DP/ALU0/s_A_LOGIC[22] ), .B2(n54204), .ZN(n54205) );
  OAI211_X1 U36727 ( .C1(\intadd_0/SUM[21] ), .C2(n55303), .A(n54206), .B(
        n54205), .ZN(n54207) );
  AOI21_X1 U36728 ( .B1(n55181), .B2(n54222), .A(n54207), .ZN(n54210) );
  INV_X1 U36729 ( .A(\DP/ALU0/s_A_LOGIC[22] ), .ZN(n54208) );
  OAI221_X1 U36730 ( .B1(\DP/ALU0/s_A_LOGIC[22] ), .B2(n53809), .C1(n54208), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[22] ), .ZN(n54209) );
  OAI211_X1 U36731 ( .C1(n54211), .C2(n55186), .A(n54210), .B(n54209), .ZN(
        \DP/RegALU3/n77 ) );
  AOI22_X1 U36732 ( .A1(n55137), .A2(n54239), .B1(n53804), .B2(n54212), .ZN(
        n54217) );
  AOI22_X1 U36733 ( .A1(n54300), .A2(\DP/ALU0/s_A_SHIFT[6] ), .B1(
        \DP/ALU0/s_A_SHIFT[29] ), .B2(n55174), .ZN(n54213) );
  OAI21_X1 U36734 ( .B1(n54411), .B2(n54214), .A(n54213), .ZN(n54215) );
  AOI211_X1 U36735 ( .C1(n54421), .C2(\DP/ALU0/s_A_SHIFT[14] ), .A(n54255), 
        .B(n54215), .ZN(n54304) );
  AOI22_X1 U36736 ( .A1(n53807), .A2(n54267), .B1(n55139), .B2(n54304), .ZN(
        n54216) );
  NAND2_X1 U36737 ( .A1(n54217), .A2(n54216), .ZN(n54238) );
  AOI22_X1 U36738 ( .A1(n55166), .A2(\intadd_1/SUM[6] ), .B1(n54286), .B2(
        n7660), .ZN(n54220) );
  NOR2_X1 U36739 ( .A1(\DP/ALU0/S_B_LOGIC[21] ), .A2(n55187), .ZN(n54218) );
  AOI22_X1 U36740 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[5] ), .B1(
        \DP/ALU0/s_A_LOGIC[21] ), .B2(n54218), .ZN(n54219) );
  OAI211_X1 U36741 ( .C1(\intadd_0/SUM[20] ), .C2(n55303), .A(n54220), .B(
        n54219), .ZN(n54221) );
  AOI21_X1 U36742 ( .B1(n55306), .B2(n54222), .A(n54221), .ZN(n54225) );
  INV_X1 U36743 ( .A(\DP/ALU0/s_A_LOGIC[21] ), .ZN(n54223) );
  OAI221_X1 U36744 ( .B1(\DP/ALU0/s_A_LOGIC[21] ), .B2(n53809), .C1(n54223), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[21] ), .ZN(n54224) );
  OAI211_X1 U36745 ( .C1(n55312), .C2(n54238), .A(n54225), .B(n54224), .ZN(
        \DP/RegALU3/n78 ) );
  AOI22_X1 U36746 ( .A1(\DP/ALU0/s_A_SHIFT[20] ), .A2(n55175), .B1(n54300), 
        .B2(\DP/ALU0/s_A_SHIFT[5] ), .ZN(n54226) );
  OAI211_X1 U36747 ( .C1(n54349), .C2(n54330), .A(n54226), .B(n54280), .ZN(
        n54227) );
  AOI21_X1 U36748 ( .B1(\DP/ALU0/s_A_SHIFT[28] ), .B2(n55174), .A(n54227), 
        .ZN(n54320) );
  AOI22_X1 U36749 ( .A1(n55137), .A2(n54256), .B1(n53804), .B2(n54228), .ZN(
        n54229) );
  OAI21_X1 U36750 ( .B1(n53760), .B2(n54284), .A(n54229), .ZN(n54230) );
  AOI21_X1 U36751 ( .B1(n55139), .B2(n54320), .A(n54230), .ZN(n54249) );
  AOI22_X1 U36752 ( .A1(n55166), .A2(\intadd_1/SUM[5] ), .B1(n54286), .B2(
        n7621), .ZN(n54233) );
  NOR2_X1 U36753 ( .A1(\DP/ALU0/S_B_LOGIC[20] ), .A2(n55187), .ZN(n54231) );
  AOI22_X1 U36754 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[4] ), .B1(
        \DP/ALU0/s_A_LOGIC[20] ), .B2(n54231), .ZN(n54232) );
  OAI211_X1 U36755 ( .C1(\intadd_0/SUM[19] ), .C2(n55303), .A(n54233), .B(
        n54232), .ZN(n54234) );
  AOI21_X1 U36756 ( .B1(n55181), .B2(n54249), .A(n54234), .ZN(n54237) );
  INV_X1 U36757 ( .A(\DP/ALU0/s_A_LOGIC[20] ), .ZN(n54235) );
  OAI221_X1 U36758 ( .B1(\DP/ALU0/s_A_LOGIC[20] ), .B2(n53809), .C1(n54235), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[20] ), .ZN(n54236) );
  OAI211_X1 U36759 ( .C1(n54238), .C2(n55186), .A(n54237), .B(n54236), .ZN(
        \DP/RegALU3/n79 ) );
  AOI22_X1 U36760 ( .A1(n55137), .A2(n54267), .B1(n53804), .B2(n54239), .ZN(
        n54244) );
  AOI22_X1 U36761 ( .A1(n55175), .A2(\DP/ALU0/s_A_SHIFT[19] ), .B1(n54300), 
        .B2(\DP/ALU0/s_A_SHIFT[4] ), .ZN(n54240) );
  OAI211_X1 U36762 ( .C1(n54349), .C2(n54241), .A(n54240), .B(n54280), .ZN(
        n54242) );
  AOI21_X1 U36763 ( .B1(\DP/ALU0/s_A_SHIFT[27] ), .B2(n53808), .A(n54242), 
        .ZN(n54328) );
  AOI22_X1 U36764 ( .A1(n53807), .A2(n54304), .B1(n55139), .B2(n54328), .ZN(
        n54243) );
  NAND2_X1 U36765 ( .A1(n54244), .A2(n54243), .ZN(n54266) );
  AOI22_X1 U36766 ( .A1(n55166), .A2(\intadd_1/SUM[4] ), .B1(n54286), .B2(
        n53708), .ZN(n54247) );
  NOR2_X1 U36767 ( .A1(\DP/ALU0/S_B_LOGIC[19] ), .A2(n55187), .ZN(n54245) );
  AOI22_X1 U36768 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[3] ), .B1(
        \DP/ALU0/s_A_LOGIC[19] ), .B2(n54245), .ZN(n54246) );
  OAI211_X1 U36769 ( .C1(\intadd_0/SUM[18] ), .C2(n55303), .A(n54247), .B(
        n54246), .ZN(n54248) );
  AOI21_X1 U36770 ( .B1(n55306), .B2(n54249), .A(n54248), .ZN(n54252) );
  INV_X1 U36771 ( .A(\DP/ALU0/s_A_LOGIC[19] ), .ZN(n54250) );
  OAI221_X1 U36772 ( .B1(\DP/ALU0/s_A_LOGIC[19] ), .B2(n53809), .C1(n54250), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[19] ), .ZN(n54251) );
  OAI211_X1 U36773 ( .C1(n55312), .C2(n54266), .A(n54252), .B(n54251), .ZN(
        \DP/RegALU3/n80 ) );
  AOI22_X1 U36774 ( .A1(\DP/ALU0/s_A_SHIFT[18] ), .A2(n55175), .B1(
        \DP/ALU0/s_A_SHIFT[26] ), .B2(n55174), .ZN(n54253) );
  OAI21_X1 U36775 ( .B1(n54349), .B2(n54362), .A(n54253), .ZN(n54254) );
  AOI211_X1 U36776 ( .C1(n54300), .C2(\DP/ALU0/s_A_SHIFT[3] ), .A(n54255), .B(
        n54254), .ZN(n54351) );
  AOI22_X1 U36777 ( .A1(n53807), .A2(n54320), .B1(n53804), .B2(n54256), .ZN(
        n54257) );
  OAI21_X1 U36778 ( .B1(n55177), .B2(n54284), .A(n54257), .ZN(n54258) );
  AOI21_X1 U36779 ( .B1(n55139), .B2(n54351), .A(n54258), .ZN(n54276) );
  AOI22_X1 U36780 ( .A1(n55166), .A2(\intadd_1/SUM[3] ), .B1(n54286), .B2(
        n7663), .ZN(n54261) );
  NOR2_X1 U36781 ( .A1(\DP/ALU0/s_A_LOGIC[18] ), .A2(n55187), .ZN(n54259) );
  AOI22_X1 U36782 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[2] ), .B1(
        \DP/ALU0/S_B_LOGIC[18] ), .B2(n54259), .ZN(n54260) );
  OAI211_X1 U36783 ( .C1(\intadd_0/SUM[17] ), .C2(n55303), .A(n54261), .B(
        n54260), .ZN(n54262) );
  AOI21_X1 U36784 ( .B1(n55181), .B2(n54276), .A(n54262), .ZN(n54265) );
  INV_X1 U36785 ( .A(\DP/ALU0/S_B_LOGIC[18] ), .ZN(n54263) );
  OAI221_X1 U36786 ( .B1(\DP/ALU0/S_B_LOGIC[18] ), .B2(n53809), .C1(n54263), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[18] ), .ZN(n54264) );
  OAI211_X1 U36787 ( .C1(n54266), .C2(n55186), .A(n54265), .B(n54264), .ZN(
        \DP/RegALU3/n81 ) );
  AOI22_X1 U36788 ( .A1(n55137), .A2(n54304), .B1(n53804), .B2(n54267), .ZN(
        n54271) );
  AOI22_X1 U36789 ( .A1(n55175), .A2(\DP/ALU0/s_A_SHIFT[17] ), .B1(n54300), 
        .B2(\DP/ALU0/s_A_SHIFT[2] ), .ZN(n54268) );
  OAI211_X1 U36790 ( .C1(n54375), .C2(n54349), .A(n54268), .B(n54280), .ZN(
        n54269) );
  AOI21_X1 U36791 ( .B1(\DP/ALU0/s_A_SHIFT[25] ), .B2(n53808), .A(n54269), 
        .ZN(n54360) );
  AOI22_X1 U36792 ( .A1(n53807), .A2(n54328), .B1(n55139), .B2(n54360), .ZN(
        n54270) );
  NAND2_X1 U36793 ( .A1(n54271), .A2(n54270), .ZN(n54295) );
  AOI22_X1 U36794 ( .A1(n55166), .A2(\intadd_1/SUM[2] ), .B1(n54286), .B2(
        n53707), .ZN(n54274) );
  NOR2_X1 U36795 ( .A1(\DP/ALU0/s_A_LOGIC[17] ), .A2(n55187), .ZN(n54272) );
  AOI22_X1 U36796 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[1] ), .B1(
        \DP/ALU0/S_B_LOGIC[17] ), .B2(n54272), .ZN(n54273) );
  OAI211_X1 U36797 ( .C1(\intadd_0/SUM[16] ), .C2(n55303), .A(n54274), .B(
        n54273), .ZN(n54275) );
  AOI21_X1 U36798 ( .B1(n55306), .B2(n54276), .A(n54275), .ZN(n54279) );
  INV_X1 U36799 ( .A(\DP/ALU0/S_B_LOGIC[17] ), .ZN(n54277) );
  OAI221_X1 U36800 ( .B1(\DP/ALU0/S_B_LOGIC[17] ), .B2(n53809), .C1(n54277), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[17] ), .ZN(n54278) );
  OAI211_X1 U36801 ( .C1(n55312), .C2(n54295), .A(n54279), .B(n54278), .ZN(
        \DP/RegALU3/n82 ) );
  AOI22_X1 U36802 ( .A1(\DP/ALU0/s_A_SHIFT[16] ), .A2(n55175), .B1(n54300), 
        .B2(\DP/ALU0/s_A_SHIFT[1] ), .ZN(n54281) );
  OAI211_X1 U36803 ( .C1(n54349), .C2(n54393), .A(n54281), .B(n54280), .ZN(
        n54282) );
  AOI21_X1 U36804 ( .B1(\DP/ALU0/s_A_SHIFT[24] ), .B2(n55174), .A(n54282), 
        .ZN(n54377) );
  AOI22_X1 U36805 ( .A1(n55137), .A2(n54320), .B1(n53807), .B2(n54351), .ZN(
        n54283) );
  OAI21_X1 U36806 ( .B1(n53761), .B2(n54284), .A(n54283), .ZN(n54285) );
  AOI21_X1 U36807 ( .B1(n55139), .B2(n54377), .A(n54285), .ZN(n54307) );
  AOI22_X1 U36808 ( .A1(n55166), .A2(\intadd_1/SUM[1] ), .B1(n54286), .B2(
        n7662), .ZN(n54290) );
  NOR2_X1 U36809 ( .A1(\DP/ALU0/s_A_LOGIC[16] ), .A2(n55187), .ZN(n54287) );
  AOI22_X1 U36810 ( .A1(n54288), .A2(\DP/ALU0/S_B_LHI[0] ), .B1(
        \DP/ALU0/S_B_LOGIC[16] ), .B2(n54287), .ZN(n54289) );
  OAI211_X1 U36811 ( .C1(\intadd_0/SUM[15] ), .C2(n55303), .A(n54290), .B(
        n54289), .ZN(n54291) );
  AOI21_X1 U36812 ( .B1(n55181), .B2(n54307), .A(n54291), .ZN(n54294) );
  INV_X1 U36813 ( .A(\DP/ALU0/S_B_LOGIC[16] ), .ZN(n54292) );
  OAI221_X1 U36814 ( .B1(\DP/ALU0/S_B_LOGIC[16] ), .B2(n53809), .C1(n54292), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[16] ), .ZN(n54293) );
  OAI211_X1 U36815 ( .C1(n54295), .C2(n55186), .A(n54294), .B(n54293), .ZN(
        \DP/RegALU3/n83 ) );
  INV_X1 U36816 ( .A(\DP/ALU0/s_A_LOGIC[15] ), .ZN(n54308) );
  NOR3_X1 U36817 ( .A1(\DP/ALU0/S_B_LOGIC[15] ), .A2(n54308), .A3(n55187), 
        .ZN(n54297) );
  OAI22_X1 U36818 ( .A1(n49809), .A2(n5463), .B1(\intadd_0/SUM[14] ), .B2(
        n55303), .ZN(n54296) );
  AOI211_X1 U36819 ( .C1(n55166), .C2(\intadd_1/SUM[0] ), .A(n54297), .B(
        n54296), .ZN(n54311) );
  INV_X1 U36820 ( .A(n55176), .ZN(n55141) );
  AOI22_X1 U36821 ( .A1(n53803), .A2(\DP/ALU0/s_A_SHIFT[8] ), .B1(n54300), 
        .B2(\DP/ALU0/s_A_SHIFT[0] ), .ZN(n54302) );
  AOI22_X1 U36822 ( .A1(n55175), .A2(\DP/ALU0/s_A_SHIFT[15] ), .B1(
        \DP/ALU0/s_A_SHIFT[23] ), .B2(n55174), .ZN(n54301) );
  OAI211_X1 U36823 ( .C1(n54303), .C2(n55141), .A(n54302), .B(n54301), .ZN(
        n54396) );
  AOI22_X1 U36824 ( .A1(n55137), .A2(n54328), .B1(n53804), .B2(n54304), .ZN(
        n54305) );
  OAI21_X1 U36825 ( .B1(n55179), .B2(n54396), .A(n54305), .ZN(n54306) );
  AOI21_X1 U36826 ( .B1(n53807), .B2(n54360), .A(n54306), .ZN(n54323) );
  AOI22_X1 U36827 ( .A1(n55181), .A2(n54323), .B1(n55306), .B2(n54307), .ZN(
        n54310) );
  OAI221_X1 U36828 ( .B1(\DP/ALU0/s_A_LOGIC[15] ), .B2(n53809), .C1(n54308), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[15] ), .ZN(n54309) );
  NAND3_X1 U36829 ( .A1(n54311), .A2(n54310), .A3(n54309), .ZN(
        \DP/RegALU3/n84 ) );
  INV_X1 U36830 ( .A(\DP/ALU0/s_A_MULT[0] ), .ZN(n55299) );
  NOR3_X1 U36831 ( .A1(\intadd_2/SUM[1] ), .A2(n54312), .A3(n55299), .ZN(
        \intadd_1/A[0] ) );
  NOR2_X1 U36832 ( .A1(\DP/ALU0/s_A_LOGIC[14] ), .A2(n55187), .ZN(n54317) );
  NAND2_X1 U36833 ( .A1(\DP/ALU0/s_A_MULT[0] ), .A2(n54313), .ZN(n54314) );
  AOI211_X1 U36834 ( .C1(\intadd_2/SUM[1] ), .C2(n54314), .A(\intadd_1/A[0] ), 
        .B(n55300), .ZN(n54316) );
  OAI22_X1 U36835 ( .A1(\intadd_0/SUM[13] ), .A2(n55303), .B1(n5463), .B2(
        n53660), .ZN(n54315) );
  AOI211_X1 U36836 ( .C1(n54317), .C2(\DP/ALU0/S_B_LOGIC[14] ), .A(n54316), 
        .B(n54315), .ZN(n54327) );
  AOI22_X1 U36837 ( .A1(n55175), .A2(\DP/ALU0/s_A_SHIFT[14] ), .B1(
        \DP/ALU0/s_A_SHIFT[30] ), .B2(n55176), .ZN(n54319) );
  AOI22_X1 U36838 ( .A1(n53802), .A2(\DP/ALU0/s_A_SHIFT[7] ), .B1(
        \DP/ALU0/s_A_SHIFT[22] ), .B2(n53808), .ZN(n54318) );
  NAND2_X1 U36839 ( .A1(n54319), .A2(n54318), .ZN(n54414) );
  AOI22_X1 U36840 ( .A1(n55137), .A2(n54351), .B1(n53804), .B2(n54320), .ZN(
        n54321) );
  OAI21_X1 U36841 ( .B1(n55179), .B2(n54414), .A(n54321), .ZN(n54322) );
  AOI21_X1 U36842 ( .B1(n53807), .B2(n54377), .A(n54322), .ZN(n54337) );
  AOI22_X1 U36843 ( .A1(n55181), .A2(n54337), .B1(n55306), .B2(n54323), .ZN(
        n54326) );
  INV_X1 U36844 ( .A(\DP/ALU0/S_B_LOGIC[14] ), .ZN(n54324) );
  OAI221_X1 U36845 ( .B1(\DP/ALU0/S_B_LOGIC[14] ), .B2(n53809), .C1(n54324), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[14] ), .ZN(n54325) );
  NAND3_X1 U36846 ( .A1(n54327), .A2(n54326), .A3(n54325), .ZN(
        \DP/RegALU3/n85 ) );
  AOI22_X1 U36847 ( .A1(n55137), .A2(n54360), .B1(n53804), .B2(n54328), .ZN(
        n54333) );
  AOI22_X1 U36848 ( .A1(n53803), .A2(\DP/ALU0/s_A_SHIFT[6] ), .B1(
        \DP/ALU0/s_A_SHIFT[29] ), .B2(n55176), .ZN(n54329) );
  OAI21_X1 U36849 ( .B1(n54411), .B2(n54330), .A(n54329), .ZN(n54331) );
  AOI21_X1 U36850 ( .B1(\DP/ALU0/s_A_SHIFT[21] ), .B2(n55174), .A(n54331), 
        .ZN(n54424) );
  NAND2_X1 U36851 ( .A1(n55139), .A2(n54424), .ZN(n54332) );
  OAI211_X1 U36852 ( .C1(n54396), .C2(n53760), .A(n54333), .B(n54332), .ZN(
        n54359) );
  OAI22_X1 U36853 ( .A1(n49810), .A2(n5463), .B1(\intadd_2/SUM[0] ), .B2(
        n55300), .ZN(n54336) );
  NAND2_X1 U36854 ( .A1(n53809), .A2(\DP/ALU0/S_B_LOGIC[13] ), .ZN(n54334) );
  OAI22_X1 U36855 ( .A1(\intadd_0/SUM[12] ), .A2(n55303), .B1(
        \DP/ALU0/s_A_LOGIC[13] ), .B2(n54334), .ZN(n54335) );
  AOI211_X1 U36856 ( .C1(n55306), .C2(n54337), .A(n54336), .B(n54335), .ZN(
        n54340) );
  INV_X1 U36857 ( .A(\DP/ALU0/S_B_LOGIC[13] ), .ZN(n54338) );
  OAI221_X1 U36858 ( .B1(\DP/ALU0/S_B_LOGIC[13] ), .B2(n53809), .C1(n54338), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[13] ), .ZN(n54339) );
  OAI211_X1 U36859 ( .C1(n54359), .C2(n55312), .A(n54340), .B(n54339), .ZN(
        \DP/RegALU3/n86 ) );
  INV_X1 U36860 ( .A(\intadd_3/SUM[1] ), .ZN(n54341) );
  NAND3_X1 U36861 ( .A1(n54341), .A2(n54342), .A3(\DP/ALU0/s_A_MULT[0] ), .ZN(
        \intadd_2/A[0] ) );
  NAND2_X1 U36862 ( .A1(\DP/ALU0/s_A_MULT[0] ), .A2(n54342), .ZN(n54343) );
  AOI21_X1 U36863 ( .B1(\intadd_3/SUM[1] ), .B2(n54343), .A(n55300), .ZN(
        n54346) );
  INV_X1 U36864 ( .A(\DP/ALU0/S_B_LOGIC[12] ), .ZN(n54354) );
  NOR3_X1 U36865 ( .A1(\DP/ALU0/s_A_LOGIC[12] ), .A2(n54354), .A3(n55187), 
        .ZN(n54345) );
  OAI22_X1 U36866 ( .A1(n49814), .A2(n5463), .B1(\intadd_0/SUM[11] ), .B2(
        n55303), .ZN(n54344) );
  AOI211_X1 U36867 ( .C1(n54346), .C2(\intadd_2/A[0] ), .A(n54345), .B(n54344), 
        .ZN(n54358) );
  AOI22_X1 U36868 ( .A1(\DP/ALU0/s_A_SHIFT[20] ), .A2(n55174), .B1(
        \DP/ALU0/s_A_SHIFT[12] ), .B2(n55175), .ZN(n54347) );
  OAI21_X1 U36869 ( .B1(n54349), .B2(n54348), .A(n54347), .ZN(n54350) );
  AOI21_X1 U36870 ( .B1(\DP/ALU0/s_A_SHIFT[28] ), .B2(n55176), .A(n54350), 
        .ZN(n54434) );
  AOI22_X1 U36871 ( .A1(n55137), .A2(n54377), .B1(n53804), .B2(n54351), .ZN(
        n54352) );
  OAI21_X1 U36872 ( .B1(n53760), .B2(n54414), .A(n54352), .ZN(n54353) );
  AOI21_X1 U36873 ( .B1(n55139), .B2(n54434), .A(n54353), .ZN(n54369) );
  AOI22_X1 U36874 ( .A1(\DP/ALU0/S_B_LOGIC[12] ), .A2(n54355), .B1(n55187), 
        .B2(n54354), .ZN(n54356) );
  AOI22_X1 U36875 ( .A1(n55181), .A2(n54369), .B1(\DP/ALU0/s_A_LOGIC[12] ), 
        .B2(n54356), .ZN(n54357) );
  OAI211_X1 U36876 ( .C1(n55186), .C2(n54359), .A(n54358), .B(n54357), .ZN(
        \DP/RegALU3/n87 ) );
  AOI22_X1 U36877 ( .A1(n53807), .A2(n54424), .B1(n53804), .B2(n54360), .ZN(
        n54365) );
  AOI22_X1 U36878 ( .A1(n54421), .A2(\DP/ALU0/s_A_SHIFT[4] ), .B1(
        \DP/ALU0/s_A_SHIFT[27] ), .B2(n55176), .ZN(n54361) );
  OAI21_X1 U36879 ( .B1(n54411), .B2(n54362), .A(n54361), .ZN(n54363) );
  AOI21_X1 U36880 ( .B1(\DP/ALU0/s_A_SHIFT[19] ), .B2(n53808), .A(n54363), 
        .ZN(n54449) );
  NAND2_X1 U36881 ( .A1(n55139), .A2(n54449), .ZN(n54364) );
  OAI211_X1 U36882 ( .C1(n54396), .C2(n55177), .A(n54365), .B(n54364), .ZN(
        n54389) );
  OAI22_X1 U36883 ( .A1(n49843), .A2(n5463), .B1(\intadd_3/SUM[0] ), .B2(
        n55300), .ZN(n54368) );
  NAND2_X1 U36884 ( .A1(n53809), .A2(\DP/ALU0/s_A_LOGIC[11] ), .ZN(n54366) );
  OAI22_X1 U36885 ( .A1(\intadd_0/SUM[10] ), .A2(n55303), .B1(
        \DP/ALU0/S_B_LOGIC[11] ), .B2(n54366), .ZN(n54367) );
  AOI211_X1 U36886 ( .C1(n55306), .C2(n54369), .A(n54368), .B(n54367), .ZN(
        n54372) );
  INV_X1 U36887 ( .A(\DP/ALU0/s_A_LOGIC[11] ), .ZN(n54370) );
  OAI221_X1 U36888 ( .B1(\DP/ALU0/s_A_LOGIC[11] ), .B2(n53809), .C1(n54370), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[11] ), .ZN(n54371) );
  OAI211_X1 U36889 ( .C1(n54389), .C2(n55312), .A(n54372), .B(n54371), .ZN(
        \DP/RegALU3/n88 ) );
  NAND3_X1 U36890 ( .A1(\DP/ALU0/s_A_MULT[0] ), .A2(n54373), .A3(
        \intadd_4/SUM[1] ), .ZN(\intadd_3/A[0] ) );
  AOI22_X1 U36891 ( .A1(n53803), .A2(\DP/ALU0/s_A_SHIFT[3] ), .B1(
        \DP/ALU0/s_A_SHIFT[26] ), .B2(n55176), .ZN(n54374) );
  OAI21_X1 U36892 ( .B1(n54375), .B2(n54411), .A(n54374), .ZN(n54376) );
  AOI21_X1 U36893 ( .B1(\DP/ALU0/s_A_SHIFT[18] ), .B2(n53808), .A(n54376), 
        .ZN(n54457) );
  AOI22_X1 U36894 ( .A1(n53807), .A2(n54434), .B1(n53804), .B2(n54377), .ZN(
        n54378) );
  OAI21_X1 U36895 ( .B1(n55177), .B2(n54414), .A(n54378), .ZN(n54379) );
  AOI21_X1 U36896 ( .B1(n55139), .B2(n54457), .A(n54379), .ZN(n54398) );
  OAI22_X1 U36897 ( .A1(n49808), .A2(n5463), .B1(\intadd_0/SUM[9] ), .B2(
        n55303), .ZN(n54385) );
  NAND2_X1 U36898 ( .A1(n53809), .A2(\DP/ALU0/S_B_LOGIC[10] ), .ZN(n54383) );
  NOR2_X1 U36899 ( .A1(n55299), .A2(n54380), .ZN(n54381) );
  OAI211_X1 U36900 ( .C1(n54381), .C2(\intadd_4/SUM[1] ), .A(n55166), .B(
        \intadd_3/A[0] ), .ZN(n54382) );
  OAI21_X1 U36901 ( .B1(\DP/ALU0/s_A_LOGIC[10] ), .B2(n54383), .A(n54382), 
        .ZN(n54384) );
  AOI211_X1 U36902 ( .C1(n55181), .C2(n54398), .A(n54385), .B(n54384), .ZN(
        n54388) );
  INV_X1 U36903 ( .A(\DP/ALU0/S_B_LOGIC[10] ), .ZN(n54386) );
  OAI221_X1 U36904 ( .B1(\DP/ALU0/S_B_LOGIC[10] ), .B2(n53809), .C1(n54386), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[10] ), .ZN(n54387) );
  OAI211_X1 U36905 ( .C1(n54389), .C2(n55186), .A(n54388), .B(n54387), .ZN(
        \DP/RegALU3/n89 ) );
  INV_X1 U36906 ( .A(\DP/ALU0/s_A_LOGIC[9] ), .ZN(n54399) );
  NOR3_X1 U36907 ( .A1(\DP/ALU0/S_B_LOGIC[9] ), .A2(n54399), .A3(n55187), .ZN(
        n54391) );
  OAI22_X1 U36908 ( .A1(n49832), .A2(n5463), .B1(\intadd_0/SUM[8] ), .B2(
        n55303), .ZN(n54390) );
  AOI211_X1 U36909 ( .C1(n55166), .C2(\intadd_4/SUM[0] ), .A(n54391), .B(
        n54390), .ZN(n54402) );
  AOI22_X1 U36910 ( .A1(n54421), .A2(\DP/ALU0/s_A_SHIFT[2] ), .B1(
        \DP/ALU0/s_A_SHIFT[17] ), .B2(n53808), .ZN(n54392) );
  OAI21_X1 U36911 ( .B1(n54411), .B2(n54393), .A(n54392), .ZN(n54394) );
  AOI21_X1 U36912 ( .B1(\DP/ALU0/s_A_SHIFT[25] ), .B2(n55176), .A(n54394), 
        .ZN(n54461) );
  AOI22_X1 U36913 ( .A1(n55137), .A2(n54424), .B1(n53807), .B2(n54449), .ZN(
        n54395) );
  OAI21_X1 U36914 ( .B1(n53761), .B2(n54396), .A(n54395), .ZN(n54397) );
  AOI21_X1 U36915 ( .B1(n55139), .B2(n54461), .A(n54397), .ZN(n54416) );
  AOI22_X1 U36916 ( .A1(n55181), .A2(n54416), .B1(n55306), .B2(n54398), .ZN(
        n54401) );
  OAI221_X1 U36917 ( .B1(\DP/ALU0/s_A_LOGIC[9] ), .B2(n53809), .C1(n54399), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[9] ), .ZN(n54400) );
  NAND3_X1 U36918 ( .A1(n54402), .A2(n54401), .A3(n54400), .ZN(
        \DP/RegALU3/n90 ) );
  NOR3_X1 U36919 ( .A1(\intadd_5/SUM[1] ), .A2(n54403), .A3(n55299), .ZN(
        \intadd_4/A[0] ) );
  NOR2_X1 U36920 ( .A1(\DP/ALU0/s_A_LOGIC[8] ), .A2(n55187), .ZN(n54408) );
  NAND2_X1 U36921 ( .A1(\DP/ALU0/s_A_MULT[0] ), .A2(n54404), .ZN(n54405) );
  AOI211_X1 U36922 ( .C1(\intadd_5/SUM[1] ), .C2(n54405), .A(\intadd_4/A[0] ), 
        .B(n55300), .ZN(n54407) );
  OAI22_X1 U36923 ( .A1(\intadd_0/SUM[7] ), .A2(n55303), .B1(n5463), .B2(
        n53661), .ZN(n54406) );
  AOI211_X1 U36924 ( .C1(n54408), .C2(\DP/ALU0/S_B_LOGIC[8] ), .A(n54407), .B(
        n54406), .ZN(n54420) );
  INV_X1 U36925 ( .A(\DP/ALU0/s_A_SHIFT[8] ), .ZN(n54410) );
  AOI22_X1 U36926 ( .A1(n53802), .A2(\DP/ALU0/s_A_SHIFT[1] ), .B1(
        \DP/ALU0/s_A_SHIFT[16] ), .B2(n53808), .ZN(n54409) );
  OAI21_X1 U36927 ( .B1(n54411), .B2(n54410), .A(n54409), .ZN(n54412) );
  AOI21_X1 U36928 ( .B1(\DP/ALU0/s_A_SHIFT[24] ), .B2(n55176), .A(n54412), 
        .ZN(n54458) );
  AOI22_X1 U36929 ( .A1(n55137), .A2(n54434), .B1(n53807), .B2(n54457), .ZN(
        n54413) );
  OAI21_X1 U36930 ( .B1(n53761), .B2(n54414), .A(n54413), .ZN(n54415) );
  AOI21_X1 U36931 ( .B1(n55139), .B2(n54458), .A(n54415), .ZN(n54430) );
  AOI22_X1 U36932 ( .A1(n55181), .A2(n54430), .B1(n55306), .B2(n54416), .ZN(
        n54419) );
  INV_X1 U36933 ( .A(\DP/ALU0/S_B_LOGIC[8] ), .ZN(n54417) );
  OAI221_X1 U36934 ( .B1(\DP/ALU0/S_B_LOGIC[8] ), .B2(n53809), .C1(n54417), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[8] ), .ZN(n54418) );
  NAND3_X1 U36935 ( .A1(n54420), .A2(n54419), .A3(n54418), .ZN(
        \DP/RegALU3/n91 ) );
  AOI22_X1 U36936 ( .A1(n55175), .A2(\DP/ALU0/s_A_SHIFT[7] ), .B1(
        \DP/ALU0/s_A_SHIFT[23] ), .B2(n55176), .ZN(n54423) );
  AOI22_X1 U36937 ( .A1(n54421), .A2(\DP/ALU0/s_A_SHIFT[0] ), .B1(
        \DP/ALU0/s_A_SHIFT[15] ), .B2(n55174), .ZN(n54422) );
  NAND2_X1 U36938 ( .A1(n54423), .A2(n54422), .ZN(n55144) );
  AOI22_X1 U36939 ( .A1(n55137), .A2(n54449), .B1(n53804), .B2(n54424), .ZN(
        n54426) );
  NAND2_X1 U36940 ( .A1(n53807), .A2(n54461), .ZN(n54425) );
  OAI211_X1 U36941 ( .C1(n55144), .C2(n55179), .A(n54426), .B(n54425), .ZN(
        n54446) );
  OAI22_X1 U36942 ( .A1(\intadd_0/SUM[6] ), .A2(n55303), .B1(n5463), .B2(
        n53662), .ZN(n54429) );
  NAND2_X1 U36943 ( .A1(n53809), .A2(\DP/ALU0/s_A_LOGIC[7] ), .ZN(n54427) );
  OAI22_X1 U36944 ( .A1(\DP/ALU0/S_B_LOGIC[7] ), .A2(n54427), .B1(
        \intadd_5/SUM[0] ), .B2(n55300), .ZN(n54428) );
  AOI211_X1 U36945 ( .C1(n55306), .C2(n54430), .A(n54429), .B(n54428), .ZN(
        n54433) );
  INV_X1 U36946 ( .A(\DP/ALU0/s_A_LOGIC[7] ), .ZN(n54431) );
  OAI221_X1 U36947 ( .B1(\DP/ALU0/s_A_LOGIC[7] ), .B2(n53809), .C1(n54431), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[7] ), .ZN(n54432) );
  OAI211_X1 U36948 ( .C1(n55312), .C2(n54446), .A(n54433), .B(n54432), .ZN(
        \DP/RegALU3/n92 ) );
  NAND3_X1 U36949 ( .A1(\DP/ALU0/s_A_MULT[0] ), .A2(n54437), .A3(
        \intadd_6/SUM[1] ), .ZN(\intadd_5/A[0] ) );
  AOI222_X1 U36950 ( .A1(n55175), .A2(\DP/ALU0/s_A_SHIFT[6] ), .B1(
        \DP/ALU0/s_A_SHIFT[14] ), .B2(n53808), .C1(\DP/ALU0/s_A_SHIFT[22] ), 
        .C2(n55176), .ZN(n55172) );
  INV_X1 U36951 ( .A(n54458), .ZN(n54475) );
  AOI22_X1 U36952 ( .A1(n55137), .A2(n54457), .B1(n53804), .B2(n54434), .ZN(
        n54435) );
  OAI21_X1 U36953 ( .B1(n53760), .B2(n54475), .A(n54435), .ZN(n54436) );
  AOI21_X1 U36954 ( .B1(n55139), .B2(n55172), .A(n54436), .ZN(n54452) );
  OAI22_X1 U36955 ( .A1(n49811), .A2(n5463), .B1(\intadd_0/SUM[5] ), .B2(
        n55303), .ZN(n54442) );
  NAND2_X1 U36956 ( .A1(n53809), .A2(\DP/ALU0/S_B_LOGIC[6] ), .ZN(n54440) );
  AND2_X1 U36957 ( .A1(\DP/ALU0/s_A_MULT[0] ), .A2(n54437), .ZN(n54438) );
  OAI211_X1 U36958 ( .C1(n54438), .C2(\intadd_6/SUM[1] ), .A(n55166), .B(
        \intadd_5/A[0] ), .ZN(n54439) );
  OAI21_X1 U36959 ( .B1(\DP/ALU0/s_A_LOGIC[6] ), .B2(n54440), .A(n54439), .ZN(
        n54441) );
  AOI211_X1 U36960 ( .C1(n55181), .C2(n54452), .A(n54442), .B(n54441), .ZN(
        n54445) );
  INV_X1 U36961 ( .A(\DP/ALU0/S_B_LOGIC[6] ), .ZN(n54443) );
  OAI221_X1 U36962 ( .B1(\DP/ALU0/S_B_LOGIC[6] ), .B2(n53809), .C1(n54443), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[6] ), .ZN(n54444) );
  OAI211_X1 U36963 ( .C1(n54446), .C2(n55186), .A(n54445), .B(n54444), .ZN(
        \DP/RegALU3/n93 ) );
  INV_X1 U36964 ( .A(\DP/ALU0/s_A_LOGIC[5] ), .ZN(n54453) );
  NOR3_X1 U36965 ( .A1(\DP/ALU0/S_B_LOGIC[5] ), .A2(n54453), .A3(n55187), .ZN(
        n54448) );
  OAI22_X1 U36966 ( .A1(n3249), .A2(n5463), .B1(\intadd_0/SUM[4] ), .B2(n55303), .ZN(n54447) );
  AOI211_X1 U36967 ( .C1(n55166), .C2(\intadd_6/SUM[0] ), .A(n54448), .B(
        n54447), .ZN(n54456) );
  AOI222_X1 U36968 ( .A1(n55175), .A2(\DP/ALU0/s_A_SHIFT[5] ), .B1(
        \DP/ALU0/s_A_SHIFT[13] ), .B2(n53808), .C1(\DP/ALU0/s_A_SHIFT[21] ), 
        .C2(n55176), .ZN(n55136) );
  AOI22_X1 U36969 ( .A1(n55137), .A2(n54461), .B1(n53804), .B2(n54449), .ZN(
        n54450) );
  OAI21_X1 U36970 ( .B1(n53760), .B2(n55144), .A(n54450), .ZN(n54451) );
  AOI21_X1 U36971 ( .B1(n55139), .B2(n55136), .A(n54451), .ZN(n55307) );
  AOI22_X1 U36972 ( .A1(n55181), .A2(n55307), .B1(n55306), .B2(n54452), .ZN(
        n54455) );
  OAI221_X1 U36973 ( .B1(\DP/ALU0/s_A_LOGIC[5] ), .B2(n53809), .C1(n54453), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[5] ), .ZN(n54454) );
  NAND3_X1 U36974 ( .A1(n54456), .A2(n54455), .A3(n54454), .ZN(
        \DP/RegALU3/n94 ) );
  AOI22_X1 U36975 ( .A1(n55137), .A2(n54458), .B1(n53804), .B2(n54457), .ZN(
        n54460) );
  AOI222_X1 U36976 ( .A1(\DP/ALU0/s_A_SHIFT[20] ), .A2(n55176), .B1(
        \DP/ALU0/s_A_SHIFT[12] ), .B2(n53808), .C1(n55175), .C2(
        \DP/ALU0/s_A_SHIFT[4] ), .ZN(n55178) );
  AOI22_X1 U36977 ( .A1(n53807), .A2(n55172), .B1(n55139), .B2(n55178), .ZN(
        n54459) );
  NAND2_X1 U36978 ( .A1(n54460), .A2(n54459), .ZN(n55313) );
  AOI222_X1 U36979 ( .A1(n55175), .A2(\DP/ALU0/s_A_SHIFT[3] ), .B1(
        \DP/ALU0/s_A_SHIFT[19] ), .B2(n55176), .C1(\DP/ALU0/s_A_SHIFT[11] ), 
        .C2(n53808), .ZN(n55135) );
  AOI22_X1 U36980 ( .A1(n53807), .A2(n55136), .B1(n53804), .B2(n54461), .ZN(
        n54462) );
  OAI21_X1 U36981 ( .B1(n55177), .B2(n55144), .A(n54462), .ZN(n54463) );
  AOI21_X1 U36982 ( .B1(n55139), .B2(n55135), .A(n54463), .ZN(n54477) );
  OAI22_X1 U36983 ( .A1(n3254), .A2(n5463), .B1(\intadd_7/SUM[0] ), .B2(n55300), .ZN(n54466) );
  NAND2_X1 U36984 ( .A1(n53809), .A2(\DP/ALU0/S_B_LOGIC[3] ), .ZN(n54464) );
  OAI22_X1 U36985 ( .A1(\intadd_0/SUM[2] ), .A2(n55303), .B1(
        \DP/ALU0/s_A_LOGIC[3] ), .B2(n54464), .ZN(n54465) );
  AOI211_X1 U36986 ( .C1(n55181), .C2(n54477), .A(n54466), .B(n54465), .ZN(
        n54469) );
  INV_X1 U36987 ( .A(\DP/ALU0/S_B_LOGIC[3] ), .ZN(n54467) );
  OAI221_X1 U36988 ( .B1(\DP/ALU0/S_B_LOGIC[3] ), .B2(n53809), .C1(n54467), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[3] ), .ZN(n54468) );
  OAI211_X1 U36989 ( .C1(n55313), .C2(n55186), .A(n54469), .B(n54468), .ZN(
        \DP/RegALU3/n96 ) );
  INV_X1 U36990 ( .A(\DP/ALU0/s_A_MULT[1] ), .ZN(n54918) );
  AOI22_X1 U36991 ( .A1(\DP/ALU0/s_A_MULT[0] ), .A2(n54918), .B1(
        \DP/ALU0/s_A_MULT[1] ), .B2(n55299), .ZN(n54915) );
  INV_X1 U36992 ( .A(n54915), .ZN(n54881) );
  NAND2_X1 U36993 ( .A1(n55299), .A2(n54918), .ZN(n54470) );
  NAND2_X1 U36994 ( .A1(\DP/ALU0/S_B_MULT[1] ), .A2(\DP/ALU0/S_B_MULT[0] ), 
        .ZN(n54859) );
  AOI222_X1 U36995 ( .A1(n54881), .A2(n54864), .B1(n54865), .B2(
        \DP/ALU0/s_A_MULT[2] ), .C1(n54885), .C2(n54863), .ZN(n54471) );
  INV_X1 U36996 ( .A(n54471), .ZN(n54479) );
  NAND3_X1 U36997 ( .A1(n54478), .A2(\DP/ALU0/s_A_MULT[0] ), .A3(n54479), .ZN(
        \intadd_7/A[0] ) );
  NOR2_X1 U36998 ( .A1(\DP/ALU0/s_A_LOGIC[2] ), .A2(n55187), .ZN(n54473) );
  OAI22_X1 U36999 ( .A1(n3247), .A2(n5463), .B1(\intadd_0/SUM[1] ), .B2(n55303), .ZN(n54472) );
  AOI21_X1 U37000 ( .B1(n54473), .B2(\DP/ALU0/S_B_LOGIC[2] ), .A(n54472), .ZN(
        n54485) );
  AOI222_X1 U37001 ( .A1(\DP/ALU0/s_A_SHIFT[18] ), .A2(n55176), .B1(
        \DP/ALU0/s_A_SHIFT[10] ), .B2(n53808), .C1(n55175), .C2(
        \DP/ALU0/s_A_SHIFT[2] ), .ZN(n55173) );
  AOI22_X1 U37002 ( .A1(n53807), .A2(n55178), .B1(n55139), .B2(n55173), .ZN(
        n54474) );
  OAI21_X1 U37003 ( .B1(n53761), .B2(n54475), .A(n54474), .ZN(n54476) );
  AOI21_X1 U37004 ( .B1(n55137), .B2(n55172), .A(n54476), .ZN(n55193) );
  AOI22_X1 U37005 ( .A1(n55181), .A2(n55193), .B1(n55306), .B2(n54477), .ZN(
        n54484) );
  AND2_X1 U37006 ( .A1(\DP/ALU0/s_A_MULT[0] ), .A2(n54478), .ZN(n54480) );
  OAI211_X1 U37007 ( .C1(n54480), .C2(n54479), .A(n55166), .B(\intadd_7/A[0] ), 
        .ZN(n54483) );
  INV_X1 U37008 ( .A(\DP/ALU0/S_B_LOGIC[2] ), .ZN(n54481) );
  OAI221_X1 U37009 ( .B1(\DP/ALU0/S_B_LOGIC[2] ), .B2(n53809), .C1(n54481), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[2] ), .ZN(n54482) );
  NAND4_X1 U37010 ( .A1(n54485), .A2(n54484), .A3(n54483), .A4(n54482), .ZN(
        \DP/RegALU3/n97 ) );
  INV_X1 U37011 ( .A(n55330), .ZN(n54490) );
  AOI221_X1 U37012 ( .B1(n53561), .B2(n55330), .C1(n53704), .C2(n54490), .A(
        n45959), .ZN(n54486) );
  NOR2_X1 U37013 ( .A1(n54486), .A2(n53820), .ZN(\DP/RegRD2/n10 ) );
  AOI221_X1 U37014 ( .B1(n53556), .B2(n54490), .C1(n53560), .C2(n55330), .A(
        n45959), .ZN(n54487) );
  NOR2_X1 U37015 ( .A1(n54487), .A2(n53822), .ZN(\DP/RegRD2/n11 ) );
  AOI221_X1 U37016 ( .B1(n53555), .B2(n54490), .C1(n53559), .C2(n55330), .A(
        n45959), .ZN(n54488) );
  NOR2_X1 U37017 ( .A1(n54488), .A2(n53819), .ZN(\DP/RegRD2/n12 ) );
  AOI221_X1 U37018 ( .B1(n53554), .B2(n54490), .C1(n53558), .C2(n55330), .A(
        n45959), .ZN(n54489) );
  NOR2_X1 U37019 ( .A1(n54489), .A2(n53819), .ZN(\DP/RegRD2/n13 ) );
  AOI221_X1 U37020 ( .B1(n53553), .B2(n54490), .C1(n53557), .C2(n55330), .A(
        n45959), .ZN(n54491) );
  NOR2_X1 U37021 ( .A1(n54491), .A2(n53822), .ZN(\DP/RegRD2/n14 ) );
  NAND2_X1 U37022 ( .A1(RST), .A2(n3019), .ZN(\DP/RegRD2/n7 ) );
  AND2_X1 U37023 ( .A1(RST), .A2(n53266), .ZN(\DP/RegRD3/n10 ) );
  AND2_X1 U37024 ( .A1(RST), .A2(n53267), .ZN(\DP/RegRD3/n11 ) );
  AND2_X1 U37025 ( .A1(RST), .A2(n53268), .ZN(\DP/RegRD3/n12 ) );
  AND2_X1 U37026 ( .A1(RST), .A2(n53269), .ZN(\DP/RegRD3/n13 ) );
  AND2_X1 U37027 ( .A1(RST), .A2(n53270), .ZN(\DP/RegRD3/n14 ) );
  AND2_X1 U37028 ( .A1(RST), .A2(n49866), .ZN(\DP/RegRD4/n10 ) );
  AND2_X1 U37029 ( .A1(RST), .A2(n49819), .ZN(\DP/RegRD4/n11 ) );
  NOR2_X1 U37030 ( .A1(n53820), .A2(n53673), .ZN(\DP/RegRD4/n12 ) );
  NOR2_X1 U37031 ( .A1(n7617), .A2(n53821), .ZN(\DP/RegRD4/n13 ) );
  NOR2_X1 U37032 ( .A1(n53819), .A2(n53693), .ZN(\DP/RegRD4/n14 ) );
  NAND2_X1 U37033 ( .A1(RST), .A2(n3021), .ZN(\DP/RegRD4/n7 ) );
  NOR2_X1 U37034 ( .A1(n53647), .A2(n53281), .ZN(n54492) );
  AOI221_X1 U37035 ( .B1(n53280), .B2(n54548), .C1(n54530), .C2(n54548), .A(
        n54492), .ZN(n55249) );
  NOR4_X1 U37036 ( .A1(\DP/RD4[2] ), .A2(\DP/RD4[3] ), .A3(\DP/RD4[4] ), .A4(
        \DP/RD4[1] ), .ZN(n54499) );
  AOI22_X1 U37037 ( .A1(\DP/RD4[4] ), .A2(n53274), .B1(\DP/RD4[0] ), .B2(
        n53273), .ZN(n54493) );
  OAI221_X1 U37038 ( .B1(\DP/RD4[4] ), .B2(n53274), .C1(\DP/RD4[0] ), .C2(
        n53273), .A(n54493), .ZN(n54498) );
  AOI22_X1 U37039 ( .A1(\DP/RD4[3] ), .A2(n53271), .B1(n53272), .B2(
        \DP/RD4[1] ), .ZN(n54494) );
  OAI221_X1 U37040 ( .B1(\DP/RD4[3] ), .B2(n53271), .C1(\DP/RD4[1] ), .C2(
        n53272), .A(n54494), .ZN(n54495) );
  AOI211_X1 U37041 ( .C1(n3015), .C2(n53275), .A(n53654), .B(n54495), .ZN(
        n54496) );
  OAI21_X1 U37042 ( .B1(n3015), .B2(n53275), .A(n54496), .ZN(n54497) );
  AOI21_X1 U37043 ( .B1(n53277), .B2(n54548), .A(n54547), .ZN(n54500) );
  OAI21_X1 U37044 ( .B1(n53647), .B2(n53276), .A(n54500), .ZN(n55214) );
  AOI22_X1 U37045 ( .A1(n54537), .A2(n53278), .B1(n55214), .B2(n54536), .ZN(
        n54596) );
  AOI22_X1 U37046 ( .A1(n55249), .A2(n54593), .B1(n54582), .B2(n54596), .ZN(
        n54505) );
  INV_X1 U37047 ( .A(n54530), .ZN(n54507) );
  OR2_X1 U37048 ( .A1(n54507), .A2(n54506), .ZN(n54502) );
  OAI21_X1 U37049 ( .B1(n54502), .B2(n54501), .A(n53647), .ZN(n54588) );
  OAI22_X1 U37050 ( .A1(n53647), .A2(n53283), .B1(n53282), .B2(n54588), .ZN(
        n55205) );
  NAND2_X1 U37051 ( .A1(n54537), .A2(n54602), .ZN(n54591) );
  OAI22_X1 U37052 ( .A1(n53279), .A2(n54606), .B1(n53318), .B2(n54591), .ZN(
        n54503) );
  AOI21_X1 U37053 ( .B1(n55205), .B2(n53805), .A(n54503), .ZN(n54504) );
  NAND2_X1 U37054 ( .A1(n54505), .A2(n54504), .ZN(DRAM_DATA_OUT[0]) );
  NOR2_X1 U37055 ( .A1(n53284), .A2(n54598), .ZN(n54508) );
  AOI211_X1 U37056 ( .C1(n53285), .C2(n53684), .A(n54508), .B(n54599), .ZN(
        n55238) );
  AOI21_X1 U37057 ( .B1(n53287), .B2(n54548), .A(n54547), .ZN(n54509) );
  OAI21_X1 U37058 ( .B1(n53647), .B2(n53286), .A(n54509), .ZN(n55209) );
  AOI22_X1 U37059 ( .A1(n54537), .A2(n53288), .B1(n55209), .B2(n54536), .ZN(
        n54557) );
  AOI22_X1 U37060 ( .A1(n55238), .A2(n54603), .B1(n54602), .B2(n54557), .ZN(
        n54512) );
  NAND2_X1 U37061 ( .A1(n54536), .A2(n54510), .ZN(n54511) );
  OAI21_X1 U37062 ( .B1(n54536), .B2(n53290), .A(n54511), .ZN(n54563) );
  NAND2_X1 U37063 ( .A1(n54563), .A2(n54582), .ZN(n54604) );
  OAI211_X1 U37064 ( .C1(n53289), .C2(n54606), .A(n54512), .B(n54604), .ZN(
        DRAM_DATA_OUT[10]) );
  NOR2_X1 U37065 ( .A1(n53295), .A2(n54598), .ZN(n54513) );
  AOI211_X1 U37066 ( .C1(n53294), .C2(n53684), .A(n54513), .B(n54599), .ZN(
        n55241) );
  AOI21_X1 U37067 ( .B1(n53292), .B2(n54548), .A(n54547), .ZN(n54514) );
  OAI21_X1 U37068 ( .B1(n53647), .B2(n53291), .A(n54514), .ZN(n55210) );
  AOI22_X1 U37069 ( .A1(n54537), .A2(n53293), .B1(n55210), .B2(n54536), .ZN(
        n54567) );
  AOI22_X1 U37070 ( .A1(n55241), .A2(n53805), .B1(n54602), .B2(n54567), .ZN(
        n54515) );
  OAI211_X1 U37071 ( .C1(n53296), .C2(n54606), .A(n54515), .B(n54604), .ZN(
        DRAM_DATA_OUT[11]) );
  NOR2_X1 U37072 ( .A1(n53301), .A2(n54598), .ZN(n54516) );
  AOI211_X1 U37073 ( .C1(n53300), .C2(n53684), .A(n54516), .B(n54599), .ZN(
        n55240) );
  AOI21_X1 U37074 ( .B1(n53298), .B2(n54548), .A(n54547), .ZN(n54517) );
  OAI21_X1 U37075 ( .B1(n53647), .B2(n53297), .A(n54517), .ZN(n55221) );
  AOI22_X1 U37076 ( .A1(n54537), .A2(n53299), .B1(n55221), .B2(n54536), .ZN(
        n54572) );
  AOI22_X1 U37077 ( .A1(n55240), .A2(n54603), .B1(n54602), .B2(n54572), .ZN(
        n54518) );
  OAI211_X1 U37078 ( .C1(n53302), .C2(n54606), .A(n54518), .B(n54604), .ZN(
        DRAM_DATA_OUT[12]) );
  AOI21_X1 U37079 ( .B1(n53307), .B2(n53684), .A(n54599), .ZN(n54519) );
  OAI21_X1 U37080 ( .B1(n53306), .B2(n54598), .A(n54519), .ZN(n55243) );
  INV_X1 U37081 ( .A(n55243), .ZN(n55097) );
  AOI21_X1 U37082 ( .B1(n53304), .B2(n54548), .A(n54547), .ZN(n54520) );
  OAI21_X1 U37083 ( .B1(n53647), .B2(n53303), .A(n54520), .ZN(n55222) );
  AOI22_X1 U37084 ( .A1(n54537), .A2(n53305), .B1(n55222), .B2(n54536), .ZN(
        n54577) );
  AOI22_X1 U37085 ( .A1(n55097), .A2(n53805), .B1(n54602), .B2(n54577), .ZN(
        n54521) );
  OAI211_X1 U37086 ( .C1(n53308), .C2(n54606), .A(n54521), .B(n54604), .ZN(
        DRAM_DATA_OUT[13]) );
  NOR2_X1 U37087 ( .A1(n53312), .A2(n54598), .ZN(n54522) );
  AOI211_X1 U37088 ( .C1(n53313), .C2(n53684), .A(n54522), .B(n54599), .ZN(
        n55237) );
  AOI21_X1 U37089 ( .B1(n53310), .B2(n54548), .A(n54547), .ZN(n54523) );
  OAI21_X1 U37090 ( .B1(n53647), .B2(n53309), .A(n54523), .ZN(n55223) );
  AOI22_X1 U37091 ( .A1(n54537), .A2(n53311), .B1(n55223), .B2(n54536), .ZN(
        n54583) );
  AOI22_X1 U37092 ( .A1(n55237), .A2(n54603), .B1(n54602), .B2(n54583), .ZN(
        n54524) );
  OAI211_X1 U37093 ( .C1(n53314), .C2(n54606), .A(n54524), .B(n54604), .ZN(
        DRAM_DATA_OUT[14]) );
  NOR2_X1 U37094 ( .A1(n53315), .A2(n54598), .ZN(n54525) );
  AOI211_X1 U37095 ( .C1(n53316), .C2(n53684), .A(n54599), .B(n54525), .ZN(
        n55236) );
  NAND2_X1 U37096 ( .A1(n55236), .A2(n53805), .ZN(n54526) );
  OAI211_X1 U37097 ( .C1(n53317), .C2(n54606), .A(n54564), .B(n54526), .ZN(
        DRAM_DATA_OUT[15]) );
  NAND2_X1 U37098 ( .A1(n55249), .A2(n54603), .ZN(n54527) );
  OAI211_X1 U37099 ( .C1(n53318), .C2(n54606), .A(n54564), .B(n54527), .ZN(
        DRAM_DATA_OUT[16]) );
  NOR2_X1 U37100 ( .A1(n53647), .A2(n53320), .ZN(n54528) );
  AOI221_X1 U37101 ( .B1(n53319), .B2(n54548), .C1(n54530), .C2(n54548), .A(
        n54528), .ZN(n55250) );
  NAND2_X1 U37102 ( .A1(n55250), .A2(n53805), .ZN(n54529) );
  OAI211_X1 U37103 ( .C1(n53328), .C2(n54606), .A(n54564), .B(n54529), .ZN(
        DRAM_DATA_OUT[17]) );
  OAI21_X1 U37104 ( .B1(n53321), .B2(n54530), .A(n54548), .ZN(n54531) );
  OAI21_X1 U37105 ( .B1(n53647), .B2(n53322), .A(n54531), .ZN(n55201) );
  INV_X1 U37106 ( .A(n55201), .ZN(n54559) );
  NAND2_X1 U37107 ( .A1(n54559), .A2(n53805), .ZN(n54532) );
  OAI211_X1 U37108 ( .C1(n53342), .C2(n54606), .A(n54564), .B(n54532), .ZN(
        DRAM_DATA_OUT[18]) );
  AOI21_X1 U37109 ( .B1(n53324), .B2(n54548), .A(n54547), .ZN(n54533) );
  OAI21_X1 U37110 ( .B1(n53647), .B2(n53323), .A(n54533), .ZN(n55220) );
  INV_X1 U37111 ( .A(n55220), .ZN(n54569) );
  NAND2_X1 U37112 ( .A1(n54569), .A2(n54603), .ZN(n54534) );
  OAI211_X1 U37113 ( .C1(n53344), .C2(n54606), .A(n54564), .B(n54534), .ZN(
        DRAM_DATA_OUT[19]) );
  AOI21_X1 U37114 ( .B1(n53326), .B2(n54548), .A(n54547), .ZN(n54535) );
  OAI21_X1 U37115 ( .B1(n53647), .B2(n53325), .A(n54535), .ZN(n55203) );
  AOI22_X1 U37116 ( .A1(n54537), .A2(n53327), .B1(n55203), .B2(n54536), .ZN(
        n54601) );
  OAI22_X1 U37117 ( .A1(n53647), .A2(n53331), .B1(n53330), .B2(n54588), .ZN(
        n55208) );
  AOI22_X1 U37118 ( .A1(n54601), .A2(n54582), .B1(n53805), .B2(n55208), .ZN(
        n54540) );
  OAI22_X1 U37119 ( .A1(n53328), .A2(n54591), .B1(n53329), .B2(n54606), .ZN(
        n54538) );
  AOI21_X1 U37120 ( .B1(n55250), .B2(n54593), .A(n54538), .ZN(n54539) );
  NAND2_X1 U37121 ( .A1(n54540), .A2(n54539), .ZN(DRAM_DATA_OUT[1]) );
  AOI21_X1 U37122 ( .B1(n53333), .B2(n54548), .A(n54547), .ZN(n54541) );
  OAI21_X1 U37123 ( .B1(n53647), .B2(n53332), .A(n54541), .ZN(n55202) );
  INV_X1 U37124 ( .A(n55202), .ZN(n54574) );
  NAND2_X1 U37125 ( .A1(n54574), .A2(n54603), .ZN(n54542) );
  OAI211_X1 U37126 ( .C1(n53348), .C2(n54606), .A(n54564), .B(n54542), .ZN(
        DRAM_DATA_OUT[20]) );
  AOI21_X1 U37127 ( .B1(n53335), .B2(n54548), .A(n54547), .ZN(n54543) );
  OAI21_X1 U37128 ( .B1(n53647), .B2(n53334), .A(n54543), .ZN(n55212) );
  INV_X1 U37129 ( .A(n55212), .ZN(n54579) );
  NAND2_X1 U37130 ( .A1(n54579), .A2(n53805), .ZN(n54544) );
  OAI211_X1 U37131 ( .C1(n53352), .C2(n54606), .A(n54564), .B(n54544), .ZN(
        DRAM_DATA_OUT[21]) );
  AOI21_X1 U37132 ( .B1(n53337), .B2(n54548), .A(n54547), .ZN(n54545) );
  OAI21_X1 U37133 ( .B1(n53647), .B2(n53336), .A(n54545), .ZN(n55213) );
  INV_X1 U37134 ( .A(n55213), .ZN(n54585) );
  NAND2_X1 U37135 ( .A1(n54585), .A2(n54603), .ZN(n54546) );
  OAI211_X1 U37136 ( .C1(n53356), .C2(n54606), .A(n54564), .B(n54546), .ZN(
        DRAM_DATA_OUT[22]) );
  AOI21_X1 U37137 ( .B1(n53339), .B2(n54548), .A(n54547), .ZN(n54549) );
  OAI21_X1 U37138 ( .B1(n53647), .B2(n53338), .A(n54549), .ZN(n55052) );
  INV_X1 U37139 ( .A(n55052), .ZN(n55219) );
  NAND2_X1 U37140 ( .A1(n55219), .A2(n53805), .ZN(n54550) );
  OAI211_X1 U37141 ( .C1(n53595), .C2(n54606), .A(n54564), .B(n54550), .ZN(
        DRAM_DATA_OUT[23]) );
  INV_X1 U37142 ( .A(n54596), .ZN(n54551) );
  OAI21_X1 U37143 ( .B1(n54551), .B2(n54566), .A(n54564), .ZN(
        DRAM_DATA_OUT[24]) );
  INV_X1 U37144 ( .A(n54601), .ZN(n54552) );
  OAI21_X1 U37145 ( .B1(n54552), .B2(n54566), .A(n54564), .ZN(
        DRAM_DATA_OUT[25]) );
  INV_X1 U37146 ( .A(n54557), .ZN(n54553) );
  OAI21_X1 U37147 ( .B1(n54553), .B2(n54566), .A(n54564), .ZN(
        DRAM_DATA_OUT[26]) );
  INV_X1 U37148 ( .A(n54567), .ZN(n54554) );
  OAI21_X1 U37149 ( .B1(n54554), .B2(n54566), .A(n54564), .ZN(
        DRAM_DATA_OUT[27]) );
  INV_X1 U37150 ( .A(n54572), .ZN(n54555) );
  OAI21_X1 U37151 ( .B1(n54555), .B2(n54566), .A(n54564), .ZN(
        DRAM_DATA_OUT[28]) );
  INV_X1 U37152 ( .A(n54577), .ZN(n54556) );
  OAI21_X1 U37153 ( .B1(n54556), .B2(n54566), .A(n54564), .ZN(
        DRAM_DATA_OUT[29]) );
  OAI22_X1 U37154 ( .A1(n53647), .A2(n53341), .B1(n53340), .B2(n54588), .ZN(
        n55336) );
  AOI22_X1 U37155 ( .A1(n54557), .A2(n54582), .B1(n54603), .B2(n55336), .ZN(
        n54561) );
  OAI22_X1 U37156 ( .A1(n53342), .A2(n54591), .B1(n53343), .B2(n54606), .ZN(
        n54558) );
  AOI21_X1 U37157 ( .B1(n54559), .B2(n54593), .A(n54558), .ZN(n54560) );
  NAND2_X1 U37158 ( .A1(n54561), .A2(n54560), .ZN(DRAM_DATA_OUT[2]) );
  INV_X1 U37159 ( .A(n54583), .ZN(n54562) );
  OAI21_X1 U37160 ( .B1(n54562), .B2(n54566), .A(n54564), .ZN(
        DRAM_DATA_OUT[30]) );
  INV_X1 U37161 ( .A(n54563), .ZN(n54565) );
  OAI21_X1 U37162 ( .B1(n54566), .B2(n54565), .A(n54564), .ZN(
        DRAM_DATA_OUT[31]) );
  OAI22_X1 U37163 ( .A1(n53647), .A2(n53347), .B1(n53346), .B2(n54588), .ZN(
        n55239) );
  AOI22_X1 U37164 ( .A1(n54567), .A2(n54582), .B1(n53805), .B2(n55239), .ZN(
        n54571) );
  OAI22_X1 U37165 ( .A1(n53344), .A2(n54591), .B1(n53345), .B2(n54606), .ZN(
        n54568) );
  AOI21_X1 U37166 ( .B1(n54569), .B2(n54593), .A(n54568), .ZN(n54570) );
  NAND2_X1 U37167 ( .A1(n54571), .A2(n54570), .ZN(DRAM_DATA_OUT[3]) );
  OAI22_X1 U37168 ( .A1(n53647), .A2(n53351), .B1(n53350), .B2(n54588), .ZN(
        n55206) );
  AOI22_X1 U37169 ( .A1(n54572), .A2(n54582), .B1(n53805), .B2(n55206), .ZN(
        n54576) );
  OAI22_X1 U37170 ( .A1(n53348), .A2(n54591), .B1(n53349), .B2(n54606), .ZN(
        n54573) );
  AOI21_X1 U37171 ( .B1(n54574), .B2(n54593), .A(n54573), .ZN(n54575) );
  NAND2_X1 U37172 ( .A1(n54576), .A2(n54575), .ZN(DRAM_DATA_OUT[4]) );
  OAI22_X1 U37173 ( .A1(n53647), .A2(n53355), .B1(n53354), .B2(n54588), .ZN(
        n55207) );
  AOI22_X1 U37174 ( .A1(n54577), .A2(n54582), .B1(n54603), .B2(n55207), .ZN(
        n54581) );
  OAI22_X1 U37175 ( .A1(n53352), .A2(n54591), .B1(n53353), .B2(n54606), .ZN(
        n54578) );
  AOI21_X1 U37176 ( .B1(n54579), .B2(n54593), .A(n54578), .ZN(n54580) );
  NAND2_X1 U37177 ( .A1(n54581), .A2(n54580), .ZN(DRAM_DATA_OUT[5]) );
  OAI22_X1 U37178 ( .A1(n53647), .A2(n53359), .B1(n53358), .B2(n54588), .ZN(
        n55334) );
  AOI22_X1 U37179 ( .A1(n54583), .A2(n54582), .B1(n53805), .B2(n55334), .ZN(
        n54587) );
  OAI22_X1 U37180 ( .A1(n53356), .A2(n54591), .B1(n53357), .B2(n54606), .ZN(
        n54584) );
  AOI21_X1 U37181 ( .B1(n54585), .B2(n54593), .A(n54584), .ZN(n54586) );
  NAND2_X1 U37182 ( .A1(n54587), .A2(n54586), .ZN(DRAM_DATA_OUT[6]) );
  INV_X1 U37183 ( .A(n54588), .ZN(n54590) );
  NOR2_X1 U37184 ( .A1(n53647), .A2(n53371), .ZN(n54589) );
  AOI21_X1 U37185 ( .B1(n49869), .B2(n54590), .A(n54589), .ZN(n55204) );
  OAI22_X1 U37186 ( .A1(n53595), .A2(n54591), .B1(n53596), .B2(n54606), .ZN(
        n54592) );
  AOI21_X1 U37187 ( .B1(n55219), .B2(n54593), .A(n54592), .ZN(n54594) );
  OAI211_X1 U37188 ( .C1(n55204), .C2(n53806), .A(n54594), .B(n54604), .ZN(
        DRAM_DATA_OUT[7]) );
  NOR2_X1 U37189 ( .A1(n53360), .A2(n54598), .ZN(n54595) );
  AOI211_X1 U37190 ( .C1(n53361), .C2(n53684), .A(n54595), .B(n54599), .ZN(
        n55242) );
  AOI22_X1 U37191 ( .A1(n55242), .A2(n53805), .B1(n54602), .B2(n54596), .ZN(
        n54597) );
  OAI211_X1 U37192 ( .C1(n53362), .C2(n54606), .A(n54597), .B(n54604), .ZN(
        DRAM_DATA_OUT[8]) );
  NOR2_X1 U37193 ( .A1(n53363), .A2(n54598), .ZN(n54600) );
  AOI211_X1 U37194 ( .C1(n53364), .C2(n53684), .A(n54600), .B(n54599), .ZN(
        n55235) );
  AOI22_X1 U37195 ( .A1(n55235), .A2(n54603), .B1(n54602), .B2(n54601), .ZN(
        n54605) );
  OAI211_X1 U37196 ( .C1(n53365), .C2(n54606), .A(n54605), .B(n54604), .ZN(
        DRAM_DATA_OUT[9]) );
  XNOR2_X1 U37197 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[1] ), .ZN(
        \intadd_0/B[0] ) );
  XNOR2_X1 U37198 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[11] ), .ZN(
        \intadd_0/B[10] ) );
  XNOR2_X1 U37199 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[12] ), .ZN(
        \intadd_0/B[11] ) );
  XNOR2_X1 U37200 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[13] ), .ZN(
        \intadd_0/B[12] ) );
  XNOR2_X1 U37201 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[14] ), .ZN(
        \intadd_0/B[13] ) );
  XNOR2_X1 U37202 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[15] ), .ZN(
        \intadd_0/B[14] ) );
  XNOR2_X1 U37203 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[16] ), .ZN(
        \intadd_0/B[15] ) );
  XNOR2_X1 U37204 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[17] ), .ZN(
        \intadd_0/B[16] ) );
  XNOR2_X1 U37205 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[18] ), .ZN(
        \intadd_0/B[17] ) );
  XNOR2_X1 U37206 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[19] ), .ZN(
        \intadd_0/B[18] ) );
  XNOR2_X1 U37207 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[20] ), .ZN(
        \intadd_0/B[19] ) );
  XNOR2_X1 U37208 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[2] ), .ZN(
        \intadd_0/B[1] ) );
  XNOR2_X1 U37209 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[21] ), .ZN(
        \intadd_0/B[20] ) );
  XNOR2_X1 U37210 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[22] ), .ZN(
        \intadd_0/B[21] ) );
  XNOR2_X1 U37211 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[23] ), .ZN(
        \intadd_0/B[22] ) );
  XNOR2_X1 U37212 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[24] ), .ZN(
        \intadd_0/B[23] ) );
  XNOR2_X1 U37213 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[25] ), .ZN(
        \intadd_0/B[24] ) );
  XNOR2_X1 U37214 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[26] ), .ZN(
        \intadd_0/B[25] ) );
  XNOR2_X1 U37215 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[27] ), .ZN(
        \intadd_0/B[26] ) );
  XNOR2_X1 U37216 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[3] ), .ZN(
        \intadd_0/B[2] ) );
  XNOR2_X1 U37217 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[4] ), .ZN(
        \intadd_0/B[3] ) );
  XNOR2_X1 U37218 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[5] ), .ZN(
        \intadd_0/B[4] ) );
  XNOR2_X1 U37219 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[6] ), .ZN(
        \intadd_0/B[5] ) );
  XNOR2_X1 U37220 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[7] ), .ZN(
        \intadd_0/B[6] ) );
  XNOR2_X1 U37221 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[8] ), .ZN(
        \intadd_0/B[7] ) );
  XNOR2_X1 U37222 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[9] ), .ZN(
        \intadd_0/B[8] ) );
  XNOR2_X1 U37223 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[10] ), .ZN(
        \intadd_0/B[9] ) );
  INV_X1 U37224 ( .A(\DP/ALU0/S_B_ADDER[0] ), .ZN(n54607) );
  AOI22_X1 U37225 ( .A1(\DP/ALU0/S_B_ADDER[0] ), .A2(\DP/ALU0/s_A_ADDER[0] ), 
        .B1(n53817), .B2(n54607), .ZN(\intadd_0/CI ) );
  NAND2_X1 U37226 ( .A1(\intadd_2/n1 ), .A2(n54608), .ZN(n54612) );
  OAI21_X1 U37227 ( .B1(\intadd_2/n1 ), .B2(n54608), .A(n54612), .ZN(n54609)
         );
  XOR2_X1 U37228 ( .A(n54610), .B(n54609), .Z(\intadd_1/A[11] ) );
  NAND2_X1 U37229 ( .A1(n54612), .A2(n54611), .ZN(n54614) );
  XNOR2_X1 U37230 ( .A(n54614), .B(n54613), .ZN(\intadd_1/A[12] ) );
  INV_X1 U37231 ( .A(n54870), .ZN(n54867) );
  AOI22_X1 U37232 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n54661), .B1(
        \DP/ALU0/s_A_MULT[10] ), .B2(n54659), .ZN(n54619) );
  NAND2_X1 U37233 ( .A1(n53642), .A2(n54869), .ZN(n54618) );
  OAI211_X1 U37234 ( .C1(n54867), .C2(n54664), .A(n54619), .B(n54618), .ZN(
        \intadd_1/B[10] ) );
  OAI21_X1 U37235 ( .B1(n54622), .B2(n54621), .A(n54620), .ZN(n54872) );
  AOI22_X1 U37236 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n54661), .B1(n53642), 
        .B2(n54870), .ZN(n54624) );
  NAND2_X1 U37237 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n54659), .ZN(n54623) );
  OAI211_X1 U37238 ( .C1(n54872), .C2(n54664), .A(n54624), .B(n54623), .ZN(
        \intadd_1/B[11] ) );
  INV_X1 U37239 ( .A(n54856), .ZN(n54876) );
  AOI22_X1 U37240 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54661), .B1(
        \DP/ALU0/s_A_MULT[12] ), .B2(n54659), .ZN(n54626) );
  INV_X1 U37241 ( .A(n54872), .ZN(n54874) );
  NAND2_X1 U37242 ( .A1(n53642), .A2(n54874), .ZN(n54625) );
  OAI211_X1 U37243 ( .C1(n54876), .C2(n54664), .A(n54626), .B(n54625), .ZN(
        \intadd_1/B[12] ) );
  INV_X1 U37244 ( .A(n54885), .ZN(n54879) );
  AOI22_X1 U37245 ( .A1(\DP/ALU0/s_A_MULT[2] ), .A2(n54661), .B1(
        \DP/ALU0/s_A_MULT[1] ), .B2(n54659), .ZN(n54628) );
  NAND2_X1 U37246 ( .A1(n53642), .A2(n54881), .ZN(n54627) );
  OAI211_X1 U37247 ( .C1(n54879), .C2(n54664), .A(n54628), .B(n54627), .ZN(
        \intadd_1/B[1] ) );
  OAI21_X1 U37248 ( .B1(n54630), .B2(n54629), .A(n54634), .ZN(n54883) );
  AOI22_X1 U37249 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n54661), .B1(
        \DP/ALU0/s_A_MULT[2] ), .B2(n54659), .ZN(n54632) );
  NAND2_X1 U37250 ( .A1(n53642), .A2(n54885), .ZN(n54631) );
  OAI211_X1 U37251 ( .C1(n54883), .C2(n54664), .A(n54632), .B(n54631), .ZN(
        \intadd_1/B[2] ) );
  INV_X1 U37252 ( .A(n54890), .ZN(n54888) );
  INV_X1 U37253 ( .A(n54883), .ZN(n54886) );
  AOI22_X1 U37254 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54661), .B1(n53642), .B2(
        n54886), .ZN(n54636) );
  NAND2_X1 U37255 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n54659), .ZN(n54635) );
  OAI211_X1 U37256 ( .C1(n54888), .C2(n54664), .A(n54636), .B(n54635), .ZN(
        \intadd_1/B[3] ) );
  INV_X1 U37257 ( .A(n54894), .ZN(n54892) );
  AOI22_X1 U37258 ( .A1(\DP/ALU0/s_A_MULT[5] ), .A2(n54661), .B1(n53642), .B2(
        n54890), .ZN(n54640) );
  NAND2_X1 U37259 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54659), .ZN(n54639) );
  OAI211_X1 U37260 ( .C1(n54892), .C2(n54664), .A(n54640), .B(n54639), .ZN(
        \intadd_1/B[4] ) );
  INV_X1 U37261 ( .A(n54898), .ZN(n54896) );
  AOI22_X1 U37262 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54661), .B1(n53642), .B2(
        n54894), .ZN(n54644) );
  NAND2_X1 U37263 ( .A1(\DP/ALU0/s_A_MULT[5] ), .A2(n54659), .ZN(n54643) );
  OAI211_X1 U37264 ( .C1(n54896), .C2(n54664), .A(n54644), .B(n54643), .ZN(
        \intadd_1/B[5] ) );
  INV_X1 U37265 ( .A(n54902), .ZN(n54900) );
  AOI22_X1 U37266 ( .A1(\DP/ALU0/s_A_MULT[7] ), .A2(n54661), .B1(n53642), .B2(
        n54898), .ZN(n54648) );
  NAND2_X1 U37267 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54659), .ZN(n54647) );
  OAI211_X1 U37268 ( .C1(n54900), .C2(n54664), .A(n54648), .B(n54647), .ZN(
        \intadd_1/B[6] ) );
  INV_X1 U37269 ( .A(n54906), .ZN(n54904) );
  AOI22_X1 U37270 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54661), .B1(n53642), .B2(
        n54902), .ZN(n54652) );
  NAND2_X1 U37271 ( .A1(\DP/ALU0/s_A_MULT[7] ), .A2(n54659), .ZN(n54651) );
  OAI211_X1 U37272 ( .C1(n54904), .C2(n54664), .A(n54652), .B(n54651), .ZN(
        \intadd_1/B[7] ) );
  INV_X1 U37273 ( .A(n54914), .ZN(n54908) );
  AOI22_X1 U37274 ( .A1(\DP/ALU0/s_A_MULT[9] ), .A2(n54661), .B1(n53642), .B2(
        n54906), .ZN(n54656) );
  NAND2_X1 U37275 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54659), .ZN(n54655) );
  OAI211_X1 U37276 ( .C1(n54908), .C2(n54664), .A(n54656), .B(n54655), .ZN(
        \intadd_1/B[8] ) );
  INV_X1 U37277 ( .A(n54869), .ZN(n54912) );
  AOI22_X1 U37278 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n54661), .B1(
        \DP/ALU0/s_A_MULT[9] ), .B2(n54659), .ZN(n54658) );
  NAND2_X1 U37279 ( .A1(n53642), .A2(n54914), .ZN(n54657) );
  OAI211_X1 U37280 ( .C1(n54912), .C2(n54664), .A(n54658), .B(n54657), .ZN(
        \intadd_1/B[9] ) );
  NOR2_X1 U37281 ( .A1(n53642), .A2(n54659), .ZN(n54663) );
  INV_X1 U37282 ( .A(n54661), .ZN(n54662) );
  OAI222_X1 U37283 ( .A1(n54915), .A2(n54664), .B1(n55299), .B2(n54663), .C1(
        n54918), .C2(n54662), .ZN(\intadd_1/CI ) );
  AOI22_X1 U37284 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n54687), .B1(
        \DP/ALU0/s_A_MULT[10] ), .B2(n54693), .ZN(n54665) );
  OAI21_X1 U37285 ( .B1(n54690), .B2(n54867), .A(n54665), .ZN(n54666) );
  AOI21_X1 U37286 ( .B1(n53644), .B2(n54869), .A(n54666), .ZN(\intadd_2/A[10] ) );
  AOI22_X1 U37287 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n54687), .B1(n53644), 
        .B2(n54870), .ZN(n54667) );
  OAI21_X1 U37288 ( .B1(n54690), .B2(n54872), .A(n54667), .ZN(n54668) );
  AOI21_X1 U37289 ( .B1(\DP/ALU0/s_A_MULT[11] ), .B2(n54693), .A(n54668), .ZN(
        \intadd_2/A[11] ) );
  AOI22_X1 U37290 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54687), .B1(
        \DP/ALU0/s_A_MULT[12] ), .B2(n54693), .ZN(n54669) );
  OAI21_X1 U37291 ( .B1(n54876), .B2(n54690), .A(n54669), .ZN(n54670) );
  AOI21_X1 U37292 ( .B1(n53644), .B2(n54874), .A(n54670), .ZN(\intadd_2/A[12] ) );
  AOI22_X1 U37293 ( .A1(\DP/ALU0/s_A_MULT[2] ), .A2(n54687), .B1(
        \DP/ALU0/s_A_MULT[1] ), .B2(n54693), .ZN(n54671) );
  OAI21_X1 U37294 ( .B1(n54690), .B2(n54879), .A(n54671), .ZN(n54672) );
  AOI21_X1 U37295 ( .B1(n53644), .B2(n54881), .A(n54672), .ZN(\intadd_2/A[1] )
         );
  AOI22_X1 U37296 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n54687), .B1(
        \DP/ALU0/s_A_MULT[2] ), .B2(n54693), .ZN(n54673) );
  OAI21_X1 U37297 ( .B1(n54690), .B2(n54883), .A(n54673), .ZN(n54674) );
  AOI21_X1 U37298 ( .B1(n53644), .B2(n54885), .A(n54674), .ZN(\intadd_2/A[2] )
         );
  AOI22_X1 U37299 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54687), .B1(n53644), .B2(
        n54886), .ZN(n54675) );
  OAI21_X1 U37300 ( .B1(n54690), .B2(n54888), .A(n54675), .ZN(n54676) );
  AOI21_X1 U37301 ( .B1(\DP/ALU0/s_A_MULT[3] ), .B2(n54693), .A(n54676), .ZN(
        \intadd_2/A[3] ) );
  AOI22_X1 U37302 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54693), .B1(n53644), .B2(
        n54890), .ZN(n54677) );
  OAI21_X1 U37303 ( .B1(n54690), .B2(n54892), .A(n54677), .ZN(n54678) );
  AOI21_X1 U37304 ( .B1(\DP/ALU0/s_A_MULT[5] ), .B2(n54687), .A(n54678), .ZN(
        \intadd_2/A[4] ) );
  AOI22_X1 U37305 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54687), .B1(n53644), .B2(
        n54894), .ZN(n54679) );
  OAI21_X1 U37306 ( .B1(n54690), .B2(n54896), .A(n54679), .ZN(n54680) );
  AOI21_X1 U37307 ( .B1(\DP/ALU0/s_A_MULT[5] ), .B2(n54693), .A(n54680), .ZN(
        \intadd_2/A[5] ) );
  AOI22_X1 U37308 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54693), .B1(n53644), .B2(
        n54898), .ZN(n54681) );
  OAI21_X1 U37309 ( .B1(n54690), .B2(n54900), .A(n54681), .ZN(n54682) );
  AOI21_X1 U37310 ( .B1(\DP/ALU0/s_A_MULT[7] ), .B2(n54687), .A(n54682), .ZN(
        \intadd_2/A[6] ) );
  AOI22_X1 U37311 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54687), .B1(n53644), .B2(
        n54902), .ZN(n54683) );
  OAI21_X1 U37312 ( .B1(n54690), .B2(n54904), .A(n54683), .ZN(n54684) );
  AOI21_X1 U37313 ( .B1(\DP/ALU0/s_A_MULT[7] ), .B2(n54693), .A(n54684), .ZN(
        \intadd_2/A[7] ) );
  AOI22_X1 U37314 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54693), .B1(n53644), .B2(
        n54906), .ZN(n54685) );
  OAI21_X1 U37315 ( .B1(n54690), .B2(n54908), .A(n54685), .ZN(n54686) );
  AOI21_X1 U37316 ( .B1(\DP/ALU0/s_A_MULT[9] ), .B2(n54687), .A(n54686), .ZN(
        \intadd_2/A[8] ) );
  AOI22_X1 U37317 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n54687), .B1(
        \DP/ALU0/s_A_MULT[9] ), .B2(n54693), .ZN(n54688) );
  OAI21_X1 U37318 ( .B1(n54690), .B2(n54912), .A(n54688), .ZN(n54689) );
  AOI21_X1 U37319 ( .B1(n53644), .B2(n54914), .A(n54689), .ZN(\intadd_2/A[9] )
         );
  OAI22_X1 U37320 ( .A1(n54918), .A2(n54691), .B1(n54690), .B2(n54915), .ZN(
        n54692) );
  AOI221_X1 U37321 ( .B1(n53644), .B2(\DP/ALU0/s_A_MULT[0] ), .C1(n54693), 
        .C2(\DP/ALU0/s_A_MULT[0] ), .A(n54692), .ZN(\intadd_2/B[0] ) );
  OAI21_X1 U37322 ( .B1(\intadd_3/n1 ), .B2(n54696), .A(n54695), .ZN(n54698)
         );
  XNOR2_X1 U37323 ( .A(n54698), .B(n54697), .ZN(\intadd_2/B[11] ) );
  INV_X1 U37324 ( .A(n54699), .ZN(n54700) );
  NOR2_X1 U37325 ( .A1(n54701), .A2(n54700), .ZN(n54702) );
  XNOR2_X1 U37326 ( .A(n54703), .B(n54702), .ZN(\intadd_2/B[12] ) );
  AOI22_X1 U37327 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n54728), .B1(
        \DP/ALU0/s_A_MULT[10] ), .B2(n54732), .ZN(n54704) );
  OAI21_X1 U37328 ( .B1(n54729), .B2(n54867), .A(n54704), .ZN(n54705) );
  AOI21_X1 U37329 ( .B1(n54733), .B2(n54869), .A(n54705), .ZN(\intadd_3/A[10] ) );
  AOI22_X1 U37330 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n54732), .B1(n54733), 
        .B2(n54870), .ZN(n54706) );
  OAI21_X1 U37331 ( .B1(n54729), .B2(n54872), .A(n54706), .ZN(n54707) );
  AOI21_X1 U37332 ( .B1(\DP/ALU0/s_A_MULT[12] ), .B2(n54728), .A(n54707), .ZN(
        \intadd_3/A[11] ) );
  AOI22_X1 U37333 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54728), .B1(n54733), 
        .B2(n54874), .ZN(n54708) );
  OAI21_X1 U37334 ( .B1(n54876), .B2(n54729), .A(n54708), .ZN(n54709) );
  AOI21_X1 U37335 ( .B1(\DP/ALU0/s_A_MULT[12] ), .B2(n54732), .A(n54709), .ZN(
        \intadd_3/A[12] ) );
  AOI22_X1 U37336 ( .A1(\DP/ALU0/s_A_MULT[2] ), .A2(n54728), .B1(
        \DP/ALU0/s_A_MULT[1] ), .B2(n54732), .ZN(n54710) );
  OAI21_X1 U37337 ( .B1(n54729), .B2(n54879), .A(n54710), .ZN(n54711) );
  AOI21_X1 U37338 ( .B1(n54733), .B2(n54881), .A(n54711), .ZN(\intadd_3/A[1] )
         );
  AOI22_X1 U37339 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n54728), .B1(
        \DP/ALU0/s_A_MULT[2] ), .B2(n54732), .ZN(n54712) );
  OAI21_X1 U37340 ( .B1(n54729), .B2(n54883), .A(n54712), .ZN(n54713) );
  AOI21_X1 U37341 ( .B1(n54733), .B2(n54885), .A(n54713), .ZN(\intadd_3/A[2] )
         );
  AOI22_X1 U37342 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n54732), .B1(n54733), .B2(
        n54886), .ZN(n54714) );
  OAI21_X1 U37343 ( .B1(n54729), .B2(n54888), .A(n54714), .ZN(n54715) );
  AOI21_X1 U37344 ( .B1(\DP/ALU0/s_A_MULT[4] ), .B2(n54728), .A(n54715), .ZN(
        \intadd_3/A[3] ) );
  AOI22_X1 U37345 ( .A1(\DP/ALU0/s_A_MULT[5] ), .A2(n54728), .B1(n54733), .B2(
        n54890), .ZN(n54716) );
  OAI21_X1 U37346 ( .B1(n54729), .B2(n54892), .A(n54716), .ZN(n54717) );
  AOI21_X1 U37347 ( .B1(\DP/ALU0/s_A_MULT[4] ), .B2(n54732), .A(n54717), .ZN(
        \intadd_3/A[4] ) );
  AOI22_X1 U37348 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54728), .B1(n54733), .B2(
        n54894), .ZN(n54718) );
  OAI21_X1 U37349 ( .B1(n54729), .B2(n54896), .A(n54718), .ZN(n54719) );
  AOI21_X1 U37350 ( .B1(\DP/ALU0/s_A_MULT[5] ), .B2(n54732), .A(n54719), .ZN(
        \intadd_3/A[5] ) );
  AOI22_X1 U37351 ( .A1(\DP/ALU0/s_A_MULT[7] ), .A2(n54728), .B1(n54733), .B2(
        n54898), .ZN(n54720) );
  OAI21_X1 U37352 ( .B1(n54729), .B2(n54900), .A(n54720), .ZN(n54721) );
  AOI21_X1 U37353 ( .B1(\DP/ALU0/s_A_MULT[6] ), .B2(n54732), .A(n54721), .ZN(
        \intadd_3/A[6] ) );
  AOI22_X1 U37354 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54728), .B1(n54733), .B2(
        n54902), .ZN(n54722) );
  OAI21_X1 U37355 ( .B1(n54729), .B2(n54904), .A(n54722), .ZN(n54723) );
  AOI21_X1 U37356 ( .B1(\DP/ALU0/s_A_MULT[7] ), .B2(n54732), .A(n54723), .ZN(
        \intadd_3/A[7] ) );
  AOI22_X1 U37357 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54732), .B1(n54733), .B2(
        n54906), .ZN(n54724) );
  OAI21_X1 U37358 ( .B1(n54729), .B2(n54908), .A(n54724), .ZN(n54725) );
  AOI21_X1 U37359 ( .B1(\DP/ALU0/s_A_MULT[9] ), .B2(n54728), .A(n54725), .ZN(
        \intadd_3/A[8] ) );
  AOI22_X1 U37360 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n54728), .B1(
        \DP/ALU0/s_A_MULT[9] ), .B2(n54732), .ZN(n54726) );
  OAI21_X1 U37361 ( .B1(n54729), .B2(n54912), .A(n54726), .ZN(n54727) );
  AOI21_X1 U37362 ( .B1(n54733), .B2(n54914), .A(n54727), .ZN(\intadd_3/A[9] )
         );
  INV_X1 U37363 ( .A(n54728), .ZN(n54730) );
  OAI22_X1 U37364 ( .A1(n54918), .A2(n54730), .B1(n54729), .B2(n54915), .ZN(
        n54731) );
  AOI221_X1 U37365 ( .B1(n54733), .B2(\DP/ALU0/s_A_MULT[0] ), .C1(n54732), 
        .C2(\DP/ALU0/s_A_MULT[0] ), .A(n54731), .ZN(\intadd_3/B[0] ) );
  INV_X1 U37366 ( .A(n54735), .ZN(n54734) );
  AOI22_X1 U37367 ( .A1(n54736), .A2(n54735), .B1(n54734), .B2(n54740), .ZN(
        n54737) );
  XNOR2_X1 U37368 ( .A(\intadd_4/n1 ), .B(n54737), .ZN(\intadd_3/B[11] ) );
  INV_X1 U37369 ( .A(\intadd_4/n1 ), .ZN(n54739) );
  OAI21_X1 U37370 ( .B1(n54740), .B2(n54739), .A(n54738), .ZN(n54742) );
  XNOR2_X1 U37371 ( .A(n54742), .B(n54741), .ZN(\intadd_3/B[12] ) );
  INV_X1 U37372 ( .A(n54744), .ZN(n54748) );
  INV_X1 U37373 ( .A(n54745), .ZN(n54743) );
  AOI22_X1 U37374 ( .A1(n54745), .A2(n54748), .B1(n54744), .B2(n54743), .ZN(
        n54746) );
  XNOR2_X1 U37375 ( .A(\intadd_5/n1 ), .B(n54746), .ZN(\intadd_4/A[11] ) );
  OAI21_X1 U37376 ( .B1(n54748), .B2(\intadd_5/n1 ), .A(n54747), .ZN(n54750)
         );
  XNOR2_X1 U37377 ( .A(n54750), .B(n54749), .ZN(\intadd_4/A[12] ) );
  AOI22_X1 U37378 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n54777), .B1(
        \DP/ALU0/s_A_MULT[10] ), .B2(n54775), .ZN(n54752) );
  NAND2_X1 U37379 ( .A1(n53640), .A2(n54869), .ZN(n54751) );
  OAI211_X1 U37380 ( .C1(n54867), .C2(n54780), .A(n54752), .B(n54751), .ZN(
        \intadd_4/B[10] ) );
  AOI22_X1 U37381 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n54777), .B1(n53640), 
        .B2(n54870), .ZN(n54754) );
  NAND2_X1 U37382 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n54775), .ZN(n54753) );
  OAI211_X1 U37383 ( .C1(n54872), .C2(n54780), .A(n54754), .B(n54753), .ZN(
        \intadd_4/B[11] ) );
  AOI22_X1 U37384 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54777), .B1(
        \DP/ALU0/s_A_MULT[12] ), .B2(n54775), .ZN(n54756) );
  NAND2_X1 U37385 ( .A1(n53640), .A2(n54874), .ZN(n54755) );
  OAI211_X1 U37386 ( .C1(n54780), .C2(n54876), .A(n54756), .B(n54755), .ZN(
        \intadd_4/B[12] ) );
  AOI22_X1 U37387 ( .A1(\DP/ALU0/s_A_MULT[2] ), .A2(n54777), .B1(
        \DP/ALU0/s_A_MULT[1] ), .B2(n54775), .ZN(n54758) );
  NAND2_X1 U37388 ( .A1(n53640), .A2(n54881), .ZN(n54757) );
  OAI211_X1 U37389 ( .C1(n54879), .C2(n54780), .A(n54758), .B(n54757), .ZN(
        \intadd_4/B[1] ) );
  AOI22_X1 U37390 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n54777), .B1(
        \DP/ALU0/s_A_MULT[2] ), .B2(n54775), .ZN(n54760) );
  NAND2_X1 U37391 ( .A1(n53640), .A2(n54885), .ZN(n54759) );
  OAI211_X1 U37392 ( .C1(n54883), .C2(n54780), .A(n54760), .B(n54759), .ZN(
        \intadd_4/B[2] ) );
  AOI22_X1 U37393 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54777), .B1(n53640), .B2(
        n54886), .ZN(n54762) );
  NAND2_X1 U37394 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n54775), .ZN(n54761) );
  OAI211_X1 U37395 ( .C1(n54888), .C2(n54780), .A(n54762), .B(n54761), .ZN(
        \intadd_4/B[3] ) );
  AOI22_X1 U37396 ( .A1(\DP/ALU0/s_A_MULT[5] ), .A2(n54777), .B1(n53640), .B2(
        n54890), .ZN(n54764) );
  NAND2_X1 U37397 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54775), .ZN(n54763) );
  OAI211_X1 U37398 ( .C1(n54892), .C2(n54780), .A(n54764), .B(n54763), .ZN(
        \intadd_4/B[4] ) );
  AOI22_X1 U37399 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54777), .B1(n53640), .B2(
        n54894), .ZN(n54766) );
  NAND2_X1 U37400 ( .A1(\DP/ALU0/s_A_MULT[5] ), .A2(n54775), .ZN(n54765) );
  OAI211_X1 U37401 ( .C1(n54896), .C2(n54780), .A(n54766), .B(n54765), .ZN(
        \intadd_4/B[5] ) );
  AOI22_X1 U37402 ( .A1(\DP/ALU0/s_A_MULT[7] ), .A2(n54777), .B1(n53640), .B2(
        n54898), .ZN(n54768) );
  NAND2_X1 U37403 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54775), .ZN(n54767) );
  OAI211_X1 U37404 ( .C1(n54900), .C2(n54780), .A(n54768), .B(n54767), .ZN(
        \intadd_4/B[6] ) );
  AOI22_X1 U37405 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54777), .B1(n53640), .B2(
        n54902), .ZN(n54770) );
  NAND2_X1 U37406 ( .A1(\DP/ALU0/s_A_MULT[7] ), .A2(n54775), .ZN(n54769) );
  OAI211_X1 U37407 ( .C1(n54904), .C2(n54780), .A(n54770), .B(n54769), .ZN(
        \intadd_4/B[7] ) );
  AOI22_X1 U37408 ( .A1(\DP/ALU0/s_A_MULT[9] ), .A2(n54777), .B1(n53640), .B2(
        n54906), .ZN(n54772) );
  NAND2_X1 U37409 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54775), .ZN(n54771) );
  OAI211_X1 U37410 ( .C1(n54908), .C2(n54780), .A(n54772), .B(n54771), .ZN(
        \intadd_4/B[8] ) );
  AOI22_X1 U37411 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n54777), .B1(
        \DP/ALU0/s_A_MULT[9] ), .B2(n54775), .ZN(n54774) );
  NAND2_X1 U37412 ( .A1(n53640), .A2(n54914), .ZN(n54773) );
  OAI211_X1 U37413 ( .C1(n54912), .C2(n54780), .A(n54774), .B(n54773), .ZN(
        \intadd_4/B[9] ) );
  NOR2_X1 U37414 ( .A1(n53640), .A2(n54775), .ZN(n54779) );
  INV_X1 U37415 ( .A(n54777), .ZN(n54778) );
  OAI222_X1 U37416 ( .A1(n54915), .A2(n54780), .B1(n55299), .B2(n54779), .C1(
        n54918), .C2(n54778), .ZN(\intadd_4/CI ) );
  AOI22_X1 U37417 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n54803), .B1(
        \DP/ALU0/s_A_MULT[10] ), .B2(n54809), .ZN(n54781) );
  OAI21_X1 U37418 ( .B1(n54806), .B2(n54867), .A(n54781), .ZN(n54782) );
  AOI21_X1 U37419 ( .B1(n53641), .B2(n54869), .A(n54782), .ZN(\intadd_5/A[10] ) );
  AOI22_X1 U37420 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n54803), .B1(n53641), 
        .B2(n54870), .ZN(n54783) );
  OAI21_X1 U37421 ( .B1(n54806), .B2(n54872), .A(n54783), .ZN(n54784) );
  AOI21_X1 U37422 ( .B1(\DP/ALU0/s_A_MULT[11] ), .B2(n54809), .A(n54784), .ZN(
        \intadd_5/A[11] ) );
  AOI22_X1 U37423 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n54809), .B1(n53641), 
        .B2(n54874), .ZN(n54785) );
  OAI21_X1 U37424 ( .B1(n54876), .B2(n54806), .A(n54785), .ZN(n54786) );
  AOI21_X1 U37425 ( .B1(\DP/ALU0/s_A_MULT[13] ), .B2(n54803), .A(n54786), .ZN(
        \intadd_5/A[12] ) );
  AOI22_X1 U37426 ( .A1(\DP/ALU0/s_A_MULT[2] ), .A2(n54803), .B1(
        \DP/ALU0/s_A_MULT[1] ), .B2(n54809), .ZN(n54787) );
  OAI21_X1 U37427 ( .B1(n54806), .B2(n54879), .A(n54787), .ZN(n54788) );
  AOI21_X1 U37428 ( .B1(n53641), .B2(n54881), .A(n54788), .ZN(\intadd_5/A[1] )
         );
  AOI22_X1 U37429 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n54803), .B1(
        \DP/ALU0/s_A_MULT[2] ), .B2(n54809), .ZN(n54789) );
  OAI21_X1 U37430 ( .B1(n54806), .B2(n54883), .A(n54789), .ZN(n54790) );
  AOI21_X1 U37431 ( .B1(n53641), .B2(n54885), .A(n54790), .ZN(\intadd_5/A[2] )
         );
  AOI22_X1 U37432 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54803), .B1(n53641), .B2(
        n54886), .ZN(n54791) );
  OAI21_X1 U37433 ( .B1(n54806), .B2(n54888), .A(n54791), .ZN(n54792) );
  AOI21_X1 U37434 ( .B1(\DP/ALU0/s_A_MULT[3] ), .B2(n54809), .A(n54792), .ZN(
        \intadd_5/A[3] ) );
  AOI22_X1 U37435 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54809), .B1(n53641), .B2(
        n54890), .ZN(n54793) );
  OAI21_X1 U37436 ( .B1(n54806), .B2(n54892), .A(n54793), .ZN(n54794) );
  AOI21_X1 U37437 ( .B1(\DP/ALU0/s_A_MULT[5] ), .B2(n54803), .A(n54794), .ZN(
        \intadd_5/A[4] ) );
  AOI22_X1 U37438 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54803), .B1(n53641), .B2(
        n54894), .ZN(n54795) );
  OAI21_X1 U37439 ( .B1(n54806), .B2(n54896), .A(n54795), .ZN(n54796) );
  AOI21_X1 U37440 ( .B1(\DP/ALU0/s_A_MULT[5] ), .B2(n54809), .A(n54796), .ZN(
        \intadd_5/A[5] ) );
  AOI22_X1 U37441 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54809), .B1(n53641), .B2(
        n54898), .ZN(n54797) );
  OAI21_X1 U37442 ( .B1(n54806), .B2(n54900), .A(n54797), .ZN(n54798) );
  AOI21_X1 U37443 ( .B1(\DP/ALU0/s_A_MULT[7] ), .B2(n54803), .A(n54798), .ZN(
        \intadd_5/A[6] ) );
  AOI22_X1 U37444 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54803), .B1(n53641), .B2(
        n54902), .ZN(n54799) );
  OAI21_X1 U37445 ( .B1(n54806), .B2(n54904), .A(n54799), .ZN(n54800) );
  AOI21_X1 U37446 ( .B1(\DP/ALU0/s_A_MULT[7] ), .B2(n54809), .A(n54800), .ZN(
        \intadd_5/A[7] ) );
  AOI22_X1 U37447 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54809), .B1(n53641), .B2(
        n54906), .ZN(n54801) );
  OAI21_X1 U37448 ( .B1(n54806), .B2(n54908), .A(n54801), .ZN(n54802) );
  AOI21_X1 U37449 ( .B1(\DP/ALU0/s_A_MULT[9] ), .B2(n54803), .A(n54802), .ZN(
        \intadd_5/A[8] ) );
  AOI22_X1 U37450 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n54803), .B1(n53641), 
        .B2(n54914), .ZN(n54804) );
  OAI21_X1 U37451 ( .B1(n54806), .B2(n54912), .A(n54804), .ZN(n54805) );
  AOI21_X1 U37452 ( .B1(\DP/ALU0/s_A_MULT[9] ), .B2(n54809), .A(n54805), .ZN(
        \intadd_5/A[9] ) );
  OAI22_X1 U37453 ( .A1(n54918), .A2(n54807), .B1(n54806), .B2(n54915), .ZN(
        n54808) );
  AOI221_X1 U37454 ( .B1(n53641), .B2(\DP/ALU0/s_A_MULT[0] ), .C1(n54809), 
        .C2(\DP/ALU0/s_A_MULT[0] ), .A(n54808), .ZN(\intadd_5/B[0] ) );
  INV_X1 U37455 ( .A(n54811), .ZN(n54812) );
  NOR2_X1 U37456 ( .A1(n54813), .A2(n54812), .ZN(n54814) );
  XNOR2_X1 U37457 ( .A(n54815), .B(n54814), .ZN(\intadd_5/B[12] ) );
  NOR3_X1 U37458 ( .A1(\intadd_7/SUM[1] ), .A2(n55298), .A3(n55299), .ZN(
        \intadd_6/A[0] ) );
  AOI21_X1 U37459 ( .B1(n54819), .B2(n54817), .A(n54816), .ZN(n54818) );
  XOR2_X1 U37460 ( .A(\intadd_7/n1 ), .B(n54818), .Z(\intadd_6/A[11] ) );
  INV_X1 U37461 ( .A(n54819), .ZN(n54821) );
  AOI21_X1 U37462 ( .B1(\intadd_7/n1 ), .B2(n54821), .A(n54820), .ZN(n54823)
         );
  XOR2_X1 U37463 ( .A(n54823), .B(n54822), .Z(\intadd_6/A[12] ) );
  AOI22_X1 U37464 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n54849), .B1(n54850), 
        .B2(n54870), .ZN(n54825) );
  AOI22_X1 U37465 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n54851), .B1(n53639), 
        .B2(n54869), .ZN(n54824) );
  NAND2_X1 U37466 ( .A1(n54825), .A2(n54824), .ZN(\intadd_6/B[10] ) );
  AOI22_X1 U37467 ( .A1(n53639), .A2(n54870), .B1(n54850), .B2(n54874), .ZN(
        n54827) );
  AOI22_X1 U37468 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n54851), .B1(
        \DP/ALU0/s_A_MULT[11] ), .B2(n54849), .ZN(n54826) );
  NAND2_X1 U37469 ( .A1(n54827), .A2(n54826), .ZN(\intadd_6/B[11] ) );
  AOI22_X1 U37470 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54851), .B1(n53639), 
        .B2(n54874), .ZN(n54829) );
  AOI22_X1 U37471 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n54849), .B1(n54856), 
        .B2(n54850), .ZN(n54828) );
  NAND2_X1 U37472 ( .A1(n54829), .A2(n54828), .ZN(\intadd_6/B[12] ) );
  AOI22_X1 U37473 ( .A1(\DP/ALU0/s_A_MULT[2] ), .A2(n54851), .B1(
        \DP/ALU0/s_A_MULT[1] ), .B2(n54849), .ZN(n54831) );
  AOI22_X1 U37474 ( .A1(n53639), .A2(n54881), .B1(n54850), .B2(n54885), .ZN(
        n54830) );
  NAND2_X1 U37475 ( .A1(n54831), .A2(n54830), .ZN(\intadd_6/B[1] ) );
  AOI22_X1 U37476 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n54851), .B1(
        \DP/ALU0/s_A_MULT[2] ), .B2(n54849), .ZN(n54833) );
  AOI22_X1 U37477 ( .A1(n53639), .A2(n54885), .B1(n54850), .B2(n54886), .ZN(
        n54832) );
  NAND2_X1 U37478 ( .A1(n54833), .A2(n54832), .ZN(\intadd_6/B[2] ) );
  AOI22_X1 U37479 ( .A1(n53639), .A2(n54886), .B1(n54850), .B2(n54890), .ZN(
        n54835) );
  AOI22_X1 U37480 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54851), .B1(
        \DP/ALU0/s_A_MULT[3] ), .B2(n54849), .ZN(n54834) );
  NAND2_X1 U37481 ( .A1(n54835), .A2(n54834), .ZN(\intadd_6/B[3] ) );
  AOI22_X1 U37482 ( .A1(n53639), .A2(n54890), .B1(n54850), .B2(n54894), .ZN(
        n54837) );
  AOI22_X1 U37483 ( .A1(\DP/ALU0/s_A_MULT[5] ), .A2(n54851), .B1(
        \DP/ALU0/s_A_MULT[4] ), .B2(n54849), .ZN(n54836) );
  NAND2_X1 U37484 ( .A1(n54837), .A2(n54836), .ZN(\intadd_6/B[4] ) );
  AOI22_X1 U37485 ( .A1(n53639), .A2(n54894), .B1(n54850), .B2(n54898), .ZN(
        n54839) );
  AOI22_X1 U37486 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54851), .B1(
        \DP/ALU0/s_A_MULT[5] ), .B2(n54849), .ZN(n54838) );
  NAND2_X1 U37487 ( .A1(n54839), .A2(n54838), .ZN(\intadd_6/B[5] ) );
  AOI22_X1 U37488 ( .A1(n53639), .A2(n54898), .B1(n54850), .B2(n54902), .ZN(
        n54841) );
  AOI22_X1 U37489 ( .A1(\DP/ALU0/s_A_MULT[7] ), .A2(n54851), .B1(
        \DP/ALU0/s_A_MULT[6] ), .B2(n54849), .ZN(n54840) );
  NAND2_X1 U37490 ( .A1(n54841), .A2(n54840), .ZN(\intadd_6/B[6] ) );
  AOI22_X1 U37491 ( .A1(n53639), .A2(n54902), .B1(n54850), .B2(n54906), .ZN(
        n54843) );
  AOI22_X1 U37492 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54851), .B1(
        \DP/ALU0/s_A_MULT[7] ), .B2(n54849), .ZN(n54842) );
  NAND2_X1 U37493 ( .A1(n54843), .A2(n54842), .ZN(\intadd_6/B[7] ) );
  AOI22_X1 U37494 ( .A1(n53639), .A2(n54906), .B1(n54850), .B2(n54914), .ZN(
        n54845) );
  AOI22_X1 U37495 ( .A1(\DP/ALU0/s_A_MULT[9] ), .A2(n54851), .B1(
        \DP/ALU0/s_A_MULT[8] ), .B2(n54849), .ZN(n54844) );
  NAND2_X1 U37496 ( .A1(n54845), .A2(n54844), .ZN(\intadd_6/B[8] ) );
  AOI22_X1 U37497 ( .A1(\DP/ALU0/s_A_MULT[9] ), .A2(n54849), .B1(n54850), .B2(
        n54869), .ZN(n54848) );
  AOI22_X1 U37498 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n54851), .B1(n53639), 
        .B2(n54914), .ZN(n54847) );
  NAND2_X1 U37499 ( .A1(n54848), .A2(n54847), .ZN(\intadd_6/B[9] ) );
  INV_X1 U37500 ( .A(n54849), .ZN(n54853) );
  AOI22_X1 U37501 ( .A1(\DP/ALU0/s_A_MULT[1] ), .A2(n54851), .B1(n54850), .B2(
        n54881), .ZN(n54852) );
  OAI221_X1 U37502 ( .B1(n55299), .B2(n54846), .C1(n55299), .C2(n54853), .A(
        n54852), .ZN(\intadd_6/CI ) );
  NOR2_X1 U37503 ( .A1(n54854), .A2(n54872), .ZN(n54855) );
  OAI222_X1 U37504 ( .A1(n54859), .A2(n54856), .B1(\DP/ALU0/s_A_MULT[13] ), 
        .B2(\DP/ALU0/S_B_MULT[1] ), .C1(n54855), .C2(\DP/ALU0/S_B_MULT[0] ), 
        .ZN(\intadd_7/A[10] ) );
  AOI222_X1 U37505 ( .A1(\DP/ALU0/s_A_MULT[14] ), .A2(n54865), .B1(n54862), 
        .B2(n54863), .C1(n54856), .C2(n54864), .ZN(\intadd_7/A[11] ) );
  OAI22_X1 U37506 ( .A1(n54860), .A2(n54859), .B1(n54858), .B2(n54857), .ZN(
        n54861) );
  AOI21_X1 U37507 ( .B1(n54862), .B2(n54864), .A(n54861), .ZN(\intadd_7/A[12] ) );
  AOI222_X1 U37508 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54865), .B1(n54864), 
        .B2(n54886), .C1(n54863), .C2(n54890), .ZN(\intadd_7/A[1] ) );
  AOI222_X1 U37509 ( .A1(\DP/ALU0/s_A_MULT[5] ), .A2(n54865), .B1(n54864), 
        .B2(n54890), .C1(n54863), .C2(n54894), .ZN(\intadd_7/A[2] ) );
  AOI222_X1 U37510 ( .A1(\DP/ALU0/s_A_MULT[6] ), .A2(n54865), .B1(n54864), 
        .B2(n54894), .C1(n54863), .C2(n54898), .ZN(\intadd_7/A[3] ) );
  AOI222_X1 U37511 ( .A1(\DP/ALU0/s_A_MULT[7] ), .A2(n54865), .B1(n54864), 
        .B2(n54898), .C1(n54863), .C2(n54902), .ZN(\intadd_7/A[4] ) );
  AOI222_X1 U37512 ( .A1(\DP/ALU0/s_A_MULT[8] ), .A2(n54865), .B1(n54864), 
        .B2(n54902), .C1(n54863), .C2(n54906), .ZN(\intadd_7/A[5] ) );
  AOI222_X1 U37513 ( .A1(\DP/ALU0/s_A_MULT[9] ), .A2(n54865), .B1(n54864), 
        .B2(n54906), .C1(n54863), .C2(n54914), .ZN(\intadd_7/A[6] ) );
  AOI222_X1 U37514 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n54865), .B1(n54864), 
        .B2(n54914), .C1(n54863), .C2(n54869), .ZN(\intadd_7/A[7] ) );
  AOI222_X1 U37515 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n54865), .B1(n54864), 
        .B2(n54869), .C1(n54863), .C2(n54870), .ZN(\intadd_7/A[8] ) );
  AOI222_X1 U37516 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n54865), .B1(n54864), 
        .B2(n54870), .C1(n54863), .C2(n54874), .ZN(\intadd_7/A[9] ) );
  AOI222_X1 U37517 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n54865), .B1(n54864), 
        .B2(n54885), .C1(n54863), .C2(n54886), .ZN(\intadd_7/B[0] ) );
  AOI22_X1 U37518 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n54910), .B1(
        \DP/ALU0/s_A_MULT[10] ), .B2(n54920), .ZN(n54866) );
  OAI21_X1 U37519 ( .B1(n54916), .B2(n54867), .A(n54866), .ZN(n54868) );
  AOI21_X1 U37520 ( .B1(n53643), .B2(n54869), .A(n54868), .ZN(\intadd_7/B[10] ) );
  AOI22_X1 U37521 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n54910), .B1(n53643), 
        .B2(n54870), .ZN(n54871) );
  OAI21_X1 U37522 ( .B1(n54916), .B2(n54872), .A(n54871), .ZN(n54873) );
  AOI21_X1 U37523 ( .B1(\DP/ALU0/s_A_MULT[11] ), .B2(n54920), .A(n54873), .ZN(
        \intadd_7/B[11] ) );
  AOI22_X1 U37524 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n54910), .B1(n53643), 
        .B2(n54874), .ZN(n54875) );
  OAI21_X1 U37525 ( .B1(n54876), .B2(n54916), .A(n54875), .ZN(n54877) );
  AOI21_X1 U37526 ( .B1(\DP/ALU0/s_A_MULT[12] ), .B2(n54920), .A(n54877), .ZN(
        \intadd_7/B[12] ) );
  AOI22_X1 U37527 ( .A1(\DP/ALU0/s_A_MULT[2] ), .A2(n54910), .B1(
        \DP/ALU0/s_A_MULT[1] ), .B2(n54920), .ZN(n54878) );
  OAI21_X1 U37528 ( .B1(n54916), .B2(n54879), .A(n54878), .ZN(n54880) );
  AOI21_X1 U37529 ( .B1(n53643), .B2(n54881), .A(n54880), .ZN(\intadd_7/B[1] )
         );
  AOI22_X1 U37530 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n54910), .B1(
        \DP/ALU0/s_A_MULT[2] ), .B2(n54920), .ZN(n54882) );
  OAI21_X1 U37531 ( .B1(n54916), .B2(n54883), .A(n54882), .ZN(n54884) );
  AOI21_X1 U37532 ( .B1(n53643), .B2(n54885), .A(n54884), .ZN(\intadd_7/B[2] )
         );
  AOI22_X1 U37533 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n54910), .B1(n53643), .B2(
        n54886), .ZN(n54887) );
  OAI21_X1 U37534 ( .B1(n54916), .B2(n54888), .A(n54887), .ZN(n54889) );
  AOI21_X1 U37535 ( .B1(\DP/ALU0/s_A_MULT[3] ), .B2(n54920), .A(n54889), .ZN(
        \intadd_7/B[3] ) );
  AOI22_X1 U37536 ( .A1(\DP/ALU0/s_A_MULT[5] ), .A2(n54910), .B1(n53643), .B2(
        n54890), .ZN(n54891) );
  OAI21_X1 U37537 ( .B1(n54916), .B2(n54892), .A(n54891), .ZN(n54893) );
  AOI21_X1 U37538 ( .B1(\DP/ALU0/s_A_MULT[4] ), .B2(n54920), .A(n54893), .ZN(
        \intadd_7/B[4] ) );
  AOI22_X1 U37539 ( .A1(\DP/ALU0/s_A_MULT[5] ), .A2(n54920), .B1(n53643), .B2(
        n54894), .ZN(n54895) );
  OAI21_X1 U37540 ( .B1(n54916), .B2(n54896), .A(n54895), .ZN(n54897) );
  AOI21_X1 U37541 ( .B1(\DP/ALU0/s_A_MULT[6] ), .B2(n54910), .A(n54897), .ZN(
        \intadd_7/B[5] ) );
  AOI22_X1 U37542 ( .A1(\DP/ALU0/s_A_MULT[7] ), .A2(n54910), .B1(n53643), .B2(
        n54898), .ZN(n54899) );
  OAI21_X1 U37543 ( .B1(n54916), .B2(n54900), .A(n54899), .ZN(n54901) );
  AOI21_X1 U37544 ( .B1(\DP/ALU0/s_A_MULT[6] ), .B2(n54920), .A(n54901), .ZN(
        \intadd_7/B[6] ) );
  AOI22_X1 U37545 ( .A1(\DP/ALU0/s_A_MULT[7] ), .A2(n54920), .B1(n53643), .B2(
        n54902), .ZN(n54903) );
  OAI21_X1 U37546 ( .B1(n54916), .B2(n54904), .A(n54903), .ZN(n54905) );
  AOI21_X1 U37547 ( .B1(\DP/ALU0/s_A_MULT[8] ), .B2(n54910), .A(n54905), .ZN(
        \intadd_7/B[7] ) );
  AOI22_X1 U37548 ( .A1(\DP/ALU0/s_A_MULT[9] ), .A2(n54910), .B1(n53643), .B2(
        n54906), .ZN(n54907) );
  OAI21_X1 U37549 ( .B1(n54916), .B2(n54908), .A(n54907), .ZN(n54909) );
  AOI21_X1 U37550 ( .B1(\DP/ALU0/s_A_MULT[8] ), .B2(n54920), .A(n54909), .ZN(
        \intadd_7/B[8] ) );
  AOI22_X1 U37551 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n54910), .B1(
        \DP/ALU0/s_A_MULT[9] ), .B2(n54920), .ZN(n54911) );
  OAI21_X1 U37552 ( .B1(n54916), .B2(n54912), .A(n54911), .ZN(n54913) );
  AOI21_X1 U37553 ( .B1(n53643), .B2(n54914), .A(n54913), .ZN(\intadd_7/B[9] )
         );
  OAI22_X1 U37554 ( .A1(n54918), .A2(n54917), .B1(n54916), .B2(n54915), .ZN(
        n54919) );
  AOI221_X1 U37555 ( .B1(n53643), .B2(\DP/ALU0/s_A_MULT[0] ), .C1(n54920), 
        .C2(\DP/ALU0/s_A_MULT[0] ), .A(n54919), .ZN(\intadd_7/CI ) );
  XNOR2_X1 U37556 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[29] ), .ZN(
        \intadd_8/B[1] ) );
  XNOR2_X1 U37557 ( .A(\DP/ALU0/s_ADD_SUB ), .B(\DP/ALU0/S_B_ADDER[30] ), .ZN(
        \intadd_8/B[2] ) );
  XNOR2_X1 U37558 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[31] ), .ZN(
        \intadd_8/B[3] ) );
  XNOR2_X1 U37559 ( .A(n53817), .B(\DP/ALU0/S_B_ADDER[28] ), .ZN(\intadd_8/CI ) );
  NOR2_X1 U37560 ( .A1(n45959), .A2(n53812), .ZN(n55290) );
  OAI21_X1 U37561 ( .B1(\IR/n61 ), .B2(n55293), .A(n55292), .ZN(n1176) );
  OAI21_X1 U37562 ( .B1(\intadd_6/n1 ), .B2(n54923), .A(n54922), .ZN(n54924)
         );
  XOR2_X1 U37563 ( .A(n54925), .B(n54924), .Z(n19108) );
  AND2_X1 U37564 ( .A1(n53611), .A2(n54926), .ZN(n20899) );
  NOR2_X1 U37565 ( .A1(w_IR_OUT[26]), .A2(n55128), .ZN(n3022) );
  NOR2_X1 U37566 ( .A1(n53678), .A2(n55128), .ZN(n3024) );
  INV_X1 U37567 ( .A(n55208), .ZN(n55027) );
  AOI22_X1 U37568 ( .A1(n53650), .A2(n55027), .B1(n53366), .B2(n53705), .ZN(
        n3026) );
  INV_X1 U37569 ( .A(n55205), .ZN(n54927) );
  AOI22_X1 U37570 ( .A1(n53650), .A2(n54927), .B1(n53367), .B2(n53705), .ZN(
        n3027) );
  NAND2_X1 U37571 ( .A1(n55332), .A2(n49955), .ZN(n54934) );
  AOI21_X1 U37572 ( .B1(n53368), .B2(n53799), .A(n54930), .ZN(n54928) );
  MUX2_X1 U37573 ( .A(n54928), .B(n55238), .S(n53650), .Z(n3028) );
  INV_X1 U37574 ( .A(n55235), .ZN(n54994) );
  OAI21_X1 U37575 ( .B1(n54932), .B2(n49958), .A(n53799), .ZN(n54929) );
  AOI22_X1 U37576 ( .A1(n53650), .A2(n54994), .B1(n54929), .B2(n53705), .ZN(
        n3029) );
  INV_X1 U37577 ( .A(n55241), .ZN(n54985) );
  OAI21_X1 U37578 ( .B1(n54930), .B2(n53369), .A(n54963), .ZN(n54931) );
  AOI22_X1 U37579 ( .A1(n53650), .A2(n54985), .B1(n54931), .B2(n53705), .ZN(
        n3032) );
  AOI21_X1 U37580 ( .B1(n53370), .B2(n54934), .A(n54932), .ZN(n54933) );
  MUX2_X1 U37581 ( .A(n54933), .B(n55242), .S(n53650), .Z(n3033) );
  OAI21_X1 U37582 ( .B1(n55332), .B2(n49955), .A(n54934), .ZN(n54935) );
  AOI22_X1 U37583 ( .A1(n53650), .A2(n55204), .B1(n54935), .B2(n53705), .ZN(
        n3034) );
  INV_X1 U37584 ( .A(n55207), .ZN(n54937) );
  OAI21_X1 U37585 ( .B1(n55134), .B2(n53372), .A(n55333), .ZN(n54936) );
  AOI22_X1 U37586 ( .A1(n53650), .A2(n54937), .B1(n54936), .B2(n53705), .ZN(
        n3036) );
  NAND2_X1 U37587 ( .A1(n54969), .A2(n53384), .ZN(n54965) );
  AOI21_X1 U37588 ( .B1(n54947), .B2(n49942), .A(n53650), .ZN(n54938) );
  INV_X1 U37589 ( .A(n54938), .ZN(n54939) );
  OAI22_X1 U37590 ( .A1(n54941), .A2(n54939), .B1(n53705), .B2(n55214), .ZN(
        n3038) );
  OAI21_X1 U37591 ( .B1(n54982), .B2(n53373), .A(n53685), .ZN(n54940) );
  AOI22_X1 U37592 ( .A1(n53650), .A2(n55222), .B1(n54940), .B2(n53705), .ZN(
        n3039) );
  OAI21_X1 U37593 ( .B1(n54941), .B2(n53374), .A(n54974), .ZN(n54942) );
  AOI22_X1 U37594 ( .A1(n53650), .A2(n55203), .B1(n54942), .B2(n53705), .ZN(
        n3040) );
  OAI21_X1 U37595 ( .B1(n54977), .B2(n53375), .A(n53694), .ZN(n54943) );
  AOI22_X1 U37596 ( .A1(n53650), .A2(n55210), .B1(n54943), .B2(n53705), .ZN(
        n3041) );
  AOI21_X1 U37597 ( .B1(n54955), .B2(n53376), .A(n53650), .ZN(n54944) );
  INV_X1 U37598 ( .A(n54944), .ZN(n54945) );
  OAI22_X1 U37599 ( .A1(n54953), .A2(n54945), .B1(n53705), .B2(n55202), .ZN(
        n3042) );
  INV_X1 U37600 ( .A(n55250), .ZN(n55078) );
  OAI21_X1 U37601 ( .B1(n54961), .B2(n53377), .A(n54957), .ZN(n54946) );
  AOI22_X1 U37602 ( .A1(n53650), .A2(n55078), .B1(n54946), .B2(n53705), .ZN(
        n3043) );
  OAI21_X1 U37603 ( .B1(n54951), .B2(n53378), .A(n54947), .ZN(n54948) );
  AOI22_X1 U37604 ( .A1(n53650), .A2(n55052), .B1(n54948), .B2(n53705), .ZN(
        n3044) );
  AOI21_X1 U37605 ( .B1(n54952), .B2(n53379), .A(n53650), .ZN(n54949) );
  INV_X1 U37606 ( .A(n54949), .ZN(n54950) );
  OAI22_X1 U37607 ( .A1(n54951), .A2(n54950), .B1(n53705), .B2(n55213), .ZN(
        n3045) );
  OAI21_X1 U37608 ( .B1(n54953), .B2(n53380), .A(n54952), .ZN(n54954) );
  AOI22_X1 U37609 ( .A1(n53650), .A2(n55212), .B1(n54954), .B2(n53705), .ZN(
        n3046) );
  OAI21_X1 U37610 ( .B1(n54960), .B2(n53381), .A(n54955), .ZN(n54956) );
  AOI22_X1 U37611 ( .A1(n53650), .A2(n55220), .B1(n54956), .B2(n53705), .ZN(
        n3047) );
  AOI21_X1 U37612 ( .B1(n54957), .B2(n53382), .A(n53650), .ZN(n54958) );
  INV_X1 U37613 ( .A(n54958), .ZN(n54959) );
  OAI22_X1 U37614 ( .A1(n54960), .A2(n54959), .B1(n53705), .B2(n55201), .ZN(
        n3048) );
  AOI21_X1 U37615 ( .B1(n49951), .B2(n54965), .A(n54961), .ZN(n54962) );
  MUX2_X1 U37616 ( .A(n54962), .B(n55249), .S(n53650), .Z(n3049) );
  AOI21_X1 U37617 ( .B1(n53383), .B2(n54963), .A(n54967), .ZN(n54964) );
  MUX2_X1 U37618 ( .A(n54964), .B(n55240), .S(n53650), .Z(n3050) );
  INV_X1 U37619 ( .A(n55236), .ZN(n55087) );
  OAI21_X1 U37620 ( .B1(n54969), .B2(n53384), .A(n54965), .ZN(n54966) );
  AOI22_X1 U37621 ( .A1(n53650), .A2(n55087), .B1(n54966), .B2(n53705), .ZN(
        n3051) );
  OAI21_X1 U37622 ( .B1(n54967), .B2(n49952), .A(n54970), .ZN(n54968) );
  AOI22_X1 U37623 ( .A1(n53650), .A2(n55243), .B1(n54968), .B2(n53705), .ZN(
        n3052) );
  AOI21_X1 U37624 ( .B1(n53385), .B2(n54970), .A(n54969), .ZN(n54971) );
  MUX2_X1 U37625 ( .A(n54971), .B(n55237), .S(n53650), .Z(n3053) );
  AOI21_X1 U37626 ( .B1(n53685), .B2(n53386), .A(n53650), .ZN(n54972) );
  INV_X1 U37627 ( .A(n54972), .ZN(n54973) );
  OAI22_X1 U37628 ( .A1(n54978), .A2(n54973), .B1(n53705), .B2(n55223), .ZN(
        n3054) );
  AOI21_X1 U37629 ( .B1(n54974), .B2(n53387), .A(n53650), .ZN(n54975) );
  INV_X1 U37630 ( .A(n54975), .ZN(n54976) );
  OAI22_X1 U37631 ( .A1(n54977), .A2(n54976), .B1(n53705), .B2(n55209), .ZN(
        n3055) );
  XNOR2_X1 U37632 ( .A(n53388), .B(n54978), .ZN(n54979) );
  AOI22_X1 U37633 ( .A1(n53650), .A2(n55215), .B1(n54979), .B2(n53705), .ZN(
        n3056) );
  AOI21_X1 U37634 ( .B1(n53694), .B2(n49937), .A(n53650), .ZN(n54980) );
  INV_X1 U37635 ( .A(n54980), .ZN(n54981) );
  OAI22_X1 U37636 ( .A1(n54982), .A2(n54981), .B1(n53705), .B2(n55221), .ZN(
        n3057) );
  OAI22_X1 U37637 ( .A1(n49843), .A2(n55116), .B1(n53511), .B2(n55120), .ZN(
        n54983) );
  AOI21_X1 U37638 ( .B1(n55118), .B2(n53462), .A(n54983), .ZN(n54984) );
  OAI21_X1 U37639 ( .B1(n54985), .B2(n55115), .A(n54984), .ZN(n3058) );
  OAI22_X1 U37640 ( .A1(n49843), .A2(n55103), .B1(n53430), .B2(n55126), .ZN(
        n54986) );
  AOI21_X1 U37641 ( .B1(n55241), .B2(n55122), .A(n54986), .ZN(n54987) );
  OAI21_X1 U37642 ( .B1(n53389), .B2(n55106), .A(n54987), .ZN(n3059) );
  AOI22_X1 U37643 ( .A1(n53461), .A2(n55118), .B1(n55099), .B2(n53756), .ZN(
        n54989) );
  NAND2_X1 U37644 ( .A1(n55238), .A2(n55100), .ZN(n54988) );
  OAI211_X1 U37645 ( .C1(n53512), .C2(n55120), .A(n54989), .B(n54988), .ZN(
        n3061) );
  OAI22_X1 U37646 ( .A1(n49808), .A2(n55103), .B1(n53429), .B2(n55126), .ZN(
        n54990) );
  AOI21_X1 U37647 ( .B1(n55238), .B2(n55122), .A(n54990), .ZN(n54991) );
  OAI21_X1 U37648 ( .B1(n53390), .B2(n55106), .A(n54991), .ZN(n3062) );
  OAI22_X1 U37649 ( .A1(n49832), .A2(n55116), .B1(n53514), .B2(n55120), .ZN(
        n54992) );
  AOI21_X1 U37650 ( .B1(n55118), .B2(n53460), .A(n54992), .ZN(n54993) );
  OAI21_X1 U37651 ( .B1(n54994), .B2(n55115), .A(n54993), .ZN(n3064) );
  OAI22_X1 U37652 ( .A1(n49832), .A2(n55103), .B1(n53428), .B2(n55126), .ZN(
        n54995) );
  AOI21_X1 U37653 ( .B1(n55235), .B2(n55122), .A(n54995), .ZN(n54996) );
  OAI21_X1 U37654 ( .B1(n53391), .B2(n55106), .A(n54996), .ZN(n3065) );
  AOI22_X1 U37655 ( .A1(n7676), .A2(n55099), .B1(n55118), .B2(n53459), .ZN(
        n54998) );
  NAND2_X1 U37656 ( .A1(n55242), .A2(n55100), .ZN(n54997) );
  OAI211_X1 U37657 ( .C1(n53507), .C2(n55120), .A(n54998), .B(n54997), .ZN(
        n3067) );
  OAI22_X1 U37658 ( .A1(n53427), .A2(n55126), .B1(n53661), .B2(n55103), .ZN(
        n54999) );
  AOI21_X1 U37659 ( .B1(n55242), .B2(n55122), .A(n54999), .ZN(n55000) );
  OAI21_X1 U37660 ( .B1(n53392), .B2(n55106), .A(n55000), .ZN(n3068) );
  OAI22_X1 U37661 ( .A1(n53508), .A2(n55120), .B1(n55116), .B2(n53662), .ZN(
        n55001) );
  AOI21_X1 U37662 ( .B1(n55118), .B2(n53458), .A(n55001), .ZN(n55002) );
  OAI21_X1 U37663 ( .B1(n55204), .B2(n55115), .A(n55002), .ZN(n3070) );
  OAI22_X1 U37664 ( .A1(n53393), .A2(n55106), .B1(n53426), .B2(n55126), .ZN(
        n55003) );
  AOI21_X1 U37665 ( .B1(n7620), .B2(n53645), .A(n55003), .ZN(n55004) );
  OAI21_X1 U37666 ( .B1(n55204), .B2(n55077), .A(n55004), .ZN(n3071) );
  AOI22_X1 U37667 ( .A1(n53457), .A2(n55118), .B1(n55099), .B2(n53757), .ZN(
        n55006) );
  NAND2_X1 U37668 ( .A1(n55100), .A2(n55334), .ZN(n55005) );
  OAI211_X1 U37669 ( .C1(n53509), .C2(n55120), .A(n55006), .B(n55005), .ZN(
        n3073) );
  OAI22_X1 U37670 ( .A1(n49811), .A2(n55103), .B1(n53425), .B2(n55126), .ZN(
        n55007) );
  AOI21_X1 U37671 ( .B1(n55122), .B2(n55334), .A(n55007), .ZN(n55008) );
  OAI21_X1 U37672 ( .B1(n53394), .B2(n55106), .A(n55008), .ZN(n3074) );
  AOI22_X1 U37673 ( .A1(n53456), .A2(n55118), .B1(n55099), .B2(DRAM_ADDR[5]), 
        .ZN(n55010) );
  NAND2_X1 U37674 ( .A1(n55100), .A2(n55207), .ZN(n55009) );
  OAI211_X1 U37675 ( .C1(n53510), .C2(n55120), .A(n55010), .B(n55009), .ZN(
        n3076) );
  OAI22_X1 U37676 ( .A1(n3249), .A2(n55103), .B1(n53424), .B2(n55126), .ZN(
        n55011) );
  AOI21_X1 U37677 ( .B1(n55122), .B2(n55207), .A(n55011), .ZN(n55012) );
  OAI21_X1 U37678 ( .B1(n53395), .B2(n55106), .A(n55012), .ZN(n3077) );
  INV_X1 U37679 ( .A(n55206), .ZN(n55132) );
  OAI22_X1 U37680 ( .A1(n3248), .A2(n55116), .B1(n53503), .B2(n55120), .ZN(
        n55013) );
  AOI21_X1 U37681 ( .B1(n55118), .B2(n53455), .A(n55013), .ZN(n55014) );
  OAI21_X1 U37682 ( .B1(n55132), .B2(n55115), .A(n55014), .ZN(n3079) );
  OAI22_X1 U37683 ( .A1(n3248), .A2(n55103), .B1(n53423), .B2(n55126), .ZN(
        n55015) );
  AOI21_X1 U37684 ( .B1(n55122), .B2(n55206), .A(n55015), .ZN(n55016) );
  OAI21_X1 U37685 ( .B1(n53396), .B2(n55106), .A(n55016), .ZN(n3080) );
  AOI22_X1 U37686 ( .A1(n53454), .A2(n55118), .B1(n55099), .B2(DRAM_ADDR[3]), 
        .ZN(n55018) );
  NAND2_X1 U37687 ( .A1(n55100), .A2(n55239), .ZN(n55017) );
  OAI211_X1 U37688 ( .C1(n53504), .C2(n55120), .A(n55018), .B(n55017), .ZN(
        n3082) );
  OAI22_X1 U37689 ( .A1(n3254), .A2(n55103), .B1(n53422), .B2(n55126), .ZN(
        n55019) );
  AOI21_X1 U37690 ( .B1(n55122), .B2(n55239), .A(n55019), .ZN(n55020) );
  OAI21_X1 U37691 ( .B1(n53397), .B2(n55106), .A(n55020), .ZN(n3083) );
  AOI22_X1 U37692 ( .A1(n53453), .A2(n55118), .B1(n55099), .B2(DRAM_ADDR[2]), 
        .ZN(n55022) );
  NAND2_X1 U37693 ( .A1(n55100), .A2(n55336), .ZN(n55021) );
  OAI211_X1 U37694 ( .C1(n53505), .C2(n55120), .A(n55022), .B(n55021), .ZN(
        n3085) );
  OAI22_X1 U37695 ( .A1(n3247), .A2(n55103), .B1(n53421), .B2(n55126), .ZN(
        n55023) );
  AOI21_X1 U37696 ( .B1(n55122), .B2(n55336), .A(n55023), .ZN(n55024) );
  OAI21_X1 U37697 ( .B1(n53398), .B2(n55106), .A(n55024), .ZN(n3086) );
  OAI22_X1 U37698 ( .A1(n3273), .A2(n55116), .B1(n53506), .B2(n55120), .ZN(
        n55025) );
  AOI21_X1 U37699 ( .B1(n55118), .B2(n53452), .A(n55025), .ZN(n55026) );
  OAI21_X1 U37700 ( .B1(n55027), .B2(n55115), .A(n55026), .ZN(n3088) );
  OAI22_X1 U37701 ( .A1(n3273), .A2(n55103), .B1(n53420), .B2(n55126), .ZN(
        n55028) );
  AOI21_X1 U37702 ( .B1(n55122), .B2(n55208), .A(n55028), .ZN(n55029) );
  OAI21_X1 U37703 ( .B1(n53399), .B2(n55106), .A(n55029), .ZN(n3089) );
  AOI22_X1 U37704 ( .A1(n53451), .A2(n55118), .B1(n55099), .B2(DRAM_ADDR[0]), 
        .ZN(n55031) );
  NAND2_X1 U37705 ( .A1(n55100), .A2(n55205), .ZN(n55030) );
  OAI211_X1 U37706 ( .C1(n53499), .C2(n55120), .A(n55031), .B(n55030), .ZN(
        n3091) );
  OAI22_X1 U37707 ( .A1(n3260), .A2(n55103), .B1(n53419), .B2(n55126), .ZN(
        n55032) );
  AOI21_X1 U37708 ( .B1(n55122), .B2(n55205), .A(n55032), .ZN(n55033) );
  OAI21_X1 U37709 ( .B1(n53400), .B2(n55106), .A(n55033), .ZN(n3092) );
  OAI22_X1 U37710 ( .A1(n53665), .A2(n55116), .B1(n55221), .B2(n55115), .ZN(
        n55034) );
  AOI21_X1 U37711 ( .B1(n55118), .B2(n53479), .A(n55034), .ZN(n55035) );
  OAI21_X1 U37712 ( .B1(n53500), .B2(n55120), .A(n55035), .ZN(n3094) );
  INV_X1 U37713 ( .A(n55221), .ZN(n55036) );
  AOI22_X1 U37714 ( .A1(n49872), .A2(n53645), .B1(n55036), .B2(n55122), .ZN(
        n55037) );
  OAI211_X1 U37715 ( .C1(n53447), .C2(n55126), .A(n55037), .B(n55124), .ZN(
        n3095) );
  OAI22_X1 U37716 ( .A1(n55210), .A2(n55115), .B1(n53672), .B2(n55116), .ZN(
        n55038) );
  AOI21_X1 U37717 ( .B1(n55118), .B2(n53478), .A(n55038), .ZN(n55039) );
  OAI21_X1 U37718 ( .B1(n53501), .B2(n55120), .A(n55039), .ZN(n3098) );
  INV_X1 U37719 ( .A(n55210), .ZN(n55040) );
  AOI22_X1 U37720 ( .A1(n55040), .A2(n55122), .B1(n7623), .B2(n53645), .ZN(
        n55041) );
  OAI211_X1 U37721 ( .C1(n53446), .C2(n55126), .A(n55041), .B(n55124), .ZN(
        n3099) );
  OAI22_X1 U37722 ( .A1(n49838), .A2(n55116), .B1(n55209), .B2(n55115), .ZN(
        n55042) );
  AOI21_X1 U37723 ( .B1(n55118), .B2(n53477), .A(n55042), .ZN(n55043) );
  OAI21_X1 U37724 ( .B1(n53502), .B2(n55120), .A(n55043), .ZN(n3101) );
  INV_X1 U37725 ( .A(n55209), .ZN(n55044) );
  AOI22_X1 U37726 ( .A1(n55044), .A2(n55122), .B1(n53645), .B2(n53648), .ZN(
        n55045) );
  OAI211_X1 U37727 ( .C1(n53445), .C2(n55126), .A(n55045), .B(n55124), .ZN(
        n3102) );
  OAI22_X1 U37728 ( .A1(n49839), .A2(n55116), .B1(n55214), .B2(n55115), .ZN(
        n55046) );
  AOI21_X1 U37729 ( .B1(n55118), .B2(n53475), .A(n55046), .ZN(n55047) );
  OAI21_X1 U37730 ( .B1(n53495), .B2(n55120), .A(n55047), .ZN(n3104) );
  OAI22_X1 U37731 ( .A1(n53443), .A2(n55126), .B1(n55214), .B2(n55077), .ZN(
        n55048) );
  AOI21_X1 U37732 ( .B1(n53645), .B2(n53706), .A(n55048), .ZN(n55049) );
  OAI21_X1 U37733 ( .B1(n53401), .B2(n55106), .A(n55049), .ZN(n3105) );
  OAI22_X1 U37734 ( .A1(n55052), .A2(n55115), .B1(n53669), .B2(n55116), .ZN(
        n55050) );
  AOI21_X1 U37735 ( .B1(n55118), .B2(n53474), .A(n55050), .ZN(n55051) );
  OAI21_X1 U37736 ( .B1(n53496), .B2(n55120), .A(n55051), .ZN(n3124) );
  OAI22_X1 U37737 ( .A1(n53442), .A2(n55126), .B1(n55052), .B2(n55077), .ZN(
        n55053) );
  AOI21_X1 U37738 ( .B1(n7661), .B2(n53645), .A(n55053), .ZN(n55054) );
  OAI21_X1 U37739 ( .B1(n53402), .B2(n55106), .A(n55054), .ZN(n3125) );
  OAI22_X1 U37740 ( .A1(n55213), .A2(n55115), .B1(n53670), .B2(n55116), .ZN(
        n55055) );
  AOI21_X1 U37741 ( .B1(n55118), .B2(n53473), .A(n55055), .ZN(n55056) );
  OAI21_X1 U37742 ( .B1(n53497), .B2(n55120), .A(n55056), .ZN(n3126) );
  OAI22_X1 U37743 ( .A1(n53441), .A2(n55126), .B1(n55213), .B2(n55077), .ZN(
        n55057) );
  AOI21_X1 U37744 ( .B1(n7622), .B2(n53645), .A(n55057), .ZN(n55058) );
  OAI21_X1 U37745 ( .B1(n53403), .B2(n55106), .A(n55058), .ZN(n3127) );
  OAI22_X1 U37746 ( .A1(n55212), .A2(n55115), .B1(n53668), .B2(n55116), .ZN(
        n55059) );
  AOI21_X1 U37747 ( .B1(n55118), .B2(n53472), .A(n55059), .ZN(n55060) );
  OAI21_X1 U37748 ( .B1(n53498), .B2(n55120), .A(n55060), .ZN(n3128) );
  OAI22_X1 U37749 ( .A1(n53440), .A2(n55126), .B1(n55212), .B2(n55077), .ZN(
        n55061) );
  AOI21_X1 U37750 ( .B1(n7660), .B2(n53645), .A(n55061), .ZN(n55062) );
  OAI21_X1 U37751 ( .B1(n53404), .B2(n55106), .A(n55062), .ZN(n3129) );
  OAI22_X1 U37752 ( .A1(n55202), .A2(n55115), .B1(n53667), .B2(n55116), .ZN(
        n55063) );
  AOI21_X1 U37753 ( .B1(n55118), .B2(n53471), .A(n55063), .ZN(n55064) );
  OAI21_X1 U37754 ( .B1(n53491), .B2(n55120), .A(n55064), .ZN(n3130) );
  OAI22_X1 U37755 ( .A1(n53439), .A2(n55126), .B1(n55202), .B2(n55077), .ZN(
        n55065) );
  AOI21_X1 U37756 ( .B1(n7621), .B2(n53645), .A(n55065), .ZN(n55066) );
  OAI21_X1 U37757 ( .B1(n53405), .B2(n55106), .A(n55066), .ZN(n3131) );
  OAI22_X1 U37758 ( .A1(n49815), .A2(n55116), .B1(n55220), .B2(n55115), .ZN(
        n55067) );
  AOI21_X1 U37759 ( .B1(n55118), .B2(n53470), .A(n55067), .ZN(n55068) );
  OAI21_X1 U37760 ( .B1(n53492), .B2(n55120), .A(n55068), .ZN(n3132) );
  OAI22_X1 U37761 ( .A1(n53438), .A2(n55126), .B1(n55220), .B2(n55077), .ZN(
        n55069) );
  AOI21_X1 U37762 ( .B1(n53645), .B2(n53708), .A(n55069), .ZN(n55070) );
  OAI21_X1 U37763 ( .B1(n53406), .B2(n55106), .A(n55070), .ZN(n3133) );
  OAI22_X1 U37764 ( .A1(n55201), .A2(n55115), .B1(n53666), .B2(n55116), .ZN(
        n55071) );
  AOI21_X1 U37765 ( .B1(n55118), .B2(n53469), .A(n55071), .ZN(n55072) );
  OAI21_X1 U37766 ( .B1(n53493), .B2(n55120), .A(n55072), .ZN(n3134) );
  OAI22_X1 U37767 ( .A1(n53437), .A2(n55126), .B1(n55201), .B2(n55077), .ZN(
        n55073) );
  AOI21_X1 U37768 ( .B1(n7663), .B2(n53645), .A(n55073), .ZN(n55074) );
  OAI21_X1 U37769 ( .B1(n53407), .B2(n55106), .A(n55074), .ZN(n3135) );
  OAI22_X1 U37770 ( .A1(n49844), .A2(n55116), .B1(n55078), .B2(n55115), .ZN(
        n55075) );
  AOI21_X1 U37771 ( .B1(n55118), .B2(n53468), .A(n55075), .ZN(n55076) );
  OAI21_X1 U37772 ( .B1(n53494), .B2(n55120), .A(n55076), .ZN(n3136) );
  OAI22_X1 U37773 ( .A1(n53436), .A2(n55126), .B1(n55078), .B2(n55077), .ZN(
        n55079) );
  AOI21_X1 U37774 ( .B1(n53645), .B2(n53707), .A(n55079), .ZN(n55080) );
  OAI21_X1 U37775 ( .B1(n53408), .B2(n55106), .A(n55080), .ZN(n3137) );
  AOI22_X1 U37776 ( .A1(n55249), .A2(n55100), .B1(n55118), .B2(n53467), .ZN(
        n55082) );
  NAND2_X1 U37777 ( .A1(n7662), .A2(n55099), .ZN(n55081) );
  OAI211_X1 U37778 ( .C1(n53487), .C2(n55120), .A(n55082), .B(n55081), .ZN(
        n3138) );
  OAI22_X1 U37779 ( .A1(n53435), .A2(n55126), .B1(n53671), .B2(n55103), .ZN(
        n55083) );
  AOI21_X1 U37780 ( .B1(n55249), .B2(n55122), .A(n55083), .ZN(n55084) );
  OAI21_X1 U37781 ( .B1(n53409), .B2(n55106), .A(n55084), .ZN(n3139) );
  OAI22_X1 U37782 ( .A1(n49809), .A2(n55116), .B1(n53488), .B2(n55120), .ZN(
        n55085) );
  AOI21_X1 U37783 ( .B1(n55118), .B2(n53466), .A(n55085), .ZN(n55086) );
  OAI21_X1 U37784 ( .B1(n55087), .B2(n55115), .A(n55086), .ZN(n3140) );
  OAI22_X1 U37785 ( .A1(n49809), .A2(n55103), .B1(n53434), .B2(n55126), .ZN(
        n55088) );
  AOI21_X1 U37786 ( .B1(n55236), .B2(n55122), .A(n55088), .ZN(n55089) );
  OAI21_X1 U37787 ( .B1(n53410), .B2(n55106), .A(n55089), .ZN(n3141) );
  AOI22_X1 U37788 ( .A1(n7624), .A2(n55099), .B1(n55118), .B2(n53465), .ZN(
        n55091) );
  NAND2_X1 U37789 ( .A1(n55237), .A2(n55100), .ZN(n55090) );
  OAI211_X1 U37790 ( .C1(n53489), .C2(n55120), .A(n55091), .B(n55090), .ZN(
        n3142) );
  OAI22_X1 U37791 ( .A1(n53433), .A2(n55126), .B1(n53660), .B2(n55103), .ZN(
        n55092) );
  AOI21_X1 U37792 ( .B1(n55237), .B2(n55122), .A(n55092), .ZN(n55093) );
  OAI21_X1 U37793 ( .B1(n53411), .B2(n55106), .A(n55093), .ZN(n3143) );
  OAI22_X1 U37794 ( .A1(n49810), .A2(n55116), .B1(n53490), .B2(n55120), .ZN(
        n55094) );
  AOI21_X1 U37795 ( .B1(n55118), .B2(n53464), .A(n55094), .ZN(n55095) );
  OAI21_X1 U37796 ( .B1(n55243), .B2(n55115), .A(n55095), .ZN(n3144) );
  OAI22_X1 U37797 ( .A1(n49810), .A2(n55103), .B1(n53432), .B2(n55126), .ZN(
        n55096) );
  AOI21_X1 U37798 ( .B1(n55097), .B2(n55122), .A(n55096), .ZN(n55098) );
  OAI21_X1 U37799 ( .B1(n53412), .B2(n55106), .A(n55098), .ZN(n3145) );
  AOI22_X1 U37800 ( .A1(n53463), .A2(n55118), .B1(n55099), .B2(n53755), .ZN(
        n55102) );
  NAND2_X1 U37801 ( .A1(n55240), .A2(n55100), .ZN(n55101) );
  OAI211_X1 U37802 ( .C1(n53483), .C2(n55120), .A(n55102), .B(n55101), .ZN(
        n3146) );
  OAI22_X1 U37803 ( .A1(n49814), .A2(n55103), .B1(n53431), .B2(n55126), .ZN(
        n55104) );
  AOI21_X1 U37804 ( .B1(n55240), .B2(n55122), .A(n55104), .ZN(n55105) );
  OAI21_X1 U37805 ( .B1(n53413), .B2(n55106), .A(n55105), .ZN(n3147) );
  OAI22_X1 U37806 ( .A1(n49834), .A2(n55116), .B1(n55115), .B2(n55223), .ZN(
        n55107) );
  AOI21_X1 U37807 ( .B1(n55118), .B2(n53481), .A(n55107), .ZN(n55108) );
  OAI21_X1 U37808 ( .B1(n53486), .B2(n55120), .A(n55108), .ZN(n3148) );
  INV_X1 U37809 ( .A(n55223), .ZN(n55109) );
  AOI22_X1 U37810 ( .A1(n55122), .A2(n55109), .B1(n53645), .B2(n53710), .ZN(
        n55110) );
  OAI211_X1 U37811 ( .C1(n53449), .C2(n55126), .A(n55110), .B(n55124), .ZN(
        n3149) );
  OAI22_X1 U37812 ( .A1(n53663), .A2(n55116), .B1(n55222), .B2(n55115), .ZN(
        n55111) );
  AOI21_X1 U37813 ( .B1(n55118), .B2(n53480), .A(n55111), .ZN(n55112) );
  OAI21_X1 U37814 ( .B1(n53484), .B2(n55120), .A(n55112), .ZN(n3150) );
  INV_X1 U37815 ( .A(n55222), .ZN(n55113) );
  AOI22_X1 U37816 ( .A1(n7625), .A2(n53645), .B1(n55113), .B2(n55122), .ZN(
        n55114) );
  OAI211_X1 U37817 ( .C1(n53448), .C2(n55126), .A(n55114), .B(n55124), .ZN(
        n3151) );
  OAI22_X1 U37818 ( .A1(n49842), .A2(n55116), .B1(n55203), .B2(n55115), .ZN(
        n55117) );
  AOI21_X1 U37819 ( .B1(n55118), .B2(n53476), .A(n55117), .ZN(n55119) );
  OAI21_X1 U37820 ( .B1(n53485), .B2(n55120), .A(n55119), .ZN(n3152) );
  INV_X1 U37821 ( .A(n55203), .ZN(n55123) );
  AOI22_X1 U37822 ( .A1(n55123), .A2(n55122), .B1(n53645), .B2(n53709), .ZN(
        n55125) );
  OAI211_X1 U37823 ( .C1(n53444), .C2(n55126), .A(n55125), .B(n55124), .ZN(
        n3153) );
  NOR2_X1 U37824 ( .A1(w_IR_OUT[30]), .A2(n55127), .ZN(n3190) );
  NOR2_X1 U37825 ( .A1(w_IR_OUT[28]), .A2(n55128), .ZN(n3191) );
  INV_X1 U37826 ( .A(n55286), .ZN(n55296) );
  NAND2_X1 U37827 ( .A1(n55342), .A2(w_PC_OUT[9]), .ZN(n55341) );
  NAND2_X1 U37828 ( .A1(n55317), .A2(w_PC_OUT[13]), .ZN(n55348) );
  NAND2_X1 U37829 ( .A1(n55349), .A2(w_PC_OUT[17]), .ZN(n55352) );
  NAND2_X1 U37830 ( .A1(n55351), .A2(w_PC_OUT[19]), .ZN(n55321) );
  NAND2_X1 U37831 ( .A1(n55355), .A2(w_PC_OUT[21]), .ZN(n55353) );
  AOI211_X1 U37832 ( .C1(n55353), .C2(n53655), .A(n55323), .B(n53815), .ZN(
        n40059) );
  AOI211_X1 U37833 ( .C1(n55321), .C2(n53658), .A(n55355), .B(n53815), .ZN(
        n40060) );
  AOI211_X1 U37834 ( .C1(n55344), .C2(n53659), .A(n55317), .B(n53815), .ZN(
        n40065) );
  AOI211_X1 U37835 ( .C1(n55341), .C2(n53656), .A(n55345), .B(n53815), .ZN(
        n43886) );
  INV_X1 U37836 ( .A(n55239), .ZN(n55130) );
  XNOR2_X1 U37837 ( .A(n49938), .B(n49939), .ZN(n55129) );
  AOI22_X1 U37838 ( .A1(n53650), .A2(n55130), .B1(n55129), .B2(n53705), .ZN(
        n43968) );
  NOR2_X1 U37839 ( .A1(n49938), .A2(n49939), .ZN(n55131) );
  OAI21_X1 U37840 ( .B1(n55131), .B2(n53743), .A(n53705), .ZN(n55133) );
  OAI22_X1 U37841 ( .A1(n55134), .A2(n55133), .B1(n55132), .B2(n53705), .ZN(
        n43969) );
  AOI211_X1 U37842 ( .C1(n55338), .C2(n53657), .A(n55342), .B(n53815), .ZN(
        n47726) );
  AOI211_X1 U37843 ( .C1(n49907), .C2(n53793), .A(n55339), .B(n53815), .ZN(
        n47727) );
  AOI22_X1 U37844 ( .A1(n55137), .A2(n55136), .B1(n53807), .B2(n55135), .ZN(
        n55143) );
  AOI22_X1 U37845 ( .A1(n55175), .A2(\DP/ALU0/s_A_SHIFT[1] ), .B1(
        \DP/ALU0/s_A_SHIFT[9] ), .B2(n55174), .ZN(n55138) );
  OAI211_X1 U37846 ( .C1(n55141), .C2(n55140), .A(n55139), .B(n55138), .ZN(
        n55142) );
  OAI211_X1 U37847 ( .C1(n55144), .C2(n53761), .A(n55143), .B(n55142), .ZN(
        n55197) );
  NAND4_X1 U37848 ( .A1(\intadd_0/SUM[25] ), .A2(\intadd_0/SUM[24] ), .A3(
        \intadd_0/SUM[23] ), .A4(\intadd_0/SUM[22] ), .ZN(n55148) );
  NAND4_X1 U37849 ( .A1(\intadd_0/SUM[21] ), .A2(\intadd_0/SUM[20] ), .A3(
        \intadd_0/SUM[19] ), .A4(\intadd_0/SUM[18] ), .ZN(n55147) );
  NAND4_X1 U37850 ( .A1(\intadd_8/SUM[2] ), .A2(\intadd_8/SUM[1] ), .A3(
        \intadd_8/SUM[0] ), .A4(\intadd_0/SUM[26] ), .ZN(n55146) );
  XNOR2_X1 U37851 ( .A(\DP/ALU0/S_B_ADDER[0] ), .B(\DP/ALU0/s_A_ADDER[0] ), 
        .ZN(n55169) );
  NAND4_X1 U37852 ( .A1(\intadd_8/SUM[3] ), .A2(n55169), .A3(\intadd_0/SUM[3] ), .A4(\intadd_0/SUM[0] ), .ZN(n55145) );
  NOR4_X1 U37853 ( .A1(n55148), .A2(n55147), .A3(n55146), .A4(n55145), .ZN(
        n55154) );
  NAND4_X1 U37854 ( .A1(\intadd_0/SUM[7] ), .A2(\intadd_0/SUM[6] ), .A3(
        \intadd_0/SUM[9] ), .A4(\intadd_0/SUM[8] ), .ZN(n55152) );
  NAND4_X1 U37855 ( .A1(\intadd_0/SUM[2] ), .A2(\intadd_0/SUM[1] ), .A3(
        \intadd_0/SUM[5] ), .A4(\intadd_0/SUM[4] ), .ZN(n55151) );
  NAND4_X1 U37856 ( .A1(\intadd_0/SUM[17] ), .A2(\intadd_0/SUM[15] ), .A3(
        \intadd_0/SUM[14] ), .A4(\intadd_0/SUM[16] ), .ZN(n55150) );
  NAND4_X1 U37857 ( .A1(\intadd_0/SUM[11] ), .A2(\intadd_0/SUM[10] ), .A3(
        \intadd_0/SUM[13] ), .A4(\intadd_0/SUM[12] ), .ZN(n55149) );
  NOR4_X1 U37858 ( .A1(n55152), .A2(n55151), .A3(n55150), .A4(n55149), .ZN(
        n55153) );
  NAND2_X1 U37859 ( .A1(n55154), .A2(n55153), .ZN(n55156) );
  XOR2_X1 U37860 ( .A(\DP/ALU0/s_SIGN ), .B(\intadd_8/n1 ), .Z(n55159) );
  NAND2_X1 U37861 ( .A1(n55159), .A2(n53646), .ZN(n55157) );
  OAI211_X1 U37862 ( .C1(w_ALU_OPCODE[2]), .C2(n55159), .A(n55157), .B(n55156), 
        .ZN(n55155) );
  OAI21_X1 U37863 ( .B1(w_ALU_OPCODE[2]), .B2(n55156), .A(n55155), .ZN(n55162)
         );
  OAI211_X1 U37864 ( .C1(n55159), .C2(n53646), .A(n55158), .B(n55157), .ZN(
        n55160) );
  OAI22_X1 U37865 ( .A1(n55163), .A2(n55162), .B1(n55161), .B2(n55160), .ZN(
        n55171) );
  NAND2_X1 U37866 ( .A1(\DP/ALU0/s_A_LOGIC[0] ), .A2(\DP/ALU0/S_B_LOGIC[0] ), 
        .ZN(n55165) );
  NAND2_X1 U37867 ( .A1(n55187), .A2(n55165), .ZN(n55164) );
  OAI221_X1 U37868 ( .B1(n55165), .B2(n55308), .C1(\DP/ALU0/s_A_LOGIC[0] ), 
        .C2(\DP/ALU0/S_B_LOGIC[0] ), .A(n55164), .ZN(n55168) );
  NAND3_X1 U37869 ( .A1(n55166), .A2(\DP/ALU0/s_A_MULT[0] ), .A3(
        \DP/ALU0/S_B_MULT[0] ), .ZN(n55167) );
  OAI211_X1 U37870 ( .C1(n55169), .C2(n55303), .A(n55168), .B(n55167), .ZN(
        n55170) );
  AOI21_X1 U37871 ( .B1(n53810), .B2(n55171), .A(n55170), .ZN(n55185) );
  OAI22_X1 U37872 ( .A1(n55173), .A2(n53760), .B1(n55172), .B2(n53761), .ZN(
        n55183) );
  AOI222_X1 U37873 ( .A1(\DP/ALU0/s_A_SHIFT[16] ), .A2(n55176), .B1(n55175), 
        .B2(\DP/ALU0/s_A_SHIFT[0] ), .C1(\DP/ALU0/s_A_SHIFT[8] ), .C2(n53808), 
        .ZN(n55180) );
  OAI22_X1 U37874 ( .A1(n55180), .A2(n55179), .B1(n55178), .B2(n55177), .ZN(
        n55182) );
  OAI21_X1 U37875 ( .B1(n55183), .B2(n55182), .A(n55181), .ZN(n55184) );
  OAI211_X1 U37876 ( .C1(n55197), .C2(n55186), .A(n55185), .B(n55184), .ZN(
        n4925) );
  INV_X1 U37877 ( .A(\DP/ALU0/s_A_LOGIC[1] ), .ZN(n55194) );
  NOR3_X1 U37878 ( .A1(\DP/ALU0/S_B_LOGIC[1] ), .A2(n55194), .A3(n55187), .ZN(
        n55192) );
  NAND2_X1 U37879 ( .A1(\DP/ALU0/s_A_MULT[1] ), .A2(\DP/ALU0/S_B_MULT[0] ), 
        .ZN(n55189) );
  NAND2_X1 U37880 ( .A1(\DP/ALU0/s_A_MULT[0] ), .A2(\DP/ALU0/S_B_MULT[1] ), 
        .ZN(n55188) );
  XNOR2_X1 U37881 ( .A(n55189), .B(n55188), .ZN(n55190) );
  OAI22_X1 U37882 ( .A1(\intadd_0/SUM[0] ), .A2(n55303), .B1(n55300), .B2(
        n55190), .ZN(n55191) );
  AOI211_X1 U37883 ( .C1(n55193), .C2(n55306), .A(n55192), .B(n55191), .ZN(
        n55196) );
  OAI221_X1 U37884 ( .B1(\DP/ALU0/s_A_LOGIC[1] ), .B2(n53809), .C1(n55194), 
        .C2(n55308), .A(\DP/ALU0/S_B_LOGIC[1] ), .ZN(n55195) );
  OAI211_X1 U37885 ( .C1(n55197), .C2(n55312), .A(n55196), .B(n55195), .ZN(
        n4926) );
  NOR2_X1 U37886 ( .A1(n53419), .A2(n53819), .ZN(n4927) );
  NOR2_X1 U37887 ( .A1(n53420), .A2(n53821), .ZN(n4928) );
  NOR2_X1 U37888 ( .A1(n53421), .A2(n53822), .ZN(n4929) );
  NOR2_X1 U37889 ( .A1(n53422), .A2(n53822), .ZN(n4930) );
  NOR2_X1 U37890 ( .A1(n53423), .A2(n53819), .ZN(n4931) );
  NOR2_X1 U37891 ( .A1(n53424), .A2(n53819), .ZN(n4932) );
  NOR2_X1 U37892 ( .A1(n53425), .A2(n53819), .ZN(n4933) );
  NOR2_X1 U37893 ( .A1(n53426), .A2(n53819), .ZN(n4934) );
  NOR2_X1 U37894 ( .A1(n53427), .A2(n53820), .ZN(n4935) );
  NOR2_X1 U37895 ( .A1(n53428), .A2(n53822), .ZN(n4936) );
  NOR2_X1 U37896 ( .A1(n53429), .A2(n53821), .ZN(n4937) );
  NOR2_X1 U37897 ( .A1(n53430), .A2(n53822), .ZN(n4938) );
  NOR2_X1 U37898 ( .A1(n53431), .A2(n53820), .ZN(n4939) );
  NOR2_X1 U37899 ( .A1(n53432), .A2(n53820), .ZN(n4940) );
  NOR2_X1 U37900 ( .A1(n53433), .A2(n53819), .ZN(n4941) );
  NOR2_X1 U37901 ( .A1(n53434), .A2(n53821), .ZN(n4942) );
  NOR2_X1 U37902 ( .A1(n53435), .A2(n53821), .ZN(n4943) );
  NOR2_X1 U37903 ( .A1(n53436), .A2(n53820), .ZN(n4944) );
  NOR2_X1 U37904 ( .A1(n53437), .A2(n53820), .ZN(n4945) );
  NOR2_X1 U37905 ( .A1(n53438), .A2(n53819), .ZN(n4946) );
  NOR2_X1 U37906 ( .A1(n53439), .A2(n53822), .ZN(n4947) );
  NOR2_X1 U37907 ( .A1(n53440), .A2(n53820), .ZN(n4948) );
  NOR2_X1 U37908 ( .A1(n53441), .A2(n53819), .ZN(n4949) );
  NOR2_X1 U37909 ( .A1(n53442), .A2(n53821), .ZN(n4950) );
  NOR2_X1 U37910 ( .A1(n53443), .A2(n53822), .ZN(n4951) );
  NOR2_X1 U37911 ( .A1(n53444), .A2(n53821), .ZN(n4952) );
  NOR2_X1 U37912 ( .A1(n53445), .A2(n53821), .ZN(n4953) );
  NOR2_X1 U37913 ( .A1(n53446), .A2(n53821), .ZN(n4954) );
  NOR2_X1 U37914 ( .A1(n53447), .A2(n53822), .ZN(n4955) );
  NOR2_X1 U37915 ( .A1(n53448), .A2(n53819), .ZN(n4956) );
  NOR2_X1 U37916 ( .A1(n53449), .A2(n53822), .ZN(n4957) );
  NOR2_X1 U37917 ( .A1(n53450), .A2(n53822), .ZN(n4958) );
  AND2_X1 U37918 ( .A1(n53810), .A2(n53451), .ZN(n4959) );
  AND2_X1 U37919 ( .A1(n53810), .A2(n53452), .ZN(n4960) );
  AND2_X1 U37920 ( .A1(n53810), .A2(n53453), .ZN(n4961) );
  AND2_X1 U37921 ( .A1(n55198), .A2(n53454), .ZN(n4962) );
  AND2_X1 U37922 ( .A1(n55198), .A2(n53455), .ZN(n4963) );
  AND2_X1 U37923 ( .A1(n55198), .A2(n53456), .ZN(n4964) );
  AND2_X1 U37924 ( .A1(n55198), .A2(n53457), .ZN(n4965) );
  AND2_X1 U37925 ( .A1(n55198), .A2(n53458), .ZN(n4966) );
  AND2_X1 U37926 ( .A1(n55198), .A2(n53459), .ZN(n4967) );
  AND2_X1 U37927 ( .A1(n55198), .A2(n53460), .ZN(n4968) );
  AND2_X1 U37928 ( .A1(n55198), .A2(n53461), .ZN(n4969) );
  AND2_X1 U37929 ( .A1(n55198), .A2(n53462), .ZN(n4970) );
  AND2_X1 U37930 ( .A1(n55198), .A2(n53463), .ZN(n4971) );
  AND2_X1 U37931 ( .A1(n55198), .A2(n53464), .ZN(n4972) );
  AND2_X1 U37932 ( .A1(n55198), .A2(n53465), .ZN(n4973) );
  AND2_X1 U37933 ( .A1(n55198), .A2(n53466), .ZN(n4974) );
  AND2_X1 U37934 ( .A1(n53810), .A2(n53467), .ZN(n4975) );
  AND2_X1 U37935 ( .A1(n53810), .A2(n53468), .ZN(n4976) );
  AND2_X1 U37936 ( .A1(n53810), .A2(n53469), .ZN(n4977) );
  AND2_X1 U37937 ( .A1(n53810), .A2(n53470), .ZN(n4978) );
  AND2_X1 U37938 ( .A1(n53810), .A2(n53471), .ZN(n4979) );
  AND2_X1 U37939 ( .A1(n53810), .A2(n53472), .ZN(n4980) );
  AND2_X1 U37940 ( .A1(n53810), .A2(n53473), .ZN(n4981) );
  AND2_X1 U37941 ( .A1(n53810), .A2(n53474), .ZN(n4982) );
  AND2_X1 U37942 ( .A1(n53810), .A2(n53475), .ZN(n4983) );
  AND2_X1 U37943 ( .A1(n53810), .A2(n53476), .ZN(n4984) );
  AND2_X1 U37944 ( .A1(n53810), .A2(n53477), .ZN(n4985) );
  AND2_X1 U37945 ( .A1(n53810), .A2(n53478), .ZN(n4986) );
  AND2_X1 U37946 ( .A1(n53810), .A2(n53479), .ZN(n4987) );
  AND2_X1 U37947 ( .A1(n53810), .A2(n53480), .ZN(n4988) );
  AND2_X1 U37948 ( .A1(n53810), .A2(n53481), .ZN(n4989) );
  AND2_X1 U37949 ( .A1(n55198), .A2(n53482), .ZN(n4990) );
  AND2_X1 U37950 ( .A1(n55199), .A2(DRAM_DATA_IN[0]), .ZN(n4992) );
  AND2_X1 U37951 ( .A1(n55199), .A2(DRAM_DATA_IN[1]), .ZN(n4993) );
  AND2_X1 U37952 ( .A1(n55199), .A2(DRAM_DATA_IN[2]), .ZN(n4994) );
  AND2_X1 U37953 ( .A1(n55199), .A2(DRAM_DATA_IN[3]), .ZN(n4995) );
  AND2_X1 U37954 ( .A1(n55199), .A2(DRAM_DATA_IN[4]), .ZN(n4996) );
  AND2_X1 U37955 ( .A1(n55199), .A2(DRAM_DATA_IN[5]), .ZN(n4997) );
  AND2_X1 U37956 ( .A1(n55199), .A2(DRAM_DATA_IN[6]), .ZN(n4998) );
  AND2_X1 U37957 ( .A1(n55199), .A2(DRAM_DATA_IN[7]), .ZN(n4999) );
  AND2_X1 U37958 ( .A1(n55199), .A2(DRAM_DATA_IN[8]), .ZN(n5000) );
  AND2_X1 U37959 ( .A1(n55199), .A2(DRAM_DATA_IN[9]), .ZN(n5001) );
  AND2_X1 U37960 ( .A1(n55199), .A2(DRAM_DATA_IN[10]), .ZN(n5002) );
  AND2_X1 U37961 ( .A1(n55199), .A2(DRAM_DATA_IN[11]), .ZN(n5003) );
  AND2_X1 U37962 ( .A1(n55199), .A2(DRAM_DATA_IN[12]), .ZN(n5004) );
  AND2_X1 U37963 ( .A1(n55199), .A2(DRAM_DATA_IN[13]), .ZN(n5005) );
  AND2_X1 U37964 ( .A1(n55199), .A2(DRAM_DATA_IN[14]), .ZN(n5006) );
  AND2_X1 U37965 ( .A1(n55199), .A2(DRAM_DATA_IN[15]), .ZN(n5007) );
  NOR2_X1 U37966 ( .A1(n53725), .A2(n55200), .ZN(n5024) );
  NOR2_X1 U37967 ( .A1(n53718), .A2(n55200), .ZN(n5025) );
  NOR2_X1 U37968 ( .A1(n53719), .A2(n55200), .ZN(n5026) );
  NOR2_X1 U37969 ( .A1(n53728), .A2(n55200), .ZN(n5027) );
  NOR2_X1 U37970 ( .A1(n53711), .A2(n55200), .ZN(n5028) );
  NOR2_X1 U37971 ( .A1(n53715), .A2(n55200), .ZN(n5029) );
  NOR2_X1 U37972 ( .A1(n53729), .A2(n55200), .ZN(n5030) );
  NOR2_X1 U37973 ( .A1(n53742), .A2(n55200), .ZN(n5031) );
  NOR2_X1 U37974 ( .A1(n53740), .A2(n55200), .ZN(n5032) );
  NOR2_X1 U37975 ( .A1(n53714), .A2(n55200), .ZN(n5033) );
  NOR2_X1 U37976 ( .A1(n53712), .A2(n55200), .ZN(n5034) );
  NOR2_X1 U37977 ( .A1(n53726), .A2(n55200), .ZN(n5035) );
  NOR2_X1 U37978 ( .A1(n53721), .A2(n55200), .ZN(n5036) );
  NOR2_X1 U37979 ( .A1(n53723), .A2(n55200), .ZN(n5037) );
  NOR2_X1 U37980 ( .A1(n53732), .A2(n55200), .ZN(n5038) );
  NOR2_X1 U37981 ( .A1(n53722), .A2(n55200), .ZN(n5039) );
  NOR2_X1 U37982 ( .A1(n53730), .A2(n55200), .ZN(n5040) );
  NOR2_X1 U37983 ( .A1(n53720), .A2(n55200), .ZN(n5041) );
  NOR2_X1 U37984 ( .A1(n53739), .A2(n55200), .ZN(n5042) );
  NOR2_X1 U37985 ( .A1(n53716), .A2(n55200), .ZN(n5043) );
  NOR2_X1 U37986 ( .A1(n53738), .A2(n55200), .ZN(n5044) );
  NOR2_X1 U37987 ( .A1(n53731), .A2(n55200), .ZN(n5045) );
  NOR2_X1 U37988 ( .A1(n53733), .A2(n55200), .ZN(n5046) );
  NOR2_X1 U37989 ( .A1(n53735), .A2(n55200), .ZN(n5047) );
  NOR2_X1 U37990 ( .A1(n53724), .A2(n55200), .ZN(n5048) );
  NOR2_X1 U37991 ( .A1(n53727), .A2(n55200), .ZN(n5049) );
  NOR2_X1 U37992 ( .A1(n53713), .A2(n55200), .ZN(n5050) );
  NOR2_X1 U37993 ( .A1(n53737), .A2(n55200), .ZN(n5051) );
  NOR2_X1 U37994 ( .A1(n53734), .A2(n55200), .ZN(n5052) );
  NOR2_X1 U37995 ( .A1(n53736), .A2(n55200), .ZN(n5053) );
  NOR2_X1 U37996 ( .A1(n53717), .A2(n55200), .ZN(n5054) );
  NOR2_X1 U37997 ( .A1(n53741), .A2(n55200), .ZN(n5055) );
  NOR2_X1 U37998 ( .A1(n3260), .A2(n55200), .ZN(n5056) );
  NOR2_X1 U37999 ( .A1(n3273), .A2(n55200), .ZN(n5057) );
  NOR2_X1 U38000 ( .A1(n3247), .A2(n55200), .ZN(n5058) );
  NOR2_X1 U38001 ( .A1(n3254), .A2(n55200), .ZN(n5059) );
  NOR2_X1 U38002 ( .A1(n3248), .A2(n55200), .ZN(n5060) );
  NOR2_X1 U38003 ( .A1(n3249), .A2(n55200), .ZN(n5061) );
  NOR2_X1 U38004 ( .A1(n49811), .A2(n53822), .ZN(n5062) );
  NOR2_X1 U38005 ( .A1(n53821), .A2(n53662), .ZN(n5063) );
  NOR2_X1 U38006 ( .A1(n53821), .A2(n53661), .ZN(n5064) );
  NOR2_X1 U38007 ( .A1(n49832), .A2(n53819), .ZN(n5065) );
  NOR2_X1 U38008 ( .A1(n49808), .A2(n53820), .ZN(n5066) );
  NOR2_X1 U38009 ( .A1(n49843), .A2(n53820), .ZN(n5067) );
  NOR2_X1 U38010 ( .A1(n49814), .A2(n53820), .ZN(n5068) );
  NOR2_X1 U38011 ( .A1(n49810), .A2(n53820), .ZN(n5069) );
  NOR2_X1 U38012 ( .A1(n53820), .A2(n53660), .ZN(n5070) );
  NOR2_X1 U38013 ( .A1(n49809), .A2(n53819), .ZN(n5071) );
  NOR2_X1 U38014 ( .A1(n53820), .A2(n53671), .ZN(n5072) );
  NOR2_X1 U38015 ( .A1(n49844), .A2(n53819), .ZN(n5073) );
  NOR2_X1 U38016 ( .A1(n53820), .A2(n53666), .ZN(n5074) );
  NOR2_X1 U38017 ( .A1(n49815), .A2(n53819), .ZN(n5075) );
  NOR2_X1 U38018 ( .A1(n53819), .A2(n53667), .ZN(n5076) );
  NOR2_X1 U38019 ( .A1(n53819), .A2(n53668), .ZN(n5077) );
  NOR2_X1 U38020 ( .A1(n53819), .A2(n53670), .ZN(n5078) );
  NOR2_X1 U38021 ( .A1(n53821), .A2(n53669), .ZN(n5079) );
  NOR2_X1 U38022 ( .A1(n49839), .A2(n53822), .ZN(n5080) );
  NOR2_X1 U38023 ( .A1(n49842), .A2(n53821), .ZN(n5081) );
  NOR2_X1 U38024 ( .A1(n49838), .A2(n53822), .ZN(n5082) );
  NOR2_X1 U38025 ( .A1(n53821), .A2(n53672), .ZN(n5083) );
  NOR2_X1 U38026 ( .A1(n53820), .A2(n53665), .ZN(n5084) );
  NOR2_X1 U38027 ( .A1(n53820), .A2(n53663), .ZN(n5085) );
  NOR2_X1 U38028 ( .A1(n49834), .A2(n53820), .ZN(n5086) );
  NOR2_X1 U38029 ( .A1(n53822), .A2(n53664), .ZN(n5087) );
  NAND4_X1 U38030 ( .A1(n55204), .A2(n55203), .A3(n55202), .A4(n55201), .ZN(
        n55218) );
  NOR4_X1 U38031 ( .A1(n55208), .A2(n55207), .A3(n55206), .A4(n55205), .ZN(
        n55211) );
  NAND3_X1 U38032 ( .A1(n55211), .A2(n55210), .A3(n55209), .ZN(n55217) );
  NAND4_X1 U38033 ( .A1(n55215), .A2(n55214), .A3(n55213), .A4(n55212), .ZN(
        n55216) );
  NOR4_X1 U38034 ( .A1(n55219), .A2(n55218), .A3(n55217), .A4(n55216), .ZN(
        n55279) );
  NAND4_X1 U38035 ( .A1(n55223), .A2(n55222), .A3(n55221), .A4(n55220), .ZN(
        n55248) );
  OAI221_X1 U38036 ( .B1(\IR/n61 ), .B2(n53515), .C1(\DP/IMMS26[25] ), .C2(
        n53693), .A(w_RF_WE3), .ZN(n55228) );
  AOI22_X1 U38037 ( .A1(\IR/n60 ), .A2(n49866), .B1(\IR/n58 ), .B2(n49819), 
        .ZN(n55224) );
  OAI221_X1 U38038 ( .B1(\IR/n60 ), .B2(n49866), .C1(\IR/n58 ), .C2(n49819), 
        .A(n55224), .ZN(n55227) );
  AOI22_X1 U38039 ( .A1(\IR/n57 ), .A2(n49857), .B1(\DP/IMMS26[23] ), .B2(
        n7617), .ZN(n55225) );
  OAI221_X1 U38040 ( .B1(\IR/n57 ), .B2(n49857), .C1(\DP/IMMS26[23] ), .C2(
        n7617), .A(n55225), .ZN(n55226) );
  NOR3_X1 U38041 ( .A1(n55228), .A2(n55227), .A3(n55226), .ZN(n55251) );
  AOI221_X1 U38042 ( .B1(\IR/n59 ), .B2(\DP/RD4[2] ), .C1(\DP/IMMS26[23] ), 
        .C2(n3015), .A(n53654), .ZN(n55234) );
  OAI22_X1 U38043 ( .A1(\IR/n57 ), .A2(\DP/RD4[0] ), .B1(\DP/RD4[3] ), .B2(
        \IR/n60 ), .ZN(n55229) );
  AOI221_X1 U38044 ( .B1(\DP/RD4[0] ), .B2(\IR/n57 ), .C1(\DP/RD4[3] ), .C2(
        \IR/n60 ), .A(n55229), .ZN(n55233) );
  OAI22_X1 U38045 ( .A1(\IR/n58 ), .A2(\DP/RD4[1] ), .B1(\DP/RD4[4] ), .B2(
        \IR/n61 ), .ZN(n55230) );
  AOI221_X1 U38046 ( .B1(\DP/RD4[1] ), .B2(\IR/n58 ), .C1(\DP/RD4[4] ), .C2(
        \IR/n61 ), .A(n55230), .ZN(n55232) );
  AND4_X1 U38047 ( .A1(\IR/n57 ), .A2(\IR/n61 ), .A3(\IR/n60 ), .A4(\IR/n59 ), 
        .ZN(n55231) );
  NAND2_X1 U38048 ( .A1(\IR/n58 ), .A2(n55231), .ZN(n55252) );
  NAND4_X1 U38049 ( .A1(n55234), .A2(n55233), .A3(n55232), .A4(n55252), .ZN(
        n55261) );
  NOR4_X1 U38050 ( .A1(n55251), .A2(n55261), .A3(n55336), .A4(n55334), .ZN(
        n55246) );
  NOR4_X1 U38051 ( .A1(n55238), .A2(n55237), .A3(n55236), .A4(n55235), .ZN(
        n55245) );
  NOR4_X1 U38052 ( .A1(n55242), .A2(n55241), .A3(n55240), .A4(n55239), .ZN(
        n55244) );
  NAND4_X1 U38053 ( .A1(n55246), .A2(n55245), .A3(n55244), .A4(n55243), .ZN(
        n55247) );
  NOR4_X1 U38054 ( .A1(n55250), .A2(n55249), .A3(n55248), .A4(n55247), .ZN(
        n55278) );
  NAND4_X1 U38055 ( .A1(n53483), .A2(n53486), .A3(n53485), .A4(n53484), .ZN(
        n55256) );
  NAND4_X1 U38056 ( .A1(n53489), .A2(n53490), .A3(n53487), .A4(n53488), .ZN(
        n55255) );
  NAND4_X1 U38057 ( .A1(n53493), .A2(n53494), .A3(n53491), .A4(n53492), .ZN(
        n55254) );
  NAND4_X1 U38058 ( .A1(n53497), .A2(n53498), .A3(n53495), .A4(n53496), .ZN(
        n55253) );
  NOR4_X1 U38059 ( .A1(n55256), .A2(n55255), .A3(n55254), .A4(n55253), .ZN(
        n55263) );
  NAND4_X1 U38060 ( .A1(n53501), .A2(n53502), .A3(n53499), .A4(n53500), .ZN(
        n55260) );
  NAND4_X1 U38061 ( .A1(n53505), .A2(n53506), .A3(n53503), .A4(n53504), .ZN(
        n55259) );
  NAND4_X1 U38062 ( .A1(n53509), .A2(n53510), .A3(n53507), .A4(n53508), .ZN(
        n55258) );
  NAND4_X1 U38063 ( .A1(n53512), .A2(n53514), .A3(n53513), .A4(n53511), .ZN(
        n55257) );
  NOR4_X1 U38064 ( .A1(n55260), .A2(n55259), .A3(n55258), .A4(n55257), .ZN(
        n55262) );
  NAND3_X1 U38065 ( .A1(n55263), .A2(n55262), .A3(n55261), .ZN(n55275) );
  NOR4_X1 U38066 ( .A1(n7620), .A2(n7624), .A3(n7676), .A4(n7662), .ZN(n55267)
         );
  NOR4_X1 U38067 ( .A1(n7663), .A2(n7621), .A3(n7660), .A4(n7622), .ZN(n55266)
         );
  NOR4_X1 U38068 ( .A1(n7625), .A2(n49872), .A3(n7661), .A4(n7623), .ZN(n55265) );
  NOR4_X1 U38069 ( .A1(n7626), .A2(DRAM_ADDR[0]), .A3(n53648), .A4(
        DRAM_ADDR[3]), .ZN(n55264) );
  NAND4_X1 U38070 ( .A1(n55267), .A2(n55266), .A3(n55265), .A4(n55264), .ZN(
        n55274) );
  NAND4_X1 U38071 ( .A1(n49815), .A2(n49811), .A3(n3248), .A4(n49814), .ZN(
        n55271) );
  NAND4_X1 U38072 ( .A1(n3273), .A2(n49810), .A3(n49842), .A4(n49839), .ZN(
        n55270) );
  NAND4_X1 U38073 ( .A1(n49834), .A2(n49843), .A3(n3249), .A4(n49809), .ZN(
        n55269) );
  NAND4_X1 U38074 ( .A1(n49832), .A2(n49844), .A3(n49808), .A4(n3247), .ZN(
        n55268) );
  NOR4_X1 U38075 ( .A1(n55271), .A2(n55270), .A3(n55269), .A4(n55268), .ZN(
        n55272) );
  NAND2_X1 U38076 ( .A1(n55276), .A2(n55272), .ZN(n55273) );
  OAI22_X1 U38077 ( .A1(n55276), .A2(n55275), .B1(n55274), .B2(n55273), .ZN(
        n55277) );
  AOI21_X1 U38078 ( .B1(n55279), .B2(n55278), .A(n55277), .ZN(n55281) );
  OAI21_X1 U38079 ( .B1(w_EQ_COND), .B2(n55281), .A(w_JUMP_EN), .ZN(n55280) );
  OAI22_X1 U38080 ( .A1(n3248), .A2(n55284), .B1(n53711), .B2(n55283), .ZN(
        n5089) );
  OAI22_X1 U38081 ( .A1(n53671), .A2(n55284), .B1(n55283), .B2(n53730), .ZN(
        n5090) );
  OAI22_X1 U38082 ( .A1(n53668), .A2(n55284), .B1(n55283), .B2(n53731), .ZN(
        n5091) );
  OAI22_X1 U38083 ( .A1(n53660), .A2(n55284), .B1(n55283), .B2(n53732), .ZN(
        n5092) );
  OAI22_X1 U38084 ( .A1(n53670), .A2(n55284), .B1(n55283), .B2(n53733), .ZN(
        n5093) );
  OAI22_X1 U38085 ( .A1(n49808), .A2(n55284), .B1(n53712), .B2(n55283), .ZN(
        n5094) );
  OAI22_X1 U38086 ( .A1(n49838), .A2(n55284), .B1(n53713), .B2(n55283), .ZN(
        n5095) );
  OAI22_X1 U38087 ( .A1(n49832), .A2(n55284), .B1(n53714), .B2(n55283), .ZN(
        n5096) );
  OAI22_X1 U38088 ( .A1(n3249), .A2(n55284), .B1(n53715), .B2(n55283), .ZN(
        n5097) );
  OAI22_X1 U38089 ( .A1(n49815), .A2(n55284), .B1(n53716), .B2(n55283), .ZN(
        n5098) );
  OAI22_X1 U38090 ( .A1(n53665), .A2(n55284), .B1(n55283), .B2(n53734), .ZN(
        n5099) );
  OAI22_X1 U38091 ( .A1(n49834), .A2(n55284), .B1(n53717), .B2(n55283), .ZN(
        n5100) );
  OAI22_X1 U38092 ( .A1(n3273), .A2(n55284), .B1(n53718), .B2(n55283), .ZN(
        n5101) );
  OAI22_X1 U38093 ( .A1(n3247), .A2(n55284), .B1(n53719), .B2(n55283), .ZN(
        n5102) );
  OAI22_X1 U38094 ( .A1(n49844), .A2(n55284), .B1(n53720), .B2(n55283), .ZN(
        n5103) );
  OAI22_X1 U38095 ( .A1(n49814), .A2(n55284), .B1(n53721), .B2(n55283), .ZN(
        n5104) );
  OAI22_X1 U38096 ( .A1(n49809), .A2(n55284), .B1(n53722), .B2(n55283), .ZN(
        n5105) );
  OAI22_X1 U38097 ( .A1(n49810), .A2(n55284), .B1(n53723), .B2(n55283), .ZN(
        n5106) );
  OAI22_X1 U38098 ( .A1(n53669), .A2(n55284), .B1(n55283), .B2(n53735), .ZN(
        n5107) );
  OAI22_X1 U38099 ( .A1(n49839), .A2(n55284), .B1(n53724), .B2(n55283), .ZN(
        n5108) );
  OAI22_X1 U38100 ( .A1(n53663), .A2(n55284), .B1(n55283), .B2(n53736), .ZN(
        n5109) );
  OAI22_X1 U38101 ( .A1(n53672), .A2(n55284), .B1(n55283), .B2(n53737), .ZN(
        n5110) );
  OAI22_X1 U38102 ( .A1(n53667), .A2(n55284), .B1(n55283), .B2(n53738), .ZN(
        n5111) );
  OAI22_X1 U38103 ( .A1(n53666), .A2(n55284), .B1(n55283), .B2(n53739), .ZN(
        n5112) );
  OAI22_X1 U38104 ( .A1(n3260), .A2(n55284), .B1(n53725), .B2(n55283), .ZN(
        n5113) );
  OAI22_X1 U38105 ( .A1(n49843), .A2(n55284), .B1(n53726), .B2(n55283), .ZN(
        n5114) );
  OAI22_X1 U38106 ( .A1(n53661), .A2(n55284), .B1(n55283), .B2(n53740), .ZN(
        n5115) );
  OAI22_X1 U38107 ( .A1(n49842), .A2(n55284), .B1(n53727), .B2(n55283), .ZN(
        n5116) );
  OAI22_X1 U38108 ( .A1(n53664), .A2(n55284), .B1(n55283), .B2(n53741), .ZN(
        n5117) );
  OAI22_X1 U38109 ( .A1(n3254), .A2(n55284), .B1(n53728), .B2(n55283), .ZN(
        n5118) );
  OAI22_X1 U38110 ( .A1(n49811), .A2(n55284), .B1(n53729), .B2(n55283), .ZN(
        n5119) );
  OAI22_X1 U38111 ( .A1(n53662), .A2(n55284), .B1(n55283), .B2(n53742), .ZN(
        n5120) );
  AND2_X1 U38112 ( .A1(n53814), .A2(IRAM_DATA[29]), .ZN(n5121) );
  AND2_X1 U38113 ( .A1(n53813), .A2(IRAM_DATA[25]), .ZN(n5122) );
  AND2_X1 U38114 ( .A1(n53813), .A2(IRAM_DATA[23]), .ZN(n5124) );
  AND2_X1 U38115 ( .A1(n53813), .A2(IRAM_DATA[28]), .ZN(n5125) );
  AND2_X1 U38116 ( .A1(n53813), .A2(IRAM_DATA[22]), .ZN(n5126) );
  AND2_X1 U38117 ( .A1(n53814), .A2(IRAM_DATA[24]), .ZN(n5127) );
  AND2_X1 U38118 ( .A1(n55354), .A2(IRAM_DATA[21]), .ZN(n5128) );
  AND2_X1 U38119 ( .A1(n53813), .A2(IRAM_DATA[0]), .ZN(n5129) );
  AND2_X1 U38120 ( .A1(n53813), .A2(IRAM_DATA[1]), .ZN(n5130) );
  AND2_X1 U38121 ( .A1(n53814), .A2(IRAM_DATA[2]), .ZN(n5131) );
  AND2_X1 U38122 ( .A1(n53813), .A2(IRAM_DATA[3]), .ZN(n5132) );
  AND2_X1 U38123 ( .A1(n53813), .A2(IRAM_DATA[4]), .ZN(n5133) );
  AND2_X1 U38124 ( .A1(n53813), .A2(IRAM_DATA[5]), .ZN(n5134) );
  AND2_X1 U38125 ( .A1(n53813), .A2(IRAM_DATA[6]), .ZN(n5135) );
  AND2_X1 U38126 ( .A1(n53813), .A2(IRAM_DATA[7]), .ZN(n5136) );
  AND2_X1 U38127 ( .A1(n53813), .A2(IRAM_DATA[8]), .ZN(n5137) );
  AND2_X1 U38128 ( .A1(n53813), .A2(IRAM_DATA[9]), .ZN(n5138) );
  AND2_X1 U38129 ( .A1(n53813), .A2(IRAM_DATA[10]), .ZN(n5139) );
  AND2_X1 U38130 ( .A1(n53813), .A2(IRAM_DATA[11]), .ZN(n5140) );
  AND2_X1 U38131 ( .A1(n53813), .A2(IRAM_DATA[12]), .ZN(n5141) );
  AND2_X1 U38132 ( .A1(n53813), .A2(IRAM_DATA[13]), .ZN(n5142) );
  AND2_X1 U38133 ( .A1(n53813), .A2(IRAM_DATA[14]), .ZN(n5143) );
  AND2_X1 U38134 ( .A1(n53813), .A2(IRAM_DATA[15]), .ZN(n5144) );
  AND2_X1 U38135 ( .A1(n53814), .A2(IRAM_DATA[16]), .ZN(n5145) );
  AND2_X1 U38136 ( .A1(n53814), .A2(IRAM_DATA[17]), .ZN(n5146) );
  AND2_X1 U38137 ( .A1(n53814), .A2(IRAM_DATA[18]), .ZN(n5147) );
  AND2_X1 U38138 ( .A1(n53814), .A2(IRAM_DATA[19]), .ZN(n5148) );
  AND2_X1 U38139 ( .A1(n53814), .A2(IRAM_DATA[20]), .ZN(n5149) );
  AND2_X1 U38140 ( .A1(n53814), .A2(IRAM_DATA[26]), .ZN(n5150) );
  AND2_X1 U38141 ( .A1(n53814), .A2(IRAM_DATA[27]), .ZN(n5151) );
  AND2_X1 U38142 ( .A1(n53814), .A2(IRAM_DATA[30]), .ZN(n5152) );
  NAND2_X1 U38143 ( .A1(n55361), .A2(w_PC_OUT[27]), .ZN(n55360) );
  NAND2_X1 U38144 ( .A1(n55359), .A2(w_PC_OUT[29]), .ZN(n55327) );
  OAI21_X1 U38145 ( .B1(n55288), .B2(w_PC_OUT[31]), .A(n53813), .ZN(n55285) );
  AOI21_X1 U38146 ( .B1(n55288), .B2(w_PC_OUT[31]), .A(n55285), .ZN(n5153) );
  NOR2_X1 U38147 ( .A1(n7226), .A2(n53815), .ZN(n5154) );
  NOR2_X1 U38148 ( .A1(n7227), .A2(n53815), .ZN(n5155) );
  AND2_X1 U38149 ( .A1(n53814), .A2(n7228), .ZN(n5156) );
  NOR2_X1 U38150 ( .A1(n7228), .A2(n7229), .ZN(n55297) );
  INV_X1 U38151 ( .A(n55297), .ZN(n55287) );
  AOI211_X1 U38152 ( .C1(n3270), .C2(n55287), .A(n55286), .B(n53815), .ZN(
        n5158) );
  AOI211_X1 U38153 ( .C1(n49845), .C2(n55327), .A(n55288), .B(n53815), .ZN(
        n5184) );
  AND2_X1 U38154 ( .A1(RST), .A2(\DP/RegA_IN[0] ), .ZN(n5186) );
  AND2_X1 U38155 ( .A1(RST), .A2(\DP/RegA_IN[1] ), .ZN(n5187) );
  AND2_X1 U38156 ( .A1(RST), .A2(\DP/RegA_IN[2] ), .ZN(n5188) );
  AND2_X1 U38157 ( .A1(RST), .A2(\DP/RegA_IN[3] ), .ZN(n5189) );
  AND2_X1 U38158 ( .A1(RST), .A2(\DP/RegA_IN[4] ), .ZN(n5190) );
  AND2_X1 U38159 ( .A1(RST), .A2(\DP/RegA_IN[5] ), .ZN(n5191) );
  AND2_X1 U38160 ( .A1(RST), .A2(\DP/RegA_IN[6] ), .ZN(n5192) );
  AND2_X1 U38161 ( .A1(RST), .A2(\DP/RegA_IN[7] ), .ZN(n5193) );
  AND2_X1 U38162 ( .A1(RST), .A2(\DP/RegA_IN[8] ), .ZN(n5194) );
  AND2_X1 U38163 ( .A1(RST), .A2(\DP/RegA_IN[9] ), .ZN(n5195) );
  AND2_X1 U38164 ( .A1(RST), .A2(\DP/RegA_IN[10] ), .ZN(n5196) );
  AND2_X1 U38165 ( .A1(RST), .A2(\DP/RegA_IN[11] ), .ZN(n5197) );
  AND2_X1 U38166 ( .A1(RST), .A2(\DP/RegA_IN[12] ), .ZN(n5198) );
  AND2_X1 U38167 ( .A1(RST), .A2(\DP/RegA_IN[13] ), .ZN(n5199) );
  AND2_X1 U38168 ( .A1(RST), .A2(\DP/RegA_IN[14] ), .ZN(n5200) );
  AND2_X1 U38169 ( .A1(RST), .A2(\DP/RegA_IN[15] ), .ZN(n5201) );
  AND2_X1 U38170 ( .A1(RST), .A2(\DP/RegA_IN[16] ), .ZN(n5202) );
  AND2_X1 U38171 ( .A1(RST), .A2(\DP/RegA_IN[17] ), .ZN(n5203) );
  AND2_X1 U38172 ( .A1(RST), .A2(\DP/RegA_IN[18] ), .ZN(n5204) );
  AND2_X1 U38173 ( .A1(RST), .A2(\DP/RegA_IN[19] ), .ZN(n5205) );
  AND2_X1 U38174 ( .A1(RST), .A2(\DP/RegA_IN[20] ), .ZN(n5206) );
  AND2_X1 U38175 ( .A1(RST), .A2(\DP/RegA_IN[21] ), .ZN(n5207) );
  AND2_X1 U38176 ( .A1(RST), .A2(\DP/RegA_IN[22] ), .ZN(n5208) );
  AND2_X1 U38177 ( .A1(RST), .A2(\DP/RegA_IN[23] ), .ZN(n5209) );
  AND2_X1 U38178 ( .A1(RST), .A2(\DP/RegA_IN[24] ), .ZN(n5210) );
  AND2_X1 U38179 ( .A1(RST), .A2(\DP/RegA_IN[25] ), .ZN(n5211) );
  AND2_X1 U38180 ( .A1(RST), .A2(\DP/RegA_IN[26] ), .ZN(n5212) );
  AND2_X1 U38181 ( .A1(RST), .A2(\DP/RegA_IN[27] ), .ZN(n5213) );
  AND2_X1 U38182 ( .A1(RST), .A2(\DP/RegA_IN[28] ), .ZN(n5214) );
  AND2_X1 U38183 ( .A1(RST), .A2(\DP/RegA_IN[29] ), .ZN(n5215) );
  AND2_X1 U38184 ( .A1(RST), .A2(\DP/RegA_IN[30] ), .ZN(n5216) );
  AND2_X1 U38185 ( .A1(RST), .A2(\DP/RegA_IN[31] ), .ZN(n5217) );
  AND2_X1 U38186 ( .A1(RST), .A2(\DP/RegB_IN[0] ), .ZN(n5218) );
  AND2_X1 U38187 ( .A1(RST), .A2(\DP/RegB_IN[1] ), .ZN(n5219) );
  AND2_X1 U38188 ( .A1(RST), .A2(\DP/RegB_IN[2] ), .ZN(n5220) );
  AND2_X1 U38189 ( .A1(RST), .A2(\DP/RegB_IN[3] ), .ZN(n5221) );
  AND2_X1 U38190 ( .A1(RST), .A2(\DP/RegB_IN[4] ), .ZN(n5222) );
  AND2_X1 U38191 ( .A1(RST), .A2(\DP/RegB_IN[5] ), .ZN(n5223) );
  AND2_X1 U38192 ( .A1(RST), .A2(\DP/RegB_IN[6] ), .ZN(n5224) );
  AND2_X1 U38193 ( .A1(RST), .A2(\DP/RegB_IN[7] ), .ZN(n5225) );
  AND2_X1 U38194 ( .A1(RST), .A2(\DP/RegB_IN[8] ), .ZN(n5226) );
  AND2_X1 U38195 ( .A1(RST), .A2(\DP/RegB_IN[9] ), .ZN(n5227) );
  AND2_X1 U38196 ( .A1(RST), .A2(\DP/RegB_IN[10] ), .ZN(n5228) );
  AND2_X1 U38197 ( .A1(RST), .A2(\DP/RegB_IN[11] ), .ZN(n5229) );
  AND2_X1 U38198 ( .A1(RST), .A2(\DP/RegB_IN[12] ), .ZN(n5230) );
  AND2_X1 U38199 ( .A1(RST), .A2(\DP/RegB_IN[13] ), .ZN(n5231) );
  AND2_X1 U38200 ( .A1(RST), .A2(\DP/RegB_IN[14] ), .ZN(n5232) );
  AND2_X1 U38201 ( .A1(RST), .A2(\DP/RegB_IN[15] ), .ZN(n5233) );
  AND2_X1 U38202 ( .A1(RST), .A2(\DP/RegB_IN[16] ), .ZN(n5234) );
  AND2_X1 U38203 ( .A1(RST), .A2(\DP/RegB_IN[17] ), .ZN(n5235) );
  AND2_X1 U38204 ( .A1(RST), .A2(\DP/RegB_IN[18] ), .ZN(n5236) );
  AND2_X1 U38205 ( .A1(RST), .A2(\DP/RegB_IN[19] ), .ZN(n5237) );
  AND2_X1 U38206 ( .A1(RST), .A2(\DP/RegB_IN[20] ), .ZN(n5238) );
  AND2_X1 U38207 ( .A1(RST), .A2(\DP/RegB_IN[21] ), .ZN(n5239) );
  AND2_X1 U38208 ( .A1(RST), .A2(\DP/RegB_IN[22] ), .ZN(n5240) );
  AND2_X1 U38209 ( .A1(RST), .A2(\DP/RegB_IN[23] ), .ZN(n5241) );
  AND2_X1 U38210 ( .A1(RST), .A2(\DP/RegB_IN[24] ), .ZN(n5242) );
  AND2_X1 U38211 ( .A1(RST), .A2(\DP/RegB_IN[25] ), .ZN(n5243) );
  AND2_X1 U38212 ( .A1(RST), .A2(\DP/RegB_IN[26] ), .ZN(n5244) );
  AND2_X1 U38213 ( .A1(RST), .A2(\DP/RegB_IN[27] ), .ZN(n5245) );
  AND2_X1 U38214 ( .A1(RST), .A2(\DP/RegB_IN[28] ), .ZN(n5246) );
  AND2_X1 U38215 ( .A1(RST), .A2(\DP/RegB_IN[29] ), .ZN(n5247) );
  AND2_X1 U38216 ( .A1(RST), .A2(\DP/RegB_IN[30] ), .ZN(n5248) );
  AND2_X1 U38217 ( .A1(RST), .A2(\DP/RegB_IN[31] ), .ZN(n5249) );
  NOR2_X1 U38218 ( .A1(n49849), .A2(n55291), .ZN(n5250) );
  NOR2_X1 U38219 ( .A1(n55291), .A2(n53686), .ZN(n5251) );
  NOR2_X1 U38220 ( .A1(n7564), .A2(n55291), .ZN(n5252) );
  NOR2_X1 U38221 ( .A1(n55291), .A2(n53649), .ZN(n5253) );
  NOR2_X1 U38222 ( .A1(n7616), .A2(n55291), .ZN(n5254) );
  NOR2_X1 U38223 ( .A1(n55291), .A2(n53687), .ZN(n5255) );
  NOR2_X1 U38224 ( .A1(n55291), .A2(n53746), .ZN(n5256) );
  NOR2_X1 U38225 ( .A1(n49908), .A2(n55291), .ZN(n5257) );
  NOR2_X1 U38226 ( .A1(n49909), .A2(n55291), .ZN(n5258) );
  NOR2_X1 U38227 ( .A1(n55291), .A2(n53747), .ZN(n5259) );
  NOR2_X1 U38228 ( .A1(n55291), .A2(n53745), .ZN(n5260) );
  NOR2_X1 U38229 ( .A1(n55291), .A2(n53748), .ZN(n5261) );
  NOR2_X1 U38230 ( .A1(n55291), .A2(n53749), .ZN(n5262) );
  NOR2_X1 U38231 ( .A1(n55291), .A2(n53750), .ZN(n5263) );
  NOR2_X1 U38232 ( .A1(n55291), .A2(n53751), .ZN(n5264) );
  NOR2_X1 U38233 ( .A1(n7667), .A2(n55291), .ZN(n5265) );
  OAI21_X1 U38234 ( .B1(n53695), .B2(n55293), .A(n55292), .ZN(n5266) );
  OAI21_X1 U38235 ( .B1(n53696), .B2(n55293), .A(n55292), .ZN(n5267) );
  OAI21_X1 U38236 ( .B1(n53697), .B2(n55293), .A(n55292), .ZN(n5268) );
  OAI21_X1 U38237 ( .B1(n53698), .B2(n55293), .A(n55292), .ZN(n5269) );
  OAI21_X1 U38238 ( .B1(n53699), .B2(n55293), .A(n55292), .ZN(n5270) );
  OAI21_X1 U38239 ( .B1(\IR/n57 ), .B2(n55293), .A(n55292), .ZN(n5271) );
  OAI21_X1 U38240 ( .B1(\IR/n58 ), .B2(n55293), .A(n55292), .ZN(n5272) );
  OAI21_X1 U38241 ( .B1(\IR/n59 ), .B2(n55293), .A(n55292), .ZN(n5273) );
  OAI21_X1 U38242 ( .B1(\IR/n60 ), .B2(n55293), .A(n55292), .ZN(n5274) );
  AND2_X1 U38243 ( .A1(n55294), .A2(n53562), .ZN(n5275) );
  AND2_X1 U38244 ( .A1(n55294), .A2(n53563), .ZN(n5276) );
  AND2_X1 U38245 ( .A1(n55294), .A2(n53564), .ZN(n5277) );
  AND2_X1 U38246 ( .A1(n55294), .A2(n53565), .ZN(n5278) );
  AND2_X1 U38247 ( .A1(n55294), .A2(n53566), .ZN(n5279) );
  AND2_X1 U38248 ( .A1(n55294), .A2(n53567), .ZN(n5280) );
  AND2_X1 U38249 ( .A1(n55294), .A2(n53568), .ZN(n5281) );
  AND2_X1 U38250 ( .A1(n55294), .A2(n53569), .ZN(n5282) );
  AND2_X1 U38251 ( .A1(n55294), .A2(n53570), .ZN(n5283) );
  AND2_X1 U38252 ( .A1(n55294), .A2(n53571), .ZN(n5284) );
  AND2_X1 U38253 ( .A1(n53811), .A2(n53572), .ZN(n5285) );
  AND2_X1 U38254 ( .A1(n53811), .A2(n53573), .ZN(n5286) );
  AND2_X1 U38255 ( .A1(n53811), .A2(n53574), .ZN(n5287) );
  AND2_X1 U38256 ( .A1(n53811), .A2(n53575), .ZN(n5288) );
  AND2_X1 U38257 ( .A1(n53811), .A2(n53576), .ZN(n5289) );
  AND2_X1 U38258 ( .A1(n53811), .A2(n53577), .ZN(n5290) );
  AND2_X1 U38259 ( .A1(n53811), .A2(n53578), .ZN(n5291) );
  AND2_X1 U38260 ( .A1(n53811), .A2(n53579), .ZN(n5292) );
  AND2_X1 U38261 ( .A1(n53811), .A2(n53580), .ZN(n5293) );
  AND2_X1 U38262 ( .A1(n53811), .A2(n53581), .ZN(n5294) );
  AND2_X1 U38263 ( .A1(n53811), .A2(n53582), .ZN(n5295) );
  AND2_X1 U38264 ( .A1(n53811), .A2(n53583), .ZN(n5296) );
  AND2_X1 U38265 ( .A1(n53811), .A2(n53584), .ZN(n5297) );
  AND2_X1 U38266 ( .A1(n53811), .A2(n53585), .ZN(n5298) );
  AND2_X1 U38267 ( .A1(n53811), .A2(n53586), .ZN(n5299) );
  AND2_X1 U38268 ( .A1(n53811), .A2(n53587), .ZN(n5300) );
  AND2_X1 U38269 ( .A1(n53811), .A2(n53588), .ZN(n5301) );
  AND2_X1 U38270 ( .A1(n53811), .A2(n53589), .ZN(n5302) );
  AND2_X1 U38271 ( .A1(n53811), .A2(n53590), .ZN(n5303) );
  AND2_X1 U38272 ( .A1(n53811), .A2(n53591), .ZN(n5304) );
  AND2_X1 U38273 ( .A1(n55294), .A2(n53592), .ZN(n5305) );
  AND2_X1 U38274 ( .A1(n55294), .A2(n53593), .ZN(n5306) );
  AOI211_X1 U38275 ( .C1(n7230), .C2(n55296), .A(n55295), .B(n53815), .ZN(
        n7478) );
  AOI211_X1 U38276 ( .C1(n7228), .C2(n7229), .A(n55297), .B(n53815), .ZN(n7489) );
  NAND2_X1 U38277 ( .A1(RST), .A2(n3018), .ZN(n897) );
  OR2_X1 U38278 ( .A1(n55299), .A2(n55298), .ZN(n55301) );
  AOI211_X1 U38279 ( .C1(\intadd_7/SUM[1] ), .C2(n55301), .A(\intadd_6/A[0] ), 
        .B(n55300), .ZN(n55305) );
  NAND2_X1 U38280 ( .A1(n53809), .A2(\DP/ALU0/S_B_LOGIC[4] ), .ZN(n55302) );
  OAI22_X1 U38281 ( .A1(\intadd_0/SUM[3] ), .A2(n55303), .B1(
        \DP/ALU0/s_A_LOGIC[4] ), .B2(n55302), .ZN(n55304) );
  AOI211_X1 U38282 ( .C1(n55307), .C2(n55306), .A(n55305), .B(n55304), .ZN(
        n55311) );
  INV_X1 U38283 ( .A(\DP/ALU0/S_B_LOGIC[4] ), .ZN(n55309) );
  OAI221_X1 U38284 ( .B1(\DP/ALU0/S_B_LOGIC[4] ), .B2(n53809), .C1(n55309), 
        .C2(n55308), .A(\DP/ALU0/s_A_LOGIC[4] ), .ZN(n55310) );
  OAI211_X1 U38285 ( .C1(n55313), .C2(n55312), .A(n55311), .B(n55310), .ZN(
        n9277) );
  OAI21_X1 U38286 ( .B1(n55316), .B2(n55315), .A(n55314), .ZN(n53612) );
  OAI211_X1 U38287 ( .C1(n55317), .C2(w_PC_OUT[13]), .A(n53814), .B(n55348), 
        .ZN(n55318) );
  INV_X1 U38288 ( .A(n55318), .ZN(n53610) );
  OAI211_X1 U38289 ( .C1(n55347), .C2(w_PC_OUT[15]), .A(n53813), .B(n55350), 
        .ZN(n55319) );
  INV_X1 U38290 ( .A(n55319), .ZN(n53609) );
  OAI211_X1 U38291 ( .C1(n55349), .C2(w_PC_OUT[17]), .A(n53814), .B(n55352), 
        .ZN(n55320) );
  INV_X1 U38292 ( .A(n55320), .ZN(n53608) );
  OAI211_X1 U38293 ( .C1(n55351), .C2(w_PC_OUT[19]), .A(n53813), .B(n55321), 
        .ZN(n55322) );
  INV_X1 U38294 ( .A(n55322), .ZN(n53607) );
  OAI211_X1 U38295 ( .C1(n55323), .C2(w_PC_OUT[23]), .A(n53813), .B(n55358), 
        .ZN(n55324) );
  INV_X1 U38296 ( .A(n55324), .ZN(n53606) );
  OAI211_X1 U38297 ( .C1(n55357), .C2(w_PC_OUT[25]), .A(n53813), .B(n55362), 
        .ZN(n55325) );
  INV_X1 U38298 ( .A(n55325), .ZN(n53605) );
  OAI211_X1 U38299 ( .C1(n55361), .C2(w_PC_OUT[27]), .A(n53813), .B(n55360), 
        .ZN(n55326) );
  INV_X1 U38300 ( .A(n55326), .ZN(n53604) );
  OAI211_X1 U38301 ( .C1(n55359), .C2(w_PC_OUT[29]), .A(n53813), .B(n55327), 
        .ZN(n55328) );
  INV_X1 U38302 ( .A(n55328), .ZN(n53603) );
  INV_X1 U38303 ( .A(\DP/ALU0/s_A_ADDER[31] ), .ZN(n51803) );
  INV_X1 U38304 ( .A(\DP/ALU0/s_A_ADDER[30] ), .ZN(n51802) );
  INV_X1 U38305 ( .A(\DP/ALU0/s_A_ADDER[29] ), .ZN(n51801) );
  INV_X1 U38306 ( .A(\DP/ALU0/s_A_ADDER[28] ), .ZN(n51800) );
  INV_X1 U38307 ( .A(\DP/ALU0/s_A_ADDER[27] ), .ZN(n51799) );
  INV_X1 U38308 ( .A(\DP/ALU0/s_A_ADDER[26] ), .ZN(n51798) );
  INV_X1 U38309 ( .A(\DP/ALU0/s_A_ADDER[25] ), .ZN(n51797) );
  INV_X1 U38310 ( .A(\DP/ALU0/s_A_ADDER[24] ), .ZN(n51796) );
  INV_X1 U38311 ( .A(\DP/ALU0/s_A_ADDER[23] ), .ZN(n51795) );
  INV_X1 U38312 ( .A(\DP/ALU0/s_A_ADDER[22] ), .ZN(n51794) );
  INV_X1 U38313 ( .A(\DP/ALU0/s_A_ADDER[21] ), .ZN(n51793) );
  INV_X1 U38314 ( .A(\DP/ALU0/s_A_ADDER[20] ), .ZN(n51792) );
  INV_X1 U38315 ( .A(\DP/ALU0/s_A_ADDER[19] ), .ZN(n51791) );
  INV_X1 U38316 ( .A(\DP/ALU0/s_A_ADDER[18] ), .ZN(n51790) );
  INV_X1 U38317 ( .A(\DP/ALU0/s_A_ADDER[17] ), .ZN(n51789) );
  INV_X1 U38318 ( .A(\DP/ALU0/s_A_ADDER[16] ), .ZN(n51788) );
  INV_X1 U38319 ( .A(\DP/ALU0/s_A_ADDER[15] ), .ZN(n51787) );
  INV_X1 U38320 ( .A(\DP/ALU0/s_A_ADDER[14] ), .ZN(n51786) );
  INV_X1 U38321 ( .A(\DP/ALU0/s_A_ADDER[13] ), .ZN(n51785) );
  INV_X1 U38322 ( .A(\DP/ALU0/s_A_ADDER[12] ), .ZN(n51784) );
  INV_X1 U38323 ( .A(\DP/ALU0/s_A_ADDER[11] ), .ZN(n51783) );
  INV_X1 U38324 ( .A(\DP/ALU0/s_A_ADDER[10] ), .ZN(n51782) );
  INV_X1 U38325 ( .A(\DP/ALU0/s_A_ADDER[9] ), .ZN(n51781) );
  INV_X1 U38326 ( .A(\DP/ALU0/s_A_ADDER[8] ), .ZN(n51780) );
  INV_X1 U38327 ( .A(\DP/ALU0/s_A_ADDER[7] ), .ZN(n51779) );
  INV_X1 U38328 ( .A(\DP/ALU0/s_A_ADDER[6] ), .ZN(n51778) );
  INV_X1 U38329 ( .A(\DP/ALU0/s_A_ADDER[5] ), .ZN(n51777) );
  INV_X1 U38330 ( .A(\DP/ALU0/s_A_ADDER[4] ), .ZN(n51776) );
  INV_X1 U38331 ( .A(\DP/ALU0/s_A_ADDER[3] ), .ZN(n51775) );
  INV_X1 U38332 ( .A(\DP/ALU0/s_A_ADDER[2] ), .ZN(n51774) );
  INV_X1 U38333 ( .A(\DP/ALU0/s_A_ADDER[1] ), .ZN(n51773) );
  INV_X1 U38334 ( .A(\intadd_7/SUM[2] ), .ZN(n51699) );
  INV_X1 U38335 ( .A(\intadd_7/SUM[3] ), .ZN(n51698) );
  INV_X1 U38336 ( .A(\intadd_7/SUM[4] ), .ZN(n51697) );
  INV_X1 U38337 ( .A(\intadd_6/SUM[2] ), .ZN(n51696) );
  INV_X1 U38338 ( .A(\intadd_7/SUM[5] ), .ZN(n51695) );
  INV_X1 U38339 ( .A(\intadd_6/SUM[3] ), .ZN(n51694) );
  INV_X1 U38340 ( .A(\intadd_7/SUM[6] ), .ZN(n51693) );
  INV_X1 U38341 ( .A(\intadd_6/SUM[4] ), .ZN(n51692) );
  INV_X1 U38342 ( .A(\intadd_5/SUM[2] ), .ZN(n51691) );
  INV_X1 U38343 ( .A(\intadd_7/SUM[7] ), .ZN(n51690) );
  INV_X1 U38344 ( .A(\intadd_6/SUM[5] ), .ZN(n51689) );
  INV_X1 U38345 ( .A(\intadd_5/SUM[3] ), .ZN(n51688) );
  INV_X1 U38346 ( .A(\intadd_7/SUM[8] ), .ZN(n51687) );
  INV_X1 U38347 ( .A(\intadd_6/SUM[6] ), .ZN(n51686) );
  INV_X1 U38348 ( .A(\intadd_5/SUM[4] ), .ZN(n51685) );
  INV_X1 U38349 ( .A(\intadd_4/SUM[2] ), .ZN(n51684) );
  INV_X1 U38350 ( .A(\intadd_7/SUM[9] ), .ZN(n51683) );
  INV_X1 U38351 ( .A(\intadd_6/SUM[7] ), .ZN(n51682) );
  INV_X1 U38352 ( .A(\intadd_5/SUM[5] ), .ZN(n51681) );
  INV_X1 U38353 ( .A(\intadd_4/SUM[3] ), .ZN(n51680) );
  INV_X1 U38354 ( .A(\intadd_7/SUM[10] ), .ZN(n51678) );
  INV_X1 U38355 ( .A(\intadd_6/SUM[8] ), .ZN(n51677) );
  INV_X1 U38356 ( .A(\intadd_5/SUM[6] ), .ZN(n51676) );
  INV_X1 U38357 ( .A(\intadd_4/SUM[4] ), .ZN(n51675) );
  INV_X1 U38358 ( .A(\intadd_7/SUM[11] ), .ZN(n51674) );
  INV_X1 U38359 ( .A(\intadd_6/SUM[9] ), .ZN(n51673) );
  INV_X1 U38360 ( .A(\intadd_5/SUM[7] ), .ZN(n51672) );
  INV_X1 U38361 ( .A(\intadd_4/SUM[5] ), .ZN(n51671) );
  INV_X1 U38362 ( .A(\intadd_7/SUM[12] ), .ZN(n51670) );
  INV_X1 U38363 ( .A(\intadd_6/SUM[10] ), .ZN(n51669) );
  INV_X1 U38364 ( .A(\intadd_5/SUM[8] ), .ZN(n51668) );
  INV_X1 U38365 ( .A(\intadd_4/SUM[6] ), .ZN(n51667) );
  INV_X1 U38366 ( .A(\intadd_2/SUM[2] ), .ZN(n51666) );
  INV_X1 U38367 ( .A(\intadd_6/SUM[11] ), .ZN(n51665) );
  INV_X1 U38368 ( .A(\intadd_5/SUM[9] ), .ZN(n51664) );
  INV_X1 U38369 ( .A(\intadd_4/SUM[7] ), .ZN(n51663) );
  INV_X1 U38370 ( .A(\intadd_2/SUM[3] ), .ZN(n51662) );
  INV_X1 U38371 ( .A(\intadd_6/SUM[12] ), .ZN(n51661) );
  INV_X1 U38372 ( .A(\intadd_5/SUM[10] ), .ZN(n51660) );
  INV_X1 U38373 ( .A(\intadd_4/SUM[8] ), .ZN(n51659) );
  INV_X1 U38374 ( .A(\intadd_2/SUM[4] ), .ZN(n51658) );
  INV_X1 U38375 ( .A(\intadd_5/SUM[11] ), .ZN(n51656) );
  INV_X1 U38376 ( .A(\intadd_4/SUM[9] ), .ZN(n51655) );
  INV_X1 U38377 ( .A(\intadd_2/SUM[5] ), .ZN(n51654) );
  INV_X1 U38378 ( .A(\intadd_5/SUM[12] ), .ZN(n51653) );
  INV_X1 U38379 ( .A(\intadd_4/SUM[10] ), .ZN(n51652) );
  INV_X1 U38380 ( .A(\intadd_2/SUM[6] ), .ZN(n51651) );
  INV_X1 U38381 ( .A(\intadd_4/SUM[11] ), .ZN(n51649) );
  INV_X1 U38382 ( .A(\intadd_2/SUM[7] ), .ZN(n51648) );
  INV_X1 U38383 ( .A(\intadd_4/SUM[12] ), .ZN(n51647) );
  INV_X1 U38384 ( .A(\intadd_2/SUM[8] ), .ZN(n51646) );
  INV_X1 U38385 ( .A(\intadd_2/SUM[9] ), .ZN(n51644) );
  INV_X1 U38386 ( .A(\intadd_2/SUM[10] ), .ZN(n51643) );
  INV_X1 U38387 ( .A(\intadd_2/SUM[11] ), .ZN(n51642) );
  INV_X1 U38388 ( .A(\intadd_2/SUM[12] ), .ZN(n51641) );
  AOI21_X1 U38389 ( .B1(n53414), .B2(n55333), .A(n55332), .ZN(n55335) );
  MUX2_X1 U38390 ( .A(n55335), .B(n55334), .S(n53650), .Z(n51623) );
  OAI22_X1 U38391 ( .A1(n53705), .A2(n55336), .B1(n49938), .B2(n53650), .ZN(
        n55337) );
  INV_X1 U38392 ( .A(n55337), .ZN(n51619) );
  OAI211_X1 U38393 ( .C1(n55339), .C2(w_PC_OUT[7]), .A(n53813), .B(n55338), 
        .ZN(n55340) );
  INV_X1 U38394 ( .A(n55340), .ZN(n51537) );
  OAI211_X1 U38395 ( .C1(n55342), .C2(w_PC_OUT[9]), .A(n53813), .B(n55341), 
        .ZN(n55343) );
  INV_X1 U38396 ( .A(n55343), .ZN(n51536) );
  OAI211_X1 U38397 ( .C1(n55345), .C2(w_PC_OUT[11]), .A(n53813), .B(n55344), 
        .ZN(n55346) );
  INV_X1 U38398 ( .A(n55346), .ZN(n51535) );
  AOI211_X1 U38399 ( .C1(n55348), .C2(n53675), .A(n55347), .B(n53815), .ZN(
        n51533) );
  AOI211_X1 U38400 ( .C1(n55350), .C2(n53690), .A(n55349), .B(n53815), .ZN(
        n51532) );
  AOI211_X1 U38401 ( .C1(n55352), .C2(n53691), .A(n55351), .B(n53815), .ZN(
        n51531) );
  OAI211_X1 U38402 ( .C1(n55355), .C2(w_PC_OUT[21]), .A(n53813), .B(n55353), 
        .ZN(n55356) );
  INV_X1 U38403 ( .A(n55356), .ZN(n51529) );
  AOI211_X1 U38404 ( .C1(n55358), .C2(n53700), .A(n55357), .B(n53815), .ZN(
        n51527) );
  AOI211_X1 U38405 ( .C1(n55360), .C2(n53676), .A(n55359), .B(n53815), .ZN(
        n51525) );
  AOI211_X1 U38406 ( .C1(n55362), .C2(n53674), .A(n55361), .B(n53815), .ZN(
        n51524) );
endmodule


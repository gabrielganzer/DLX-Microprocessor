
module REGISTER_GENERIC_WIDTH32_0 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n96, n97, n98, n99, n102, n44, n69, n34, n35, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292;

  DFF_X1 \DOUT_reg[7]  ( .D(n70), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n71), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[3]  ( .D(n74), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[31]  ( .D(n75), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[25]  ( .D(n82), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[8]  ( .D(n69), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[11]  ( .D(n97), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  DFF_X1 \DOUT_reg[18]  ( .D(n90), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[20]  ( .D(n87), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[27]  ( .D(n80), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[29]  ( .D(n78), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[24]  ( .D(n83), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n84), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[13]  ( .D(n102), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[15]  ( .D(n93), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[12]  ( .D(n96), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[17]  ( .D(n91), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[2]  ( .D(n77), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n88), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[30]  ( .D(n76), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[28]  ( .D(n79), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[19]  ( .D(n89), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[5]  ( .D(n72), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[9]  ( .D(n68), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[26]  ( .D(n81), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[10]  ( .D(n98), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[22]  ( .D(n85), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[14]  ( .D(n94), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[21]  ( .D(n86), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[16]  ( .D(n92), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[4]  ( .D(n73), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  BUF_X1 U3 ( .A(n35), .Z(n256) );
  BUF_X1 U4 ( .A(n34), .Z(n259) );
  BUF_X1 U5 ( .A(n34), .Z(n257) );
  BUF_X1 U6 ( .A(n34), .Z(n258) );
  BUF_X1 U7 ( .A(n35), .Z(n255) );
  BUF_X1 U8 ( .A(n35), .Z(n254) );
  OAI22_X1 U9 ( .A1(n52), .A2(n259), .B1(n256), .B2(n275), .ZN(n92) );
  INV_X1 U10 ( .A(DIN[16]), .ZN(n275) );
  OAI22_X1 U11 ( .A1(n50), .A2(n259), .B1(n256), .B2(n277), .ZN(n94) );
  INV_X1 U12 ( .A(DIN[14]), .ZN(n277) );
  OAI22_X1 U13 ( .A1(n46), .A2(n259), .B1(n256), .B2(n281), .ZN(n98) );
  INV_X1 U14 ( .A(DIN[10]), .ZN(n281) );
  OAI22_X1 U15 ( .A1(n55), .A2(n258), .B1(n256), .B2(n272), .ZN(n89) );
  INV_X1 U16 ( .A(DIN[19]), .ZN(n272) );
  OAI22_X1 U17 ( .A1(n53), .A2(n259), .B1(n256), .B2(n274), .ZN(n91) );
  INV_X1 U18 ( .A(DIN[17]), .ZN(n274) );
  OAI22_X1 U19 ( .A1(n48), .A2(n259), .B1(n256), .B2(n279), .ZN(n96) );
  INV_X1 U20 ( .A(DIN[12]), .ZN(n279) );
  OAI22_X1 U21 ( .A1(n51), .A2(n259), .B1(n256), .B2(n276), .ZN(n93) );
  INV_X1 U22 ( .A(DIN[15]), .ZN(n276) );
  OAI22_X1 U23 ( .A1(n54), .A2(n259), .B1(n256), .B2(n273), .ZN(n90) );
  INV_X1 U24 ( .A(DIN[18]), .ZN(n273) );
  OAI22_X1 U25 ( .A1(n36), .A2(n259), .B1(n256), .B2(n291), .ZN(n99) );
  INV_X1 U26 ( .A(DIN[0]), .ZN(n291) );
  OAI22_X1 U27 ( .A1(n47), .A2(n259), .B1(n256), .B2(n280), .ZN(n97) );
  INV_X1 U28 ( .A(DIN[11]), .ZN(n280) );
  OAI22_X1 U29 ( .A1(n40), .A2(n257), .B1(n254), .B2(n287), .ZN(n73) );
  INV_X1 U30 ( .A(DIN[4]), .ZN(n287) );
  OAI22_X1 U31 ( .A1(n57), .A2(n258), .B1(n255), .B2(n270), .ZN(n86) );
  INV_X1 U32 ( .A(DIN[21]), .ZN(n270) );
  OAI22_X1 U33 ( .A1(n58), .A2(n258), .B1(n255), .B2(n269), .ZN(n85) );
  INV_X1 U34 ( .A(DIN[22]), .ZN(n269) );
  OAI22_X1 U35 ( .A1(n45), .A2(n257), .B1(n254), .B2(n282), .ZN(n68) );
  INV_X1 U36 ( .A(DIN[9]), .ZN(n282) );
  OAI22_X1 U37 ( .A1(n41), .A2(n257), .B1(n254), .B2(n286), .ZN(n72) );
  INV_X1 U38 ( .A(DIN[5]), .ZN(n286) );
  OAI22_X1 U39 ( .A1(n37), .A2(n258), .B1(n255), .B2(n290), .ZN(n88) );
  INV_X1 U40 ( .A(DIN[1]), .ZN(n290) );
  OAI22_X1 U41 ( .A1(n38), .A2(n257), .B1(n254), .B2(n289), .ZN(n77) );
  INV_X1 U42 ( .A(DIN[2]), .ZN(n289) );
  OAI22_X1 U43 ( .A1(n49), .A2(n257), .B1(n254), .B2(n278), .ZN(n102) );
  INV_X1 U44 ( .A(DIN[13]), .ZN(n278) );
  OAI22_X1 U45 ( .A1(n59), .A2(n258), .B1(n255), .B2(n268), .ZN(n84) );
  INV_X1 U46 ( .A(DIN[23]), .ZN(n268) );
  OAI22_X1 U47 ( .A1(n56), .A2(n258), .B1(n255), .B2(n271), .ZN(n87) );
  INV_X1 U48 ( .A(DIN[20]), .ZN(n271) );
  OAI22_X1 U49 ( .A1(n44), .A2(n257), .B1(n254), .B2(n283), .ZN(n69) );
  INV_X1 U50 ( .A(DIN[8]), .ZN(n283) );
  OAI22_X1 U51 ( .A1(n39), .A2(n257), .B1(n254), .B2(n288), .ZN(n74) );
  INV_X1 U52 ( .A(DIN[3]), .ZN(n288) );
  OAI22_X1 U53 ( .A1(n42), .A2(n257), .B1(n254), .B2(n285), .ZN(n71) );
  INV_X1 U54 ( .A(DIN[6]), .ZN(n285) );
  OAI22_X1 U55 ( .A1(n43), .A2(n257), .B1(n254), .B2(n284), .ZN(n70) );
  INV_X1 U56 ( .A(DIN[7]), .ZN(n284) );
  OAI22_X1 U57 ( .A1(n62), .A2(n258), .B1(n255), .B2(n265), .ZN(n81) );
  INV_X1 U58 ( .A(DIN[26]), .ZN(n265) );
  OAI22_X1 U59 ( .A1(n64), .A2(n258), .B1(n255), .B2(n263), .ZN(n79) );
  INV_X1 U60 ( .A(DIN[28]), .ZN(n263) );
  OAI22_X1 U61 ( .A1(n66), .A2(n257), .B1(n254), .B2(n261), .ZN(n76) );
  INV_X1 U62 ( .A(DIN[30]), .ZN(n261) );
  OAI22_X1 U63 ( .A1(n60), .A2(n258), .B1(n255), .B2(n267), .ZN(n83) );
  INV_X1 U64 ( .A(DIN[24]), .ZN(n267) );
  OAI22_X1 U65 ( .A1(n65), .A2(n258), .B1(n255), .B2(n262), .ZN(n78) );
  INV_X1 U66 ( .A(DIN[29]), .ZN(n262) );
  OAI22_X1 U67 ( .A1(n63), .A2(n258), .B1(n255), .B2(n264), .ZN(n80) );
  INV_X1 U68 ( .A(DIN[27]), .ZN(n264) );
  OAI22_X1 U69 ( .A1(n61), .A2(n258), .B1(n255), .B2(n266), .ZN(n82) );
  INV_X1 U70 ( .A(DIN[25]), .ZN(n266) );
  OAI22_X1 U71 ( .A1(n67), .A2(n257), .B1(n254), .B2(n260), .ZN(n75) );
  INV_X1 U72 ( .A(DIN[31]), .ZN(n260) );
  NAND2_X1 U73 ( .A1(RST), .A2(n257), .ZN(n35) );
  NAND2_X1 U74 ( .A1(n292), .A2(RST), .ZN(n34) );
  INV_X1 U75 ( .A(EN), .ZN(n292) );
endmodule


module REGISTER_GENERIC_WIDTH32_12 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294;

  DFF_X1 \DOUT_reg[30]  ( .D(n69), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[27]  ( .D(n72), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n73), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[20]  ( .D(n79), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n80), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n81), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n83), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n84), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n89), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n90), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n91), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n92), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n93), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n94), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n95), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n96), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n97), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n98), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  DFF_X1 \DOUT_reg[21]  ( .D(n78), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[24]  ( .D(n75), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[22]  ( .D(n77), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[28]  ( .D(n71), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[31]  ( .D(n68), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[25]  ( .D(n74), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[29]  ( .D(n70), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  BUF_X1 U3 ( .A(n35), .Z(n258) );
  BUF_X1 U4 ( .A(n34), .Z(n261) );
  BUF_X1 U5 ( .A(n34), .Z(n259) );
  BUF_X1 U6 ( .A(n34), .Z(n260) );
  BUF_X1 U7 ( .A(n35), .Z(n257) );
  BUF_X1 U8 ( .A(n35), .Z(n256) );
  OAI22_X1 U9 ( .A1(n36), .A2(n261), .B1(n258), .B2(n294), .ZN(n99) );
  INV_X1 U10 ( .A(DIN[0]), .ZN(n294) );
  OAI22_X1 U11 ( .A1(n37), .A2(n261), .B1(n258), .B2(n293), .ZN(n98) );
  INV_X1 U12 ( .A(DIN[1]), .ZN(n293) );
  OAI22_X1 U13 ( .A1(n38), .A2(n261), .B1(n258), .B2(n292), .ZN(n97) );
  INV_X1 U14 ( .A(DIN[2]), .ZN(n292) );
  OAI22_X1 U15 ( .A1(n39), .A2(n261), .B1(n258), .B2(n291), .ZN(n96) );
  INV_X1 U16 ( .A(DIN[3]), .ZN(n291) );
  OAI22_X1 U17 ( .A1(n40), .A2(n261), .B1(n258), .B2(n290), .ZN(n95) );
  INV_X1 U18 ( .A(DIN[4]), .ZN(n290) );
  OAI22_X1 U19 ( .A1(n41), .A2(n261), .B1(n258), .B2(n289), .ZN(n94) );
  INV_X1 U20 ( .A(DIN[5]), .ZN(n289) );
  OAI22_X1 U21 ( .A1(n42), .A2(n261), .B1(n258), .B2(n288), .ZN(n93) );
  INV_X1 U22 ( .A(DIN[6]), .ZN(n288) );
  OAI22_X1 U23 ( .A1(n43), .A2(n261), .B1(n258), .B2(n287), .ZN(n92) );
  INV_X1 U24 ( .A(DIN[7]), .ZN(n287) );
  OAI22_X1 U25 ( .A1(n44), .A2(n261), .B1(n258), .B2(n286), .ZN(n91) );
  INV_X1 U26 ( .A(DIN[8]), .ZN(n286) );
  OAI22_X1 U27 ( .A1(n45), .A2(n260), .B1(n258), .B2(n285), .ZN(n90) );
  INV_X1 U28 ( .A(DIN[9]), .ZN(n285) );
  OAI22_X1 U29 ( .A1(n65), .A2(n259), .B1(n256), .B2(n265), .ZN(n70) );
  INV_X1 U30 ( .A(DIN[29]), .ZN(n265) );
  OAI22_X1 U31 ( .A1(n61), .A2(n259), .B1(n256), .B2(n269), .ZN(n74) );
  INV_X1 U32 ( .A(DIN[25]), .ZN(n269) );
  OAI22_X1 U33 ( .A1(n67), .A2(n259), .B1(n256), .B2(n263), .ZN(n68) );
  INV_X1 U34 ( .A(DIN[31]), .ZN(n263) );
  OAI22_X1 U35 ( .A1(n59), .A2(n259), .B1(n256), .B2(n271), .ZN(n76) );
  INV_X1 U36 ( .A(DIN[23]), .ZN(n271) );
  OAI22_X1 U37 ( .A1(n64), .A2(n259), .B1(n256), .B2(n266), .ZN(n71) );
  INV_X1 U38 ( .A(DIN[28]), .ZN(n266) );
  OAI22_X1 U39 ( .A1(n58), .A2(n259), .B1(n256), .B2(n272), .ZN(n77) );
  INV_X1 U40 ( .A(DIN[22]), .ZN(n272) );
  OAI22_X1 U41 ( .A1(n60), .A2(n259), .B1(n256), .B2(n270), .ZN(n75) );
  INV_X1 U42 ( .A(DIN[24]), .ZN(n270) );
  OAI22_X1 U43 ( .A1(n57), .A2(n259), .B1(n256), .B2(n273), .ZN(n78) );
  INV_X1 U44 ( .A(DIN[21]), .ZN(n273) );
  OAI22_X1 U45 ( .A1(n46), .A2(n260), .B1(n257), .B2(n284), .ZN(n89) );
  INV_X1 U46 ( .A(DIN[10]), .ZN(n284) );
  OAI22_X1 U47 ( .A1(n47), .A2(n260), .B1(n257), .B2(n283), .ZN(n88) );
  INV_X1 U48 ( .A(DIN[11]), .ZN(n283) );
  OAI22_X1 U49 ( .A1(n48), .A2(n260), .B1(n257), .B2(n282), .ZN(n87) );
  INV_X1 U50 ( .A(DIN[12]), .ZN(n282) );
  OAI22_X1 U51 ( .A1(n49), .A2(n260), .B1(n257), .B2(n281), .ZN(n86) );
  INV_X1 U52 ( .A(DIN[13]), .ZN(n281) );
  OAI22_X1 U53 ( .A1(n50), .A2(n260), .B1(n257), .B2(n280), .ZN(n85) );
  INV_X1 U54 ( .A(DIN[14]), .ZN(n280) );
  OAI22_X1 U55 ( .A1(n51), .A2(n260), .B1(n257), .B2(n279), .ZN(n84) );
  INV_X1 U56 ( .A(DIN[15]), .ZN(n279) );
  OAI22_X1 U57 ( .A1(n52), .A2(n260), .B1(n257), .B2(n278), .ZN(n83) );
  INV_X1 U58 ( .A(DIN[16]), .ZN(n278) );
  OAI22_X1 U59 ( .A1(n53), .A2(n260), .B1(n257), .B2(n277), .ZN(n82) );
  INV_X1 U60 ( .A(DIN[17]), .ZN(n277) );
  OAI22_X1 U61 ( .A1(n54), .A2(n260), .B1(n257), .B2(n276), .ZN(n81) );
  INV_X1 U62 ( .A(DIN[18]), .ZN(n276) );
  OAI22_X1 U63 ( .A1(n55), .A2(n260), .B1(n257), .B2(n275), .ZN(n80) );
  INV_X1 U64 ( .A(DIN[19]), .ZN(n275) );
  OAI22_X1 U65 ( .A1(n56), .A2(n260), .B1(n257), .B2(n274), .ZN(n79) );
  INV_X1 U66 ( .A(DIN[20]), .ZN(n274) );
  OAI22_X1 U67 ( .A1(n62), .A2(n259), .B1(n256), .B2(n268), .ZN(n73) );
  INV_X1 U68 ( .A(DIN[26]), .ZN(n268) );
  OAI22_X1 U69 ( .A1(n63), .A2(n259), .B1(n256), .B2(n267), .ZN(n72) );
  INV_X1 U70 ( .A(DIN[27]), .ZN(n267) );
  OAI22_X1 U71 ( .A1(n66), .A2(n259), .B1(n256), .B2(n264), .ZN(n69) );
  INV_X1 U72 ( .A(DIN[30]), .ZN(n264) );
  NAND2_X1 U73 ( .A1(RST), .A2(n259), .ZN(n35) );
  NAND2_X1 U74 ( .A1(n262), .A2(RST), .ZN(n34) );
  INV_X1 U75 ( .A(EN), .ZN(n262) );
endmodule


module DLX_CU_WIDTH32_LENGTH5 ( CLK, RST, IR_IN, EN1, EN2, RF_RD1, RF_RD2, 
        MuxIMM_SEL, SIGN_EN, EN3, MuxA_SEL, MuxB_SEL, EQ_COND, JUMP_EN, RF_WE3, 
    .ALU_OPCODE({\ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , 
        \ALU_OPCODE[1] , \ALU_OPCODE[0] }), EN4, RF_WE4, DRAM_WE, SIGN_LD_EN, 
        MuxLD_SEL, MuxSW_SEL, MuxWB_SEL, RF_WE, JUMP_LINK );
  input [31:0] IR_IN;
  output [2:0] MuxLD_SEL;
  output [2:0] MuxSW_SEL;
  input CLK, RST;
  output EN1, EN2, RF_RD1, RF_RD2, MuxIMM_SEL, SIGN_EN, EN3, MuxA_SEL,
         MuxB_SEL, EQ_COND, JUMP_EN, RF_WE3, \ALU_OPCODE[4] , \ALU_OPCODE[3] ,
         \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] , EN4, RF_WE4,
         DRAM_WE, SIGN_LD_EN, MuxWB_SEL, RF_WE, JUMP_LINK;
  wire   IR_IN_31, IR_IN_30, IR_IN_29, IR_IN_28, IR_IN_27, IR_IN_26, RF_WE4,
         cw3_11, cw3_10, cw3_9, n47, n62, n142, n145, n138, n139, n140, n143,
         n43, n44, n45, n46, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n141, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406;
  wire   [4:0] ALU_OPCODE;
  wire   [21:0] cw1;
  wire   [16:0] cw2;
  wire   [7:0] cw3;
  wire   [2:0] cw4;
  wire   [4:0] aluOpcode1;
  wire   [4:0] aluOpcode2;
  wire   [21:0] cw;
  wire   [4:0] aluOpcodei;
  assign IR_IN_31 = IR_IN[31];
  assign IR_IN_30 = IR_IN[30];
  assign IR_IN_29 = IR_IN[29];
  assign IR_IN_28 = IR_IN[28];
  assign IR_IN_27 = IR_IN[27];
  assign IR_IN_26 = IR_IN[26];
  assign MuxLD_SEL[2] = RF_WE4;

  DFFR_X1 \cw1_reg[22]  ( .D(1'b1), .CK(CLK), .RN(n359), .Q(EN1) );
  DFFR_X1 \cw1_reg[21]  ( .D(cw[21]), .CK(CLK), .RN(n361), .Q(cw1[21]) );
  DFFR_X1 \cw1_reg[20]  ( .D(cw[20]), .CK(CLK), .RN(n359), .Q(cw1[20]) );
  SDFFR_X1 \cw1_reg[19]  ( .D(n371), .SI(1'b1), .SE(n141), .CK(CLK), .RN(n367), 
        .Q(cw1[19]) );
  DFFR_X1 \cw1_reg[18]  ( .D(cw[18]), .CK(CLK), .RN(n363), .Q(cw1[18]) );
  DFFR_X1 \cw1_reg[17]  ( .D(cw[17]), .CK(CLK), .RN(n359), .Q(cw1[17]) );
  DFFR_X1 \cw1_reg[16]  ( .D(cw[21]), .CK(CLK), .RN(n361), .Q(cw1[16]) );
  SDFFR_X1 \cw1_reg[15]  ( .D(n145), .SI(1'b1), .SE(n62), .CK(CLK), .RN(n367), 
        .Q(cw1[15]) );
  DFFR_X1 \cw1_reg[14]  ( .D(n371), .CK(CLK), .RN(n364), .Q(cw1[14]) );
  DFFR_X1 \cw1_reg[13]  ( .D(n138), .CK(CLK), .RN(n365), .Q(cw1[13]) );
  DFFR_X1 \cw1_reg[12]  ( .D(n372), .CK(CLK), .RN(n365), .Q(cw1[12]) );
  DFFR_X1 \cw1_reg[11]  ( .D(cw[21]), .CK(CLK), .RN(n362), .Q(cw1[11]) );
  DFFR_X1 \cw1_reg[10]  ( .D(n141), .CK(CLK), .RN(n363), .Q(cw1[10]) );
  SDFFR_X1 \cw1_reg[9]  ( .D(1'b0), .SI(n388), .SE(n47), .CK(CLK), .RN(n367), 
        .Q(cw1[9]) );
  DFFR_X1 \cw1_reg[8]  ( .D(n380), .CK(CLK), .RN(n366), .Q(cw1[8]) );
  DFFR_X1 \cw1_reg[7]  ( .D(n381), .CK(CLK), .RN(n366), .Q(cw1[7]) );
  DFFR_X1 \cw1_reg[6]  ( .D(cw[6]), .CK(CLK), .RN(n361), .Q(cw1[6]) );
  DFFR_X1 \cw1_reg[5]  ( .D(n139), .CK(CLK), .RN(n362), .Q(cw1[5]) );
  DFFR_X1 \cw1_reg[4]  ( .D(n140), .CK(CLK), .RN(n363), .Q(cw1[4]) );
  DFFR_X1 \cw1_reg[3]  ( .D(cw[3]), .CK(CLK), .RN(n360), .Q(cw1[3]) );
  DFFR_X1 \cw1_reg[2]  ( .D(n379), .CK(CLK), .RN(n366), .Q(cw1[2]) );
  DFFR_X1 \cw1_reg[1]  ( .D(n142), .CK(CLK), .RN(n360), .Q(cw1[1]) );
  DFFR_X1 \cw1_reg[0]  ( .D(n143), .CK(CLK), .RN(n363), .Q(cw1[0]) );
  DFFR_X1 \cw2_reg[21]  ( .D(cw1[21]), .CK(CLK), .RN(n361), .Q(EN2) );
  DFFR_X1 \cw2_reg[20]  ( .D(cw1[20]), .CK(CLK), .RN(n359), .Q(RF_RD1) );
  DFFR_X1 \cw2_reg[19]  ( .D(cw1[19]), .CK(CLK), .RN(n364), .Q(RF_RD2) );
  DFFR_X1 \cw2_reg[17]  ( .D(cw1[17]), .CK(CLK), .RN(n359), .Q(SIGN_EN) );
  DFFR_X1 \cw2_reg[16]  ( .D(cw1[16]), .CK(CLK), .RN(n361), .Q(cw2[16]) );
  DFFR_X1 \cw2_reg[15]  ( .D(cw1[15]), .CK(CLK), .RN(n365), .Q(cw2[15]) );
  DFFR_X1 \cw2_reg[14]  ( .D(cw1[14]), .CK(CLK), .RN(n364), .Q(cw2[14]) );
  DFFR_X1 \cw2_reg[13]  ( .D(cw1[13]), .CK(CLK), .RN(n365), .Q(cw2[13]) );
  DFFR_X1 \cw2_reg[12]  ( .D(cw1[12]), .CK(CLK), .RN(n364), .Q(cw2[12]) );
  DFFR_X1 \cw2_reg[11]  ( .D(cw1[11]), .CK(CLK), .RN(n361), .Q(cw2[11]) );
  DFFR_X1 \cw2_reg[10]  ( .D(cw1[10]), .CK(CLK), .RN(n363), .Q(cw2[10]) );
  DFFR_X1 \cw2_reg[9]  ( .D(cw1[9]), .CK(CLK), .RN(n364), .Q(cw2[9]) );
  DFFR_X1 \cw2_reg[8]  ( .D(cw1[8]), .CK(CLK), .RN(n366), .Q(cw2[8]) );
  DFFR_X1 \cw2_reg[7]  ( .D(cw1[7]), .CK(CLK), .RN(n367), .Q(cw2[7]) );
  DFFR_X1 \cw2_reg[6]  ( .D(cw1[6]), .CK(CLK), .RN(n361), .Q(cw2[6]) );
  DFFR_X1 \cw2_reg[5]  ( .D(cw1[5]), .CK(CLK), .RN(n362), .Q(cw2[5]) );
  DFFR_X1 \cw2_reg[4]  ( .D(cw1[4]), .CK(CLK), .RN(n363), .Q(cw2[4]) );
  DFFR_X1 \cw2_reg[3]  ( .D(cw1[3]), .CK(CLK), .RN(n360), .Q(cw2[3]) );
  DFFR_X1 \cw2_reg[2]  ( .D(cw1[2]), .CK(CLK), .RN(n366), .Q(cw2[2]) );
  DFFR_X1 \cw2_reg[1]  ( .D(cw1[1]), .CK(CLK), .RN(n360), .Q(cw2[1]) );
  DFFR_X1 \cw2_reg[0]  ( .D(cw1[0]), .CK(CLK), .RN(n363), .Q(cw2[0]) );
  DFFR_X1 \cw3_reg[16]  ( .D(cw2[16]), .CK(CLK), .RN(n361), .Q(EN3) );
  DFFR_X1 \cw3_reg[13]  ( .D(cw2[13]), .CK(CLK), .RN(n365), .Q(EQ_COND) );
  DFFR_X1 \cw3_reg[12]  ( .D(cw2[12]), .CK(CLK), .RN(n365), .Q(JUMP_EN) );
  DFFR_X1 \cw3_reg[11]  ( .D(cw2[11]), .CK(CLK), .RN(n360), .Q(cw3_11) );
  DFFR_X1 \cw3_reg[10]  ( .D(cw2[10]), .CK(CLK), .RN(n363), .Q(cw3_10) );
  DFFR_X1 \cw3_reg[9]  ( .D(cw2[9]), .CK(CLK), .RN(n364), .Q(cw3_9) );
  DFFR_X1 \cw3_reg[8]  ( .D(cw2[8]), .CK(CLK), .RN(n366), .Q(RF_WE3) );
  DFFR_X1 \cw3_reg[7]  ( .D(cw2[7]), .CK(CLK), .RN(n360), .Q(cw3[7]) );
  DFFR_X1 \cw3_reg[6]  ( .D(cw2[6]), .CK(CLK), .RN(n359), .Q(cw3[6]) );
  DFFR_X1 \cw3_reg[5]  ( .D(cw2[5]), .CK(CLK), .RN(n362), .Q(cw3[5]) );
  DFFR_X1 \cw3_reg[4]  ( .D(cw2[4]), .CK(CLK), .RN(n363), .Q(cw3[4]) );
  DFFR_X1 \cw3_reg[3]  ( .D(cw2[3]), .CK(CLK), .RN(n360), .Q(cw3[3]) );
  DFFR_X1 \cw3_reg[2]  ( .D(cw2[2]), .CK(CLK), .RN(n366), .Q(cw3[2]) );
  DFFR_X1 \cw3_reg[1]  ( .D(cw2[1]), .CK(CLK), .RN(n362), .Q(cw3[1]) );
  DFFR_X1 \cw3_reg[0]  ( .D(cw2[0]), .CK(CLK), .RN(n363), .Q(cw3[0]) );
  DFFR_X1 \cw4_reg[11]  ( .D(cw3_11), .CK(CLK), .RN(n360), .Q(EN4) );
  DFFR_X1 \cw4_reg[10]  ( .D(cw3_10), .CK(CLK), .RN(n363), .Q(DRAM_WE) );
  DFFR_X1 \cw4_reg[9]  ( .D(cw3_9), .CK(CLK), .RN(n364), .Q(SIGN_LD_EN) );
  DFFR_X1 \cw4_reg[8]  ( .D(RF_WE3), .CK(CLK), .RN(n365), .Q(RF_WE4) );
  DFFR_X1 \cw4_reg[7]  ( .D(cw3[7]), .CK(CLK), .RN(n360), .Q(MuxLD_SEL[1]) );
  DFFR_X1 \cw4_reg[6]  ( .D(cw3[6]), .CK(CLK), .RN(n360), .Q(MuxLD_SEL[0]) );
  DFFR_X1 \cw4_reg[5]  ( .D(cw3[5]), .CK(CLK), .RN(n362), .Q(MuxSW_SEL[2]) );
  DFFR_X1 \cw4_reg[4]  ( .D(cw3[4]), .CK(CLK), .RN(n364), .Q(MuxSW_SEL[1]) );
  DFFR_X1 \cw4_reg[3]  ( .D(cw3[3]), .CK(CLK), .RN(n359), .Q(MuxSW_SEL[0]) );
  DFFR_X1 \cw4_reg[2]  ( .D(cw3[2]), .CK(CLK), .RN(n366), .Q(cw4[2]) );
  DFFR_X1 \cw4_reg[1]  ( .D(cw3[1]), .CK(CLK), .RN(n361), .Q(cw4[1]) );
  DFFR_X1 \cw4_reg[0]  ( .D(cw3[0]), .CK(CLK), .RN(n365), .Q(cw4[0]) );
  DFFR_X1 \cw5_reg[1]  ( .D(cw4[1]), .CK(CLK), .RN(n361), .Q(RF_WE) );
  DFFR_X1 \aluOpcode1_reg[4]  ( .D(aluOpcodei[4]), .CK(CLK), .RN(n365), .Q(
        aluOpcode1[4]) );
  DFFR_X1 \aluOpcode1_reg[3]  ( .D(aluOpcodei[3]), .CK(CLK), .RN(n359), .Q(
        aluOpcode1[3]) );
  DFFR_X1 \aluOpcode1_reg[2]  ( .D(aluOpcodei[2]), .CK(CLK), .RN(n360), .Q(
        aluOpcode1[2]) );
  DFFR_X1 \aluOpcode1_reg[1]  ( .D(aluOpcodei[1]), .CK(CLK), .RN(n364), .Q(
        aluOpcode1[1]) );
  DFFR_X1 \aluOpcode1_reg[0]  ( .D(aluOpcodei[0]), .CK(CLK), .RN(n366), .Q(
        aluOpcode1[0]) );
  DFFR_X1 \aluOpcode2_reg[4]  ( .D(aluOpcode1[4]), .CK(CLK), .RN(n365), .Q(
        aluOpcode2[4]) );
  DFFR_X1 \aluOpcode3_reg[4]  ( .D(aluOpcode2[4]), .CK(CLK), .RN(n365), .Q(
        ALU_OPCODE[4]) );
  DFFR_X1 \aluOpcode2_reg[3]  ( .D(aluOpcode1[3]), .CK(CLK), .RN(n359), .Q(
        aluOpcode2[3]) );
  DFFR_X1 \aluOpcode3_reg[3]  ( .D(aluOpcode2[3]), .CK(CLK), .RN(n362), .Q(
        ALU_OPCODE[3]) );
  DFFR_X1 \aluOpcode2_reg[2]  ( .D(aluOpcode1[2]), .CK(CLK), .RN(n359), .Q(
        aluOpcode2[2]) );
  DFFR_X1 \aluOpcode3_reg[2]  ( .D(aluOpcode2[2]), .CK(CLK), .RN(n359), .Q(
        ALU_OPCODE[2]) );
  DFFR_X1 \aluOpcode2_reg[1]  ( .D(aluOpcode1[1]), .CK(CLK), .RN(n364), .Q(
        aluOpcode2[1]) );
  DFFR_X1 \aluOpcode3_reg[1]  ( .D(aluOpcode2[1]), .CK(CLK), .RN(n364), .Q(
        ALU_OPCODE[1]) );
  DFFR_X1 \aluOpcode2_reg[0]  ( .D(aluOpcode1[0]), .CK(CLK), .RN(n366), .Q(
        aluOpcode2[0]) );
  DFFR_X1 \aluOpcode3_reg[0]  ( .D(aluOpcode2[0]), .CK(CLK), .RN(n366), .Q(
        ALU_OPCODE[0]) );
  DFFR_X1 \cw3_reg[14]  ( .D(cw2[14]), .CK(CLK), .RN(n362), .Q(MuxB_SEL) );
  DFFR_X1 \cw3_reg[15]  ( .D(cw2[15]), .CK(CLK), .RN(n362), .Q(MuxA_SEL) );
  DFFR_X1 \cw2_reg[18]  ( .D(cw1[18]), .CK(CLK), .RN(n361), .Q(MuxIMM_SEL) );
  DFFR_X1 \cw5_reg[2]  ( .D(cw4[2]), .CK(CLK), .RN(n362), .Q(MuxWB_SEL) );
  DFFR_X1 \cw5_reg[0]  ( .D(cw4[0]), .CK(CLK), .RN(n362), .Q(JUMP_LINK) );
  NAND3_X1 U141 ( .A1(n49), .A2(n50), .A3(n51), .ZN(cw[6]) );
  NAND3_X1 U142 ( .A1(n48), .A2(n53), .A3(n49), .ZN(cw[21]) );
  NAND3_X1 U143 ( .A1(n68), .A2(n69), .A3(IR_IN[5]), .ZN(n67) );
  NAND3_X1 U144 ( .A1(n368), .A2(IR_IN[0]), .A3(n89), .ZN(n85) );
  NAND3_X1 U145 ( .A1(n105), .A2(n106), .A3(n107), .ZN(n104) );
  NAND3_X1 U146 ( .A1(n394), .A2(n71), .A3(n61), .ZN(n107) );
  NAND3_X1 U147 ( .A1(IR_IN_29), .A2(IR_IN_31), .A3(n120), .ZN(n119) );
  NAND3_X1 U148 ( .A1(n368), .A2(n398), .A3(n122), .ZN(n106) );
  NAND3_X1 U149 ( .A1(n133), .A2(n402), .A3(IR_IN_29), .ZN(n45) );
  NAND3_X1 U150 ( .A1(n44), .A2(n43), .A3(n50), .ZN(n56) );
  NAND3_X1 U151 ( .A1(n133), .A2(n406), .A3(n46), .ZN(n43) );
  NAND3_X1 U152 ( .A1(n103), .A2(n406), .A3(n133), .ZN(n44) );
  NAND3_X1 U153 ( .A1(n108), .A2(n131), .A3(n120), .ZN(n55) );
  NAND3_X1 U154 ( .A1(n95), .A2(n131), .A3(n120), .ZN(n72) );
  NAND3_X1 U155 ( .A1(n393), .A2(n401), .A3(n61), .ZN(n98) );
  NAND3_X1 U156 ( .A1(n136), .A2(n397), .A3(n368), .ZN(n126) );
  NAND3_X1 U157 ( .A1(n402), .A2(n378), .A3(n131), .ZN(n134) );
  OR3_X1 U3 ( .A1(n56), .A2(n143), .A3(n370), .ZN(n142) );
  INV_X1 U7 ( .A(n49), .ZN(n370) );
  INV_X1 U8 ( .A(n57), .ZN(n384) );
  INV_X1 U9 ( .A(n53), .ZN(n372) );
  INV_X1 U10 ( .A(n48), .ZN(n379) );
  NOR3_X1 U11 ( .A1(n57), .A2(n371), .A3(n58), .ZN(n49) );
  INV_X1 U12 ( .A(n132), .ZN(n390) );
  NOR2_X1 U13 ( .A1(n389), .A2(n134), .ZN(n61) );
  NOR3_X1 U14 ( .A1(n143), .A2(n62), .A3(n377), .ZN(n53) );
  NOR2_X1 U15 ( .A1(n56), .A2(n141), .ZN(n48) );
  NOR2_X1 U16 ( .A1(n385), .A2(n387), .ZN(n57) );
  INV_X1 U17 ( .A(n95), .ZN(n387) );
  OAI21_X1 U18 ( .B1(n80), .B2(n81), .A(n106), .ZN(n96) );
  AOI21_X1 U19 ( .B1(n382), .B2(n81), .A(n387), .ZN(n115) );
  NAND2_X1 U20 ( .A1(n90), .A2(n390), .ZN(n75) );
  NOR2_X1 U21 ( .A1(n387), .A2(n134), .ZN(n145) );
  INV_X1 U22 ( .A(n52), .ZN(n375) );
  INV_X1 U23 ( .A(n97), .ZN(n368) );
  NAND2_X1 U24 ( .A1(n373), .A2(n72), .ZN(n143) );
  INV_X1 U25 ( .A(n145), .ZN(n373) );
  NOR3_X1 U26 ( .A1(n52), .A2(n372), .A3(n141), .ZN(n51) );
  INV_X1 U27 ( .A(n55), .ZN(n377) );
  INV_X1 U28 ( .A(n66), .ZN(n394) );
  INV_X1 U29 ( .A(n81), .ZN(n376) );
  INV_X1 U30 ( .A(n65), .ZN(n393) );
  AND2_X1 U31 ( .A1(n77), .A2(n387), .ZN(n80) );
  NAND2_X1 U32 ( .A1(n47), .A2(n95), .ZN(n50) );
  INV_X1 U33 ( .A(n44), .ZN(n380) );
  INV_X1 U34 ( .A(n43), .ZN(n381) );
  NAND2_X1 U35 ( .A1(n60), .A2(n384), .ZN(cw[18]) );
  OAI21_X1 U36 ( .B1(n386), .B2(n385), .A(n91), .ZN(n84) );
  NOR2_X1 U37 ( .A1(n103), .A2(n46), .ZN(n132) );
  NAND4_X1 U38 ( .A1(n374), .A2(n75), .A3(n382), .A4(n76), .ZN(n58) );
  INV_X1 U39 ( .A(n83), .ZN(n385) );
  INV_X1 U40 ( .A(n109), .ZN(n405) );
  OR4_X1 U41 ( .A1(n142), .A2(n62), .A3(n52), .A4(n54), .ZN(cw[3]) );
  OAI21_X1 U42 ( .B1(n387), .B2(n45), .A(n55), .ZN(n54) );
  INV_X1 U43 ( .A(n79), .ZN(n374) );
  OAI211_X1 U44 ( .C1(n80), .C2(n375), .A(n81), .B(n82), .ZN(n79) );
  AOI21_X1 U45 ( .B1(n83), .B2(n390), .A(n84), .ZN(n82) );
  NOR4_X1 U46 ( .A1(n378), .A2(n402), .A3(n406), .A4(n403), .ZN(n90) );
  NOR3_X1 U47 ( .A1(n402), .A2(n404), .A3(n378), .ZN(n52) );
  OAI222_X1 U48 ( .A1(n386), .A2(n375), .B1(n88), .B2(n399), .C1(n77), .C2(
        n385), .ZN(n129) );
  NAND4_X1 U49 ( .A1(n369), .A2(n383), .A3(n100), .A4(n101), .ZN(aluOpcodei[2]) );
  AOI22_X1 U50 ( .A1(n376), .A2(n108), .B1(n83), .B2(n46), .ZN(n100) );
  INV_X1 U51 ( .A(n84), .ZN(n383) );
  AOI221_X1 U52 ( .B1(n102), .B2(n368), .C1(n90), .C2(n103), .A(n104), .ZN(
        n101) );
  AOI21_X1 U53 ( .B1(n387), .B2(n132), .A(n45), .ZN(n141) );
  NOR2_X1 U54 ( .A1(n392), .A2(n388), .ZN(n95) );
  NOR2_X1 U55 ( .A1(n108), .A2(n103), .ZN(n77) );
  OAI21_X1 U56 ( .B1(n134), .B2(n386), .A(n73), .ZN(n62) );
  NOR2_X1 U57 ( .A1(n398), .A2(n400), .ZN(n71) );
  NOR3_X1 U58 ( .A1(n405), .A2(n389), .A3(n402), .ZN(n114) );
  NAND4_X1 U59 ( .A1(n68), .A2(n401), .A3(n397), .A4(n396), .ZN(n66) );
  NOR3_X1 U60 ( .A1(n396), .A2(n116), .A3(n88), .ZN(n113) );
  AOI21_X1 U61 ( .B1(n99), .B2(n401), .A(n102), .ZN(n116) );
  NAND2_X1 U62 ( .A1(n109), .A2(n120), .ZN(n81) );
  NAND4_X1 U63 ( .A1(n71), .A2(n68), .A3(n396), .A4(n395), .ZN(n65) );
  INV_X1 U64 ( .A(n103), .ZN(n389) );
  INV_X1 U65 ( .A(n108), .ZN(n386) );
  INV_X1 U66 ( .A(n121), .ZN(n382) );
  OAI211_X1 U67 ( .C1(n77), .C2(n382), .A(n374), .B(n78), .ZN(cw[17]) );
  AND3_X1 U68 ( .A1(n384), .A2(n48), .A3(n73), .ZN(n78) );
  NOR2_X1 U69 ( .A1(n70), .A2(n88), .ZN(n87) );
  NOR2_X1 U70 ( .A1(n391), .A2(n45), .ZN(n140) );
  INV_X1 U71 ( .A(n46), .ZN(n391) );
  NOR2_X1 U72 ( .A1(n389), .A2(n45), .ZN(n139) );
  NAND4_X1 U73 ( .A1(n369), .A2(n110), .A3(n111), .A4(n112), .ZN(aluOpcodei[1]) );
  NAND2_X1 U74 ( .A1(n90), .A2(n46), .ZN(n110) );
  AOI21_X1 U75 ( .B1(n368), .B2(n117), .A(n118), .ZN(n111) );
  NOR4_X1 U76 ( .A1(n57), .A2(n113), .A3(n114), .A4(n115), .ZN(n112) );
  NAND4_X1 U77 ( .A1(n126), .A2(n76), .A3(n127), .A4(n128), .ZN(aluOpcodei[0])
         );
  AND3_X1 U78 ( .A1(n98), .A2(n53), .A3(n48), .ZN(n127) );
  AOI211_X1 U79 ( .C1(n121), .C2(n390), .A(n129), .B(n96), .ZN(n128) );
  NAND2_X1 U80 ( .A1(n130), .A2(n396), .ZN(n97) );
  INV_X1 U81 ( .A(n99), .ZN(n399) );
  INV_X1 U82 ( .A(n131), .ZN(n404) );
  AND3_X1 U83 ( .A1(n402), .A2(n406), .A3(n133), .ZN(n47) );
  INV_X1 U84 ( .A(n59), .ZN(n371) );
  AND4_X1 U85 ( .A1(n72), .A2(n48), .A3(n73), .A4(n74), .ZN(n60) );
  NOR2_X1 U86 ( .A1(n377), .A2(n58), .ZN(n74) );
  NAND2_X1 U87 ( .A1(n60), .A2(n59), .ZN(cw[20]) );
  NOR2_X1 U88 ( .A1(n392), .A2(IR_IN_27), .ZN(n46) );
  NOR3_X1 U89 ( .A1(n402), .A2(IR_IN_30), .A3(n405), .ZN(n83) );
  NOR2_X1 U90 ( .A1(IR_IN_26), .A2(IR_IN_27), .ZN(n103) );
  INV_X1 U91 ( .A(IR_IN_28), .ZN(n402) );
  NOR2_X1 U92 ( .A1(n406), .A2(IR_IN_31), .ZN(n109) );
  NAND4_X1 U93 ( .A1(n109), .A2(IR_IN_30), .A3(IR_IN_28), .A4(n390), .ZN(n91)
         );
  INV_X1 U94 ( .A(IR_IN_29), .ZN(n406) );
  INV_X1 U95 ( .A(IR_IN_26), .ZN(n392) );
  NOR3_X1 U96 ( .A1(IR_IN[6]), .A2(IR_IN[10]), .A3(n137), .ZN(n68) );
  OR3_X1 U97 ( .A1(IR_IN[9]), .A2(IR_IN[8]), .A3(IR_IN[7]), .ZN(n137) );
  NOR3_X1 U98 ( .A1(IR_IN_28), .A2(IR_IN_30), .A3(n405), .ZN(n121) );
  NOR3_X1 U99 ( .A1(n398), .A2(IR_IN[1]), .A3(n401), .ZN(n102) );
  NOR2_X1 U100 ( .A1(IR_IN_29), .A2(IR_IN_31), .ZN(n131) );
  NOR2_X1 U101 ( .A1(n378), .A2(IR_IN_28), .ZN(n120) );
  AOI21_X1 U102 ( .B1(n400), .B2(IR_IN[2]), .A(n99), .ZN(n70) );
  NOR2_X1 U103 ( .A1(n388), .A2(IR_IN_26), .ZN(n108) );
  NAND2_X1 U104 ( .A1(n61), .A2(n63), .ZN(n59) );
  OAI221_X1 U105 ( .B1(n64), .B2(n65), .C1(n398), .C2(n66), .A(n67), .ZN(n63)
         );
  NOR2_X1 U106 ( .A1(n397), .A2(n401), .ZN(n64) );
  NAND4_X1 U107 ( .A1(IR_IN_28), .A2(n131), .A3(n390), .A4(n378), .ZN(n73) );
  NOR4_X1 U108 ( .A1(IR_IN_30), .A2(n404), .A3(n389), .A4(n402), .ZN(n138) );
  NOR2_X1 U109 ( .A1(n400), .A2(IR_IN[2]), .ZN(n99) );
  INV_X1 U110 ( .A(IR_IN[3]), .ZN(n397) );
  NAND4_X1 U111 ( .A1(n120), .A2(IR_IN_29), .A3(IR_IN_31), .A4(n135), .ZN(n76)
         );
  NAND2_X1 U112 ( .A1(n387), .A2(n386), .ZN(n135) );
  INV_X1 U113 ( .A(IR_IN[2]), .ZN(n398) );
  INV_X1 U114 ( .A(IR_IN[0]), .ZN(n401) );
  NOR2_X1 U115 ( .A1(n403), .A2(IR_IN_30), .ZN(n133) );
  OAI22_X1 U116 ( .A1(IR_IN[2]), .A2(IR_IN[1]), .B1(IR_IN[0]), .B2(n398), .ZN(
        n136) );
  OAI22_X1 U117 ( .A1(n70), .A2(n397), .B1(IR_IN[4]), .B2(n71), .ZN(n69) );
  INV_X1 U118 ( .A(IR_IN_30), .ZN(n378) );
  NAND2_X1 U119 ( .A1(n130), .A2(IR_IN[3]), .ZN(n88) );
  AOI21_X1 U120 ( .B1(n382), .B2(n119), .A(n386), .ZN(n118) );
  NOR2_X1 U121 ( .A1(n397), .A2(IR_IN[0]), .ZN(n122) );
  INV_X1 U122 ( .A(IR_IN[1]), .ZN(n400) );
  INV_X1 U123 ( .A(IR_IN[4]), .ZN(n396) );
  OAI21_X1 U124 ( .B1(n122), .B2(n399), .A(n123), .ZN(n117) );
  OAI211_X1 U125 ( .C1(IR_IN[2]), .C2(IR_IN[3]), .A(n401), .B(n400), .ZN(n123)
         );
  INV_X1 U126 ( .A(IR_IN_31), .ZN(n403) );
  OR4_X1 U127 ( .A1(n88), .A2(n398), .A3(IR_IN[0]), .A4(IR_IN[1]), .ZN(n105)
         );
  INV_X1 U128 ( .A(IR_IN_27), .ZN(n388) );
  NAND4_X1 U129 ( .A1(n75), .A2(n76), .A3(n85), .A4(n86), .ZN(aluOpcodei[4])
         );
  AOI22_X1 U130 ( .A1(n87), .A2(IR_IN[4]), .B1(n376), .B2(n46), .ZN(n86) );
  NOR3_X1 U131 ( .A1(n397), .A2(IR_IN[2]), .A3(IR_IN[1]), .ZN(n89) );
  NAND4_X1 U132 ( .A1(n384), .A2(n91), .A3(n92), .A4(n93), .ZN(aluOpcodei[3])
         );
  NAND4_X1 U133 ( .A1(n61), .A2(n393), .A3(IR_IN[0]), .A4(n397), .ZN(n92) );
  AOI221_X1 U134 ( .B1(IR_IN[3]), .B2(n94), .C1(n52), .C2(n95), .A(n96), .ZN(
        n93) );
  OAI21_X1 U135 ( .B1(n70), .B2(n97), .A(n98), .ZN(n94) );
  AND3_X1 U136 ( .A1(IR_IN[5]), .A2(n68), .A3(n61), .ZN(n130) );
  INV_X1 U137 ( .A(IR_IN[5]), .ZN(n395) );
  INV_X1 U138 ( .A(n124), .ZN(n369) );
  OAI221_X1 U139 ( .B1(n389), .B2(n81), .C1(n77), .C2(n375), .A(n125), .ZN(
        n124) );
  NAND4_X1 U140 ( .A1(n61), .A2(n394), .A3(IR_IN[2]), .A4(n395), .ZN(n125) );
  CLKBUF_X1 U158 ( .A(RST), .Z(n356) );
  CLKBUF_X1 U159 ( .A(RST), .Z(n357) );
  CLKBUF_X1 U160 ( .A(RST), .Z(n358) );
  CLKBUF_X1 U161 ( .A(n356), .Z(n359) );
  CLKBUF_X1 U162 ( .A(n356), .Z(n360) );
  CLKBUF_X1 U163 ( .A(n356), .Z(n361) );
  CLKBUF_X1 U164 ( .A(n357), .Z(n362) );
  CLKBUF_X1 U165 ( .A(n357), .Z(n363) );
  CLKBUF_X1 U166 ( .A(n357), .Z(n364) );
  CLKBUF_X1 U167 ( .A(n358), .Z(n365) );
  CLKBUF_X1 U168 ( .A(n358), .Z(n366) );
  CLKBUF_X1 U169 ( .A(n358), .Z(n367) );
endmodule


module REGISTER_GENERIC_WIDTH32_11 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294;

  DFF_X1 \DOUT_reg[30]  ( .D(n69), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[29]  ( .D(n70), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[28]  ( .D(n71), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[27]  ( .D(n72), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n73), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[25]  ( .D(n74), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[24]  ( .D(n75), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[22]  ( .D(n77), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[21]  ( .D(n78), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[20]  ( .D(n79), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n80), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n81), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n83), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n84), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n89), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n90), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n91), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n92), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n93), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n94), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n95), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n96), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n97), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n98), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  DFF_X1 \DOUT_reg[31]  ( .D(n68), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  BUF_X1 U3 ( .A(n35), .Z(n258) );
  BUF_X1 U4 ( .A(n35), .Z(n257) );
  BUF_X1 U5 ( .A(n35), .Z(n256) );
  BUF_X1 U6 ( .A(n34), .Z(n261) );
  NAND2_X1 U7 ( .A1(RST), .A2(n259), .ZN(n35) );
  BUF_X1 U8 ( .A(n34), .Z(n259) );
  BUF_X1 U9 ( .A(n34), .Z(n260) );
  OAI22_X1 U10 ( .A1(n55), .A2(n260), .B1(n257), .B2(n280), .ZN(n80) );
  INV_X1 U11 ( .A(DIN[19]), .ZN(n280) );
  OAI22_X1 U12 ( .A1(n59), .A2(n259), .B1(n256), .B2(n278), .ZN(n76) );
  INV_X1 U13 ( .A(DIN[23]), .ZN(n278) );
  OAI22_X1 U14 ( .A1(n63), .A2(n259), .B1(n256), .B2(n276), .ZN(n72) );
  INV_X1 U15 ( .A(DIN[27]), .ZN(n276) );
  OAI22_X1 U16 ( .A1(n67), .A2(n259), .B1(n256), .B2(n275), .ZN(n68) );
  INV_X1 U17 ( .A(DIN[31]), .ZN(n275) );
  OAI22_X1 U18 ( .A1(n56), .A2(n260), .B1(n257), .B2(n269), .ZN(n79) );
  INV_X1 U19 ( .A(DIN[20]), .ZN(n269) );
  OAI22_X1 U20 ( .A1(n60), .A2(n259), .B1(n256), .B2(n271), .ZN(n75) );
  INV_X1 U21 ( .A(DIN[24]), .ZN(n271) );
  OAI22_X1 U22 ( .A1(n64), .A2(n259), .B1(n256), .B2(n273), .ZN(n71) );
  INV_X1 U23 ( .A(DIN[28]), .ZN(n273) );
  OAI22_X1 U24 ( .A1(n66), .A2(n259), .B1(n256), .B2(n274), .ZN(n69) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n274) );
  OAI22_X1 U26 ( .A1(n58), .A2(n259), .B1(n256), .B2(n279), .ZN(n77) );
  INV_X1 U27 ( .A(DIN[22]), .ZN(n279) );
  OAI22_X1 U28 ( .A1(n57), .A2(n259), .B1(n256), .B2(n268), .ZN(n78) );
  INV_X1 U29 ( .A(DIN[21]), .ZN(n268) );
  OAI22_X1 U30 ( .A1(n61), .A2(n259), .B1(n256), .B2(n270), .ZN(n74) );
  INV_X1 U31 ( .A(DIN[25]), .ZN(n270) );
  OAI22_X1 U32 ( .A1(n65), .A2(n259), .B1(n256), .B2(n272), .ZN(n70) );
  INV_X1 U33 ( .A(DIN[29]), .ZN(n272) );
  OAI22_X1 U34 ( .A1(n62), .A2(n259), .B1(n256), .B2(n277), .ZN(n73) );
  INV_X1 U35 ( .A(DIN[26]), .ZN(n277) );
  OAI22_X1 U36 ( .A1(n54), .A2(n260), .B1(n257), .B2(n281), .ZN(n81) );
  INV_X1 U37 ( .A(DIN[18]), .ZN(n281) );
  NAND2_X1 U38 ( .A1(n262), .A2(RST), .ZN(n34) );
  INV_X1 U39 ( .A(EN), .ZN(n262) );
  OAI22_X1 U40 ( .A1(n36), .A2(n261), .B1(n258), .B2(n292), .ZN(n99) );
  INV_X1 U41 ( .A(DIN[0]), .ZN(n292) );
  OAI22_X1 U42 ( .A1(n37), .A2(n261), .B1(n258), .B2(n294), .ZN(n98) );
  INV_X1 U43 ( .A(DIN[1]), .ZN(n294) );
  OAI22_X1 U44 ( .A1(n38), .A2(n261), .B1(n258), .B2(n293), .ZN(n97) );
  INV_X1 U45 ( .A(DIN[2]), .ZN(n293) );
  OAI22_X1 U46 ( .A1(n39), .A2(n261), .B1(n258), .B2(n291), .ZN(n96) );
  INV_X1 U47 ( .A(DIN[3]), .ZN(n291) );
  OAI22_X1 U48 ( .A1(n40), .A2(n261), .B1(n258), .B2(n289), .ZN(n95) );
  INV_X1 U49 ( .A(DIN[4]), .ZN(n289) );
  OAI22_X1 U50 ( .A1(n41), .A2(n261), .B1(n258), .B2(n290), .ZN(n94) );
  INV_X1 U51 ( .A(DIN[5]), .ZN(n290) );
  OAI22_X1 U52 ( .A1(n42), .A2(n261), .B1(n258), .B2(n288), .ZN(n93) );
  INV_X1 U53 ( .A(DIN[6]), .ZN(n288) );
  OAI22_X1 U54 ( .A1(n43), .A2(n261), .B1(n258), .B2(n263), .ZN(n92) );
  INV_X1 U55 ( .A(DIN[7]), .ZN(n263) );
  OAI22_X1 U56 ( .A1(n44), .A2(n261), .B1(n258), .B2(n287), .ZN(n91) );
  INV_X1 U57 ( .A(DIN[8]), .ZN(n287) );
  OAI22_X1 U58 ( .A1(n45), .A2(n260), .B1(n258), .B2(n286), .ZN(n90) );
  INV_X1 U59 ( .A(DIN[9]), .ZN(n286) );
  OAI22_X1 U60 ( .A1(n47), .A2(n260), .B1(n257), .B2(n285), .ZN(n88) );
  INV_X1 U61 ( .A(DIN[11]), .ZN(n285) );
  OAI22_X1 U62 ( .A1(n51), .A2(n260), .B1(n257), .B2(n282), .ZN(n84) );
  INV_X1 U63 ( .A(DIN[15]), .ZN(n282) );
  OAI22_X1 U64 ( .A1(n53), .A2(n260), .B1(n257), .B2(n266), .ZN(n82) );
  INV_X1 U65 ( .A(DIN[17]), .ZN(n266) );
  OAI22_X1 U66 ( .A1(n48), .A2(n260), .B1(n257), .B2(n265), .ZN(n87) );
  INV_X1 U67 ( .A(DIN[12]), .ZN(n265) );
  OAI22_X1 U68 ( .A1(n52), .A2(n260), .B1(n257), .B2(n267), .ZN(n83) );
  INV_X1 U69 ( .A(DIN[16]), .ZN(n267) );
  OAI22_X1 U70 ( .A1(n50), .A2(n260), .B1(n257), .B2(n283), .ZN(n85) );
  INV_X1 U71 ( .A(DIN[14]), .ZN(n283) );
  OAI22_X1 U72 ( .A1(n46), .A2(n260), .B1(n257), .B2(n284), .ZN(n89) );
  INV_X1 U73 ( .A(DIN[10]), .ZN(n284) );
  OAI22_X1 U74 ( .A1(n49), .A2(n260), .B1(n257), .B2(n264), .ZN(n86) );
  INV_X1 U75 ( .A(DIN[13]), .ZN(n264) );
endmodule


module MUX21_GENERIC_NBIT32_0 ( S1, S0, SEL, Y );
  input [31:0] S1;
  input [31:0] S0;
  output [31:0] Y;
  input SEL;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250;

  INV_X1 U1 ( .A(n250), .ZN(n240) );
  INV_X1 U2 ( .A(n250), .ZN(n241) );
  INV_X1 U3 ( .A(n51), .ZN(Y[14]) );
  AOI22_X1 U4 ( .A1(S0[14]), .A2(n241), .B1(S1[14]), .B2(n245), .ZN(n51) );
  INV_X1 U5 ( .A(n38), .ZN(Y[27]) );
  AOI22_X1 U6 ( .A1(S0[27]), .A2(n240), .B1(S1[27]), .B2(n242), .ZN(n38) );
  INV_X1 U7 ( .A(n37), .ZN(Y[28]) );
  AOI22_X1 U8 ( .A1(S0[28]), .A2(n241), .B1(S1[28]), .B2(n242), .ZN(n37) );
  INV_X1 U9 ( .A(n34), .ZN(Y[31]) );
  AOI22_X1 U10 ( .A1(S0[31]), .A2(n241), .B1(n249), .B2(S1[31]), .ZN(n34) );
  INV_X1 U11 ( .A(n52), .ZN(Y[13]) );
  AOI22_X1 U12 ( .A1(S0[13]), .A2(n241), .B1(S1[13]), .B2(n246), .ZN(n52) );
  INV_X1 U13 ( .A(n50), .ZN(Y[15]) );
  AOI22_X1 U14 ( .A1(S0[15]), .A2(n241), .B1(S1[15]), .B2(n245), .ZN(n50) );
  BUF_X1 U15 ( .A(n239), .Z(n248) );
  BUF_X1 U16 ( .A(n238), .Z(n247) );
  BUF_X1 U17 ( .A(n238), .Z(n245) );
  BUF_X1 U18 ( .A(n237), .Z(n244) );
  BUF_X1 U19 ( .A(n238), .Z(n246) );
  BUF_X1 U20 ( .A(n237), .Z(n243) );
  BUF_X1 U21 ( .A(n237), .Z(n242) );
  BUF_X1 U22 ( .A(n239), .Z(n250) );
  BUF_X1 U23 ( .A(n239), .Z(n249) );
  INV_X1 U24 ( .A(n61), .ZN(Y[4]) );
  AOI22_X1 U25 ( .A1(S0[4]), .A2(n240), .B1(S1[4]), .B2(n248), .ZN(n61) );
  INV_X1 U26 ( .A(n60), .ZN(Y[5]) );
  AOI22_X1 U27 ( .A1(S0[5]), .A2(n240), .B1(S1[5]), .B2(n248), .ZN(n60) );
  INV_X1 U28 ( .A(n59), .ZN(Y[6]) );
  AOI22_X1 U29 ( .A1(S0[6]), .A2(n240), .B1(S1[6]), .B2(n248), .ZN(n59) );
  INV_X1 U30 ( .A(n58), .ZN(Y[7]) );
  AOI22_X1 U31 ( .A1(S0[7]), .A2(n240), .B1(S1[7]), .B2(n247), .ZN(n58) );
  INV_X1 U32 ( .A(n57), .ZN(Y[8]) );
  AOI22_X1 U33 ( .A1(S0[8]), .A2(n240), .B1(S1[8]), .B2(n247), .ZN(n57) );
  INV_X1 U34 ( .A(n54), .ZN(Y[11]) );
  AOI22_X1 U35 ( .A1(S0[11]), .A2(n240), .B1(S1[11]), .B2(n246), .ZN(n54) );
  INV_X1 U36 ( .A(n53), .ZN(Y[12]) );
  AOI22_X1 U37 ( .A1(S0[12]), .A2(n241), .B1(S1[12]), .B2(n246), .ZN(n53) );
  INV_X1 U38 ( .A(n49), .ZN(Y[16]) );
  AOI22_X1 U39 ( .A1(S0[16]), .A2(n241), .B1(S1[16]), .B2(n245), .ZN(n49) );
  INV_X1 U40 ( .A(n47), .ZN(Y[18]) );
  AOI22_X1 U41 ( .A1(S0[18]), .A2(n241), .B1(S1[18]), .B2(n244), .ZN(n47) );
  INV_X1 U42 ( .A(n46), .ZN(Y[19]) );
  AOI22_X1 U43 ( .A1(S0[19]), .A2(n241), .B1(S1[19]), .B2(n244), .ZN(n46) );
  INV_X1 U44 ( .A(n44), .ZN(Y[21]) );
  AOI22_X1 U45 ( .A1(S0[21]), .A2(n241), .B1(S1[21]), .B2(n244), .ZN(n44) );
  INV_X1 U46 ( .A(n43), .ZN(Y[22]) );
  AOI22_X1 U47 ( .A1(S0[22]), .A2(n241), .B1(S1[22]), .B2(n243), .ZN(n43) );
  INV_X1 U48 ( .A(n63), .ZN(Y[2]) );
  AOI22_X1 U49 ( .A1(S0[2]), .A2(n240), .B1(S1[2]), .B2(n249), .ZN(n63) );
  INV_X1 U50 ( .A(n40), .ZN(Y[25]) );
  AOI22_X1 U51 ( .A1(S0[25]), .A2(n240), .B1(S1[25]), .B2(n243), .ZN(n40) );
  INV_X1 U52 ( .A(n39), .ZN(Y[26]) );
  AOI22_X1 U53 ( .A1(S0[26]), .A2(n241), .B1(S1[26]), .B2(n243), .ZN(n39) );
  INV_X1 U54 ( .A(n36), .ZN(Y[29]) );
  AOI22_X1 U55 ( .A1(S0[29]), .A2(n240), .B1(S1[29]), .B2(n242), .ZN(n36) );
  INV_X1 U56 ( .A(n35), .ZN(Y[30]) );
  AOI22_X1 U57 ( .A1(S0[30]), .A2(n241), .B1(S1[30]), .B2(n242), .ZN(n35) );
  INV_X1 U58 ( .A(n42), .ZN(Y[23]) );
  AOI22_X1 U59 ( .A1(S0[23]), .A2(n241), .B1(S1[23]), .B2(n246), .ZN(n42) );
  INV_X1 U60 ( .A(n41), .ZN(Y[24]) );
  AOI22_X1 U61 ( .A1(S0[24]), .A2(n240), .B1(S1[24]), .B2(n243), .ZN(n41) );
  BUF_X1 U62 ( .A(SEL), .Z(n239) );
  BUF_X1 U63 ( .A(SEL), .Z(n238) );
  BUF_X1 U64 ( .A(SEL), .Z(n237) );
  INV_X1 U65 ( .A(n62), .ZN(Y[3]) );
  AOI22_X1 U66 ( .A1(S0[3]), .A2(n240), .B1(S1[3]), .B2(n248), .ZN(n62) );
  INV_X1 U67 ( .A(n56), .ZN(Y[9]) );
  AOI22_X1 U68 ( .A1(S0[9]), .A2(n240), .B1(S1[9]), .B2(n247), .ZN(n56) );
  INV_X1 U69 ( .A(n55), .ZN(Y[10]) );
  AOI22_X1 U70 ( .A1(S0[10]), .A2(n240), .B1(S1[10]), .B2(n247), .ZN(n55) );
  INV_X1 U71 ( .A(n48), .ZN(Y[17]) );
  AOI22_X1 U72 ( .A1(S0[17]), .A2(n241), .B1(S1[17]), .B2(n245), .ZN(n48) );
  INV_X1 U73 ( .A(n45), .ZN(Y[20]) );
  AOI22_X1 U74 ( .A1(S0[20]), .A2(n241), .B1(S1[20]), .B2(n244), .ZN(n45) );
  INV_X1 U75 ( .A(n65), .ZN(Y[0]) );
  AOI22_X1 U76 ( .A1(S0[0]), .A2(n240), .B1(S1[0]), .B2(n249), .ZN(n65) );
  INV_X1 U77 ( .A(n64), .ZN(Y[1]) );
  AOI22_X1 U78 ( .A1(S0[1]), .A2(n240), .B1(S1[1]), .B2(n249), .ZN(n64) );
endmodule


module REGISTER_FILE_WIDTH32_LENGTH5 ( CLK, RST, EN, RD1, RD2, WR, DATAIN, 
        OUT1, OUT2, ADD_WR, ADD_RD1, ADD_RD2 );
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input CLK, RST, EN, RD1, RD2, WR;
  wire   n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8411, n8413, n8415, n8417,
         n8419, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8461, n8463, n8465, n8467, n8469,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8565,
         n8567, n8569, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573;

  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n3626), .CK(CLK), .Q(n9600), .QN(n11847)
         );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n3625), .CK(CLK), .Q(n9597), .QN(n11846)
         );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n3624), .CK(CLK), .Q(n9594), .QN(n11845)
         );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n3623), .CK(CLK), .Q(n9591), .QN(n11844)
         );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n3622), .CK(CLK), .Q(n9588), .QN(n11843)
         );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n3621), .CK(CLK), .Q(n9585), .QN(n11842)
         );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n3620), .CK(CLK), .Q(n9582), .QN(n11841)
         );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n3619), .CK(CLK), .Q(n8521), .QN(n11840)
         );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n3618), .CK(CLK), .Q(n8518), .QN(n11959)
         );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n3617), .CK(CLK), .Q(n8517), .QN(n11958)
         );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n3616), .CK(CLK), .Q(n8516), .QN(n11957)
         );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n3615), .CK(CLK), .Q(n8515), .QN(n11956)
         );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n3614), .CK(CLK), .Q(n8514), .QN(n11955)
         );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n3613), .CK(CLK), .Q(n8513), .QN(n11954)
         );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n3612), .CK(CLK), .Q(n8512), .QN(n11953)
         );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n3611), .CK(CLK), .Q(n8511), .QN(n11952)
         );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n3610), .CK(CLK), .Q(n8510), .QN(n11951)
         );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n3609), .CK(CLK), .Q(n8509), .QN(n11950)
         );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n3608), .CK(CLK), .Q(n8508), .QN(n11949)
         );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n3607), .CK(CLK), .Q(n8507), .QN(n11948)
         );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n3606), .CK(CLK), .Q(n8506), .QN(n11866)
         );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n3605), .CK(CLK), .Q(n8505), .QN(n11865)
         );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n3604), .CK(CLK), .Q(n8504), .QN(n11864)
         );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n3603), .CK(CLK), .Q(n8503), .QN(n11863)
         );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n3602), .CK(CLK), .Q(n11518), .QN(n9983)
         );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n3601), .CK(CLK), .Q(n11514), .QN(n9982)
         );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n3600), .CK(CLK), .Q(n11510), .QN(n9981)
         );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n3599), .CK(CLK), .Q(n11506), .QN(n9980)
         );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n3598), .CK(CLK), .Q(n11502), .QN(n9979)
         );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n3597), .CK(CLK), .Q(n11498), .QN(n9978)
         );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n3596), .CK(CLK), .Q(n11494), .QN(n9977)
         );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n3595), .CK(CLK), .Q(n11490), .QN(n9976)
         );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n3594), .CK(CLK), .Q(n9912), .QN(n11783)
         );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n3593), .CK(CLK), .Q(n9909), .QN(n11782)
         );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n3592), .CK(CLK), .Q(n9906), .QN(n11781)
         );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n3591), .CK(CLK), .Q(n9903), .QN(n11780)
         );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n3590), .CK(CLK), .Q(n9900), .QN(n11779)
         );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n3589), .CK(CLK), .Q(n9897), .QN(n11778)
         );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n3588), .CK(CLK), .Q(n9894), .QN(n11777)
         );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n3587), .CK(CLK), .Q(n8065), .QN(n11776)
         );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n3586), .CK(CLK), .Q(n8062), .QN(n11775)
         );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n3585), .CK(CLK), .Q(n8061), .QN(n11774)
         );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n3584), .CK(CLK), .Q(n8060), .QN(n11703)
         );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n3583), .CK(CLK), .Q(n8059), .QN(n11702)
         );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n3582), .CK(CLK), .Q(n8058), .QN(n11701)
         );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n3581), .CK(CLK), .Q(n8057), .QN(n11700)
         );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n3580), .CK(CLK), .Q(n8056), .QN(n11699)
         );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n3579), .CK(CLK), .Q(n8055), .QN(n11698)
         );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n3578), .CK(CLK), .Q(n8054), .QN(n11697)
         );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n3577), .CK(CLK), .Q(n8053), .QN(n11696)
         );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n3576), .CK(CLK), .Q(n8052), .QN(n11695)
         );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n3575), .CK(CLK), .Q(n8051), .QN(n11694)
         );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n3574), .CK(CLK), .Q(n8050), .QN(n11693)
         );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n3573), .CK(CLK), .Q(n8049), .QN(n11692)
         );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n3572), .CK(CLK), .Q(n8048), .QN(n11691)
         );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n3571), .CK(CLK), .Q(n8047), .QN(n11690)
         );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n3570), .CK(CLK), .Q(n8046), .QN(n11689)
         );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n3569), .CK(CLK), .Q(n8045), .QN(n11688)
         );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n3568), .CK(CLK), .Q(n8044), .QN(n11687)
         );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n3567), .CK(CLK), .Q(n8043), .QN(n11686)
         );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n3566), .CK(CLK), .Q(n8042), .QN(n11685)
         );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n3565), .CK(CLK), .Q(n8041), .QN(n11684)
         );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n3564), .CK(CLK), .Q(n8040), .QN(n11683)
         );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n3563), .CK(CLK), .Q(n8039), .QN(n11682)
         );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n4273), .CK(CLK), .QN(n11051) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n4274), .CK(CLK), .QN(n11049) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n4275), .CK(CLK), .QN(n11047) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n4276), .CK(CLK), .QN(n11045) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n4277), .CK(CLK), .QN(n11043) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n4278), .CK(CLK), .QN(n11041) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n4279), .CK(CLK), .QN(n11039) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n4280), .CK(CLK), .QN(n11037) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n4281), .CK(CLK), .QN(n11191) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n4282), .CK(CLK), .QN(n11187) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n4283), .CK(CLK), .QN(n11183) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n4284), .CK(CLK), .QN(n11179) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n4285), .CK(CLK), .QN(n11175) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n4286), .CK(CLK), .QN(n11170) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n4287), .CK(CLK), .QN(n11165) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n4288), .CK(CLK), .QN(n11160) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n4289), .CK(CLK), .QN(n11155) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n4290), .CK(CLK), .QN(n11150) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n4291), .CK(CLK), .QN(n11145) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n4292), .CK(CLK), .QN(n11140) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n4293), .CK(CLK), .QN(n11135) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n4294), .CK(CLK), .QN(n11130) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n4295), .CK(CLK), .QN(n11125) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n4296), .CK(CLK), .QN(n11120) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n4297), .CK(CLK), .QN(n11116) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n4298), .CK(CLK), .QN(n11112) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n4299), .CK(CLK), .QN(n11108) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n4300), .CK(CLK), .QN(n11104) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n4301), .CK(CLK), .QN(n11100) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n4302), .CK(CLK), .QN(n11096) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n4303), .CK(CLK), .QN(n11092) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n4304), .CK(CLK), .QN(n11088) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n4305), .CK(CLK), .QN(n11307) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n4306), .CK(CLK), .QN(n11305) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n4307), .CK(CLK), .QN(n11303) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n4308), .CK(CLK), .QN(n11301) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n4309), .CK(CLK), .QN(n11299) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n4310), .CK(CLK), .QN(n11297) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n4311), .CK(CLK), .QN(n11295) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n4312), .CK(CLK), .QN(n11293) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n4313), .CK(CLK), .QN(n11447) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n4314), .CK(CLK), .QN(n11443) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n4315), .CK(CLK), .QN(n11439) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n4316), .CK(CLK), .QN(n11435) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n4317), .CK(CLK), .QN(n11431) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n4318), .CK(CLK), .QN(n11426) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n4319), .CK(CLK), .QN(n11421) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n4320), .CK(CLK), .QN(n11416) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n4321), .CK(CLK), .QN(n11411) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n4322), .CK(CLK), .QN(n11406) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n4323), .CK(CLK), .QN(n11401) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n4324), .CK(CLK), .QN(n11396) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n4325), .CK(CLK), .QN(n11391) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n4326), .CK(CLK), .QN(n11386) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n4327), .CK(CLK), .QN(n11381) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n4328), .CK(CLK), .QN(n11376) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n4329), .CK(CLK), .QN(n11372) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n4330), .CK(CLK), .QN(n11368) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n4331), .CK(CLK), .QN(n11364) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n4332), .CK(CLK), .QN(n11360) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n4333), .CK(CLK), .QN(n11356) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n4334), .CK(CLK), .QN(n11352) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n4335), .CK(CLK), .QN(n11348) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n4336), .CK(CLK), .QN(n11344) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n3498), .CK(CLK), .Q(n9572), .QN(n11839)
         );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n3497), .CK(CLK), .Q(n9570), .QN(n11838)
         );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n3496), .CK(CLK), .Q(n9568), .QN(n11837)
         );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n3495), .CK(CLK), .Q(n9566), .QN(n11836)
         );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n3494), .CK(CLK), .Q(n9564), .QN(n11835)
         );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n3493), .CK(CLK), .Q(n9562), .QN(n11834)
         );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n3492), .CK(CLK), .Q(n9560), .QN(n11833)
         );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n3491), .CK(CLK), .Q(n8520), .QN(n11832)
         );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n3490), .CK(CLK), .Q(n8493), .QN(n11947)
         );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n3489), .CK(CLK), .Q(n8492), .QN(n11946)
         );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n3488), .CK(CLK), .Q(n8491), .QN(n11945)
         );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n3487), .CK(CLK), .Q(n8490), .QN(n11944)
         );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n3486), .CK(CLK), .Q(n8489), .QN(n11943)
         );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n3485), .CK(CLK), .Q(n8488), .QN(n11942)
         );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n3484), .CK(CLK), .Q(n8487), .QN(n11941)
         );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n3483), .CK(CLK), .Q(n8486), .QN(n11940)
         );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n3482), .CK(CLK), .Q(n8485), .QN(n11939)
         );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n3481), .CK(CLK), .Q(n8484), .QN(n11938)
         );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n3480), .CK(CLK), .Q(n8483), .QN(n11937)
         );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n3479), .CK(CLK), .Q(n8482), .QN(n11936)
         );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n3478), .CK(CLK), .Q(n8481), .QN(n11862)
         );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n3477), .CK(CLK), .Q(n8480), .QN(n11861)
         );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n3476), .CK(CLK), .Q(n8479), .QN(n11860)
         );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n3475), .CK(CLK), .Q(n8478), .QN(n11859)
         );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n3474), .CK(CLK), .Q(n11484), .QN(n9975)
         );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n3473), .CK(CLK), .Q(n11482), .QN(n9974)
         );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n3472), .CK(CLK), .Q(n11480), .QN(n9973)
         );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n3471), .CK(CLK), .Q(n11478), .QN(n9972)
         );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n3470), .CK(CLK), .Q(n11476), .QN(n9971)
         );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n3469), .CK(CLK), .Q(n11474), .QN(n9970)
         );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n3468), .CK(CLK), .Q(n11472), .QN(n9969)
         );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n3467), .CK(CLK), .Q(n11470), .QN(n9968)
         );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n3466), .CK(CLK), .Q(n9884), .QN(n11773)
         );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n3465), .CK(CLK), .Q(n9882), .QN(n11772)
         );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n3464), .CK(CLK), .Q(n9880), .QN(n11771)
         );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n3463), .CK(CLK), .Q(n9878), .QN(n11770)
         );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n3462), .CK(CLK), .Q(n9876), .QN(n11769)
         );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n3461), .CK(CLK), .Q(n9874), .QN(n11768)
         );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n3460), .CK(CLK), .Q(n9872), .QN(n11767)
         );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n3459), .CK(CLK), .Q(n8064), .QN(n11766)
         );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n3458), .CK(CLK), .Q(n8037), .QN(n11765)
         );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n3457), .CK(CLK), .Q(n8036), .QN(n11764)
         );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n3456), .CK(CLK), .Q(n8035), .QN(n11681)
         );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n3455), .CK(CLK), .Q(n8034), .QN(n11680)
         );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n3454), .CK(CLK), .Q(n8033), .QN(n11679)
         );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n3453), .CK(CLK), .Q(n8032), .QN(n11678)
         );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n3452), .CK(CLK), .Q(n8031), .QN(n11677)
         );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n3451), .CK(CLK), .Q(n8030), .QN(n11676)
         );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n3450), .CK(CLK), .Q(n8029), .QN(n11675)
         );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n3449), .CK(CLK), .Q(n8028), .QN(n11674)
         );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n3448), .CK(CLK), .Q(n8027), .QN(n11673)
         );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n3447), .CK(CLK), .Q(n8026), .QN(n11672)
         );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n3446), .CK(CLK), .Q(n8025), .QN(n11671)
         );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n3445), .CK(CLK), .Q(n8024), .QN(n11670)
         );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n3444), .CK(CLK), .Q(n8023), .QN(n11669)
         );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n3443), .CK(CLK), .Q(n8022), .QN(n11668)
         );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n3442), .CK(CLK), .Q(n8021), .QN(n11667)
         );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n3441), .CK(CLK), .Q(n8020), .QN(n11666)
         );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n3440), .CK(CLK), .Q(n8019), .QN(n11665)
         );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n3439), .CK(CLK), .Q(n8018), .QN(n11664)
         );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n3438), .CK(CLK), .Q(n8017), .QN(n11663)
         );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n3437), .CK(CLK), .Q(n8016), .QN(n11662)
         );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n3436), .CK(CLK), .Q(n8015), .QN(n11661)
         );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n3435), .CK(CLK), .Q(n8014), .QN(n11660)
         );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n4337), .CK(CLK), .QN(n11068) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n4338), .CK(CLK), .QN(n11067) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n4339), .CK(CLK), .QN(n11066) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n4340), .CK(CLK), .QN(n11065) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n4341), .CK(CLK), .QN(n11064) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n4342), .CK(CLK), .QN(n11063) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n4343), .CK(CLK), .QN(n11062) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n4344), .CK(CLK), .QN(n11061) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n4345), .CK(CLK), .QN(n11012) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n4346), .CK(CLK), .QN(n11011) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n4347), .CK(CLK), .QN(n11010) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n4348), .CK(CLK), .QN(n11009) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n4349), .CK(CLK), .QN(n11008) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n4350), .CK(CLK), .QN(n11007) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n4351), .CK(CLK), .QN(n11006) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n4352), .CK(CLK), .QN(n11005) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n4353), .CK(CLK), .QN(n11004) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n4354), .CK(CLK), .QN(n11003) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n4355), .CK(CLK), .QN(n11002) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n4356), .CK(CLK), .QN(n11001) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n4357), .CK(CLK), .QN(n11000) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n4358), .CK(CLK), .QN(n10999) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n4359), .CK(CLK), .QN(n10998) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n4360), .CK(CLK), .QN(n10997) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n4361), .CK(CLK), .QN(n11035) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n4362), .CK(CLK), .QN(n11033) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n4363), .CK(CLK), .QN(n11031) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n4364), .CK(CLK), .QN(n11029) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n4365), .CK(CLK), .QN(n11027) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n4366), .CK(CLK), .QN(n11025) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n4367), .CK(CLK), .QN(n11023) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n4368), .CK(CLK), .QN(n11021) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n4369), .CK(CLK), .QN(n11324) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n4370), .CK(CLK), .QN(n11323) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n4371), .CK(CLK), .QN(n11322) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n4372), .CK(CLK), .QN(n11321) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n4373), .CK(CLK), .QN(n11320) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n4374), .CK(CLK), .QN(n11319) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n4375), .CK(CLK), .QN(n11318) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n4376), .CK(CLK), .QN(n11317) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n4377), .CK(CLK), .QN(n11268) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n4378), .CK(CLK), .QN(n11267) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n4379), .CK(CLK), .QN(n11266) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n4380), .CK(CLK), .QN(n11265) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n4381), .CK(CLK), .QN(n11264) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n4382), .CK(CLK), .QN(n11263) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n4383), .CK(CLK), .QN(n11262) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n4384), .CK(CLK), .QN(n11261) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n4385), .CK(CLK), .QN(n11260) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n4386), .CK(CLK), .QN(n11259) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n4387), .CK(CLK), .QN(n11258) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n4388), .CK(CLK), .QN(n11257) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n4389), .CK(CLK), .QN(n11256) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n4390), .CK(CLK), .QN(n11255) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n4391), .CK(CLK), .QN(n11254) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n4392), .CK(CLK), .QN(n11253) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n4393), .CK(CLK), .QN(n11291) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n4394), .CK(CLK), .QN(n11289) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n4395), .CK(CLK), .QN(n11287) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n4396), .CK(CLK), .QN(n11285) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n4397), .CK(CLK), .QN(n11283) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n4398), .CK(CLK), .QN(n11281) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n4399), .CK(CLK), .QN(n11279) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n4400), .CK(CLK), .QN(n11277) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n3370), .CK(CLK), .QN(n11316) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n3369), .CK(CLK), .QN(n11315) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n3368), .CK(CLK), .QN(n11314) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n3367), .CK(CLK), .QN(n11313) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n3366), .CK(CLK), .QN(n11312) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n3365), .CK(CLK), .QN(n11311) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n3364), .CK(CLK), .QN(n11310) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n3363), .CK(CLK), .QN(n11309) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n3362), .CK(CLK), .QN(n11231) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n3361), .CK(CLK), .QN(n11230) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n3360), .CK(CLK), .QN(n11229) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n3359), .CK(CLK), .QN(n11228) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n3358), .CK(CLK), .QN(n11227) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n3357), .CK(CLK), .QN(n11226) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n3356), .CK(CLK), .QN(n11225) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n3355), .CK(CLK), .QN(n11224) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n3354), .CK(CLK), .QN(n11223) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n3353), .CK(CLK), .QN(n11222) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n3352), .CK(CLK), .QN(n11221) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n3351), .CK(CLK), .QN(n11220) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n3350), .CK(CLK), .QN(n11219) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n3349), .CK(CLK), .QN(n11218) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n3348), .CK(CLK), .QN(n11217) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n3347), .CK(CLK), .QN(n11216) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n3346), .CK(CLK), .QN(n11246) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n3345), .CK(CLK), .QN(n11245) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n3344), .CK(CLK), .QN(n11244) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n3343), .CK(CLK), .QN(n11243) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n3342), .CK(CLK), .QN(n11242) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n3341), .CK(CLK), .QN(n11241) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n3340), .CK(CLK), .QN(n11240) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n3339), .CK(CLK), .QN(n11239) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n3338), .CK(CLK), .QN(n11060) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n3337), .CK(CLK), .QN(n11059) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n3336), .CK(CLK), .QN(n11058) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n3335), .CK(CLK), .QN(n11057) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n3334), .CK(CLK), .QN(n11056) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n3333), .CK(CLK), .QN(n11055) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n3332), .CK(CLK), .QN(n11054) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n3331), .CK(CLK), .QN(n11053) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n3330), .CK(CLK), .QN(n10975) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n3329), .CK(CLK), .QN(n10974) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n3328), .CK(CLK), .QN(n10973) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n3327), .CK(CLK), .QN(n10972) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n3326), .CK(CLK), .QN(n10971) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n3325), .CK(CLK), .QN(n10970) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n3324), .CK(CLK), .QN(n10969) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n3323), .CK(CLK), .QN(n10968) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n3322), .CK(CLK), .QN(n10967) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n3321), .CK(CLK), .QN(n10966) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n3320), .CK(CLK), .QN(n10965) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n3319), .CK(CLK), .QN(n10964) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n3318), .CK(CLK), .QN(n10963) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n3317), .CK(CLK), .QN(n10962) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n3316), .CK(CLK), .QN(n10961) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n3315), .CK(CLK), .QN(n10960) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n3314), .CK(CLK), .QN(n10990) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n3313), .CK(CLK), .QN(n10989) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n3312), .CK(CLK), .QN(n10988) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n3311), .CK(CLK), .QN(n10987) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n3310), .CK(CLK), .QN(n10986) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n3309), .CK(CLK), .QN(n10985) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n3308), .CK(CLK), .QN(n10984) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n3307), .CK(CLK), .QN(n10983) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n3306), .CK(CLK), .Q(n9911), .QN(n11763)
         );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n3305), .CK(CLK), .Q(n9908), .QN(n11762)
         );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n3304), .CK(CLK), .Q(n9905), .QN(n11761)
         );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n3303), .CK(CLK), .Q(n9902), .QN(n11760)
         );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n3302), .CK(CLK), .Q(n9899), .QN(n11759)
         );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n3301), .CK(CLK), .Q(n9896), .QN(n11758)
         );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n3300), .CK(CLK), .Q(n9893), .QN(n11757)
         );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n3299), .CK(CLK), .Q(n8013), .QN(n11756)
         );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n3298), .CK(CLK), .Q(n8011), .QN(n11755)
         );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n3297), .CK(CLK), .Q(n8009), .QN(n11754)
         );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n3296), .CK(CLK), .Q(n8007), .QN(n11659)
         );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n3295), .CK(CLK), .Q(n8005), .QN(n11658)
         );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n3294), .CK(CLK), .Q(n8003), .QN(n11657)
         );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n3293), .CK(CLK), .Q(n8001), .QN(n11656)
         );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n3292), .CK(CLK), .Q(n7999), .QN(n11655)
         );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n3291), .CK(CLK), .Q(n7997), .QN(n11654)
         );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n3290), .CK(CLK), .Q(n7995), .QN(n11653)
         );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n3289), .CK(CLK), .Q(n7993), .QN(n11652)
         );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n3288), .CK(CLK), .Q(n7991), .QN(n11651)
         );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n3287), .CK(CLK), .Q(n7989), .QN(n11650)
         );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n3286), .CK(CLK), .Q(n7987), .QN(n11649)
         );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n3285), .CK(CLK), .Q(n7985), .QN(n11648)
         );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n3284), .CK(CLK), .Q(n7983), .QN(n11647)
         );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n3283), .CK(CLK), .Q(n7981), .QN(n11646)
         );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n3282), .CK(CLK), .Q(n7979), .QN(n11645)
         );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n3281), .CK(CLK), .Q(n7977), .QN(n11644)
         );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n3280), .CK(CLK), .Q(n7975), .QN(n11643)
         );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n3279), .CK(CLK), .Q(n7973), .QN(n11642)
         );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n3278), .CK(CLK), .Q(n7971), .QN(n11641)
         );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n3277), .CK(CLK), .Q(n7969), .QN(n11640)
         );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n3276), .CK(CLK), .Q(n7967), .QN(n11639)
         );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n3275), .CK(CLK), .Q(n7965), .QN(n11638)
         );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n3274), .CK(CLK), .Q(n9599), .QN(n11831)
         );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n3273), .CK(CLK), .Q(n9596), .QN(n11830)
         );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n3272), .CK(CLK), .Q(n9593), .QN(n11829)
         );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n3271), .CK(CLK), .Q(n9590), .QN(n11828)
         );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n3270), .CK(CLK), .Q(n9587), .QN(n11827)
         );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n3269), .CK(CLK), .Q(n9584), .QN(n11826)
         );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n3268), .CK(CLK), .Q(n9581), .QN(n11825)
         );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n3267), .CK(CLK), .Q(n8469), .QN(n11824)
         );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n3266), .CK(CLK), .Q(n8467), .QN(n11935)
         );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n3265), .CK(CLK), .Q(n8465), .QN(n11934)
         );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n3264), .CK(CLK), .Q(n8463), .QN(n11933)
         );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n3263), .CK(CLK), .Q(n8461), .QN(n11932)
         );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n3262), .CK(CLK), .Q(n8459), .QN(n11931)
         );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n3261), .CK(CLK), .Q(n8457), .QN(n11930)
         );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n3260), .CK(CLK), .Q(n8455), .QN(n11929)
         );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n3259), .CK(CLK), .Q(n8453), .QN(n11928)
         );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n3258), .CK(CLK), .Q(n8451), .QN(n11927)
         );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n3257), .CK(CLK), .Q(n8449), .QN(n11926)
         );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n3256), .CK(CLK), .Q(n8447), .QN(n11925)
         );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n3255), .CK(CLK), .Q(n8445), .QN(n11924)
         );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n3254), .CK(CLK), .Q(n8443), .QN(n11858)
         );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n3253), .CK(CLK), .Q(n8441), .QN(n11857)
         );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n3252), .CK(CLK), .Q(n8439), .QN(n11856)
         );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n3251), .CK(CLK), .Q(n8437), .QN(n11855)
         );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n3250), .CK(CLK), .Q(n11463), .QN(n9967)
         );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n3249), .CK(CLK), .Q(n11462), .QN(n9966)
         );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n3248), .CK(CLK), .Q(n11461), .QN(n9965)
         );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n3247), .CK(CLK), .Q(n11460), .QN(n9964)
         );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n3246), .CK(CLK), .Q(n11459), .QN(n9963)
         );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n3245), .CK(CLK), .Q(n11458), .QN(n9962)
         );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n3244), .CK(CLK), .Q(n11457), .QN(n9961)
         );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n3243), .CK(CLK), .Q(n11456), .QN(n9960)
         );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n3242), .CK(CLK), .QN(n11339) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n3241), .CK(CLK), .QN(n11337) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n3240), .CK(CLK), .QN(n11335) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n3239), .CK(CLK), .QN(n11333) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n3238), .CK(CLK), .QN(n11331) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n3237), .CK(CLK), .QN(n11329) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n3236), .CK(CLK), .QN(n11327) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n3235), .CK(CLK), .QN(n11325) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n3234), .CK(CLK), .QN(n11206) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n3233), .CK(CLK), .QN(n11205) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n3232), .CK(CLK), .QN(n11204) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n3231), .CK(CLK), .QN(n11203) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n3230), .CK(CLK), .QN(n11202) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n3229), .CK(CLK), .QN(n11201) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n3228), .CK(CLK), .QN(n11200) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n3227), .CK(CLK), .QN(n11199) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n3226), .CK(CLK), .QN(n11198) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n3225), .CK(CLK), .QN(n11197) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n3224), .CK(CLK), .QN(n11196) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n3223), .CK(CLK), .QN(n11195) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n3222), .CK(CLK), .QN(n11194) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n3221), .CK(CLK), .QN(n11193) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n3220), .CK(CLK), .QN(n11192) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n3219), .CK(CLK), .QN(n11375) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n3218), .CK(CLK), .QN(n11214) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n3217), .CK(CLK), .QN(n11213) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n3216), .CK(CLK), .QN(n11212) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n3215), .CK(CLK), .QN(n11211) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n3214), .CK(CLK), .QN(n11210) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n3213), .CK(CLK), .QN(n11209) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n3212), .CK(CLK), .QN(n11208) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n3211), .CK(CLK), .QN(n11207) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n3210), .CK(CLK), .QN(n11083) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n3209), .CK(CLK), .QN(n11081) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n3208), .CK(CLK), .QN(n11079) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n3207), .CK(CLK), .QN(n11077) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n3206), .CK(CLK), .QN(n11075) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n3205), .CK(CLK), .QN(n11073) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n3204), .CK(CLK), .QN(n11071) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n3203), .CK(CLK), .QN(n11069) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n3202), .CK(CLK), .QN(n10950) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n3201), .CK(CLK), .QN(n10949) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n3200), .CK(CLK), .QN(n10948) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n3199), .CK(CLK), .QN(n10947) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n3198), .CK(CLK), .QN(n10946) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n3197), .CK(CLK), .QN(n10945) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n3196), .CK(CLK), .QN(n10944) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n3195), .CK(CLK), .QN(n10943) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n3194), .CK(CLK), .QN(n10942) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n3193), .CK(CLK), .QN(n10941) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n3192), .CK(CLK), .QN(n10940) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n3191), .CK(CLK), .QN(n10939) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n3190), .CK(CLK), .QN(n10938) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n3189), .CK(CLK), .QN(n10937) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n3188), .CK(CLK), .QN(n10936) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n3187), .CK(CLK), .QN(n11119) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n3186), .CK(CLK), .QN(n10958) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n3185), .CK(CLK), .QN(n10957) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n3184), .CK(CLK), .QN(n10956) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n3183), .CK(CLK), .QN(n10955) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n3182), .CK(CLK), .QN(n10954) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n3181), .CK(CLK), .QN(n10953) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n3180), .CK(CLK), .QN(n10952) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n3179), .CK(CLK), .QN(n10951) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n3178), .CK(CLK), .Q(n9870), .QN(n11753)
         );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n3177), .CK(CLK), .Q(n9869), .QN(n11752)
         );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n3176), .CK(CLK), .Q(n9868), .QN(n11751)
         );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n3175), .CK(CLK), .Q(n9867), .QN(n11750)
         );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n3174), .CK(CLK), .Q(n9866), .QN(n11749)
         );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n3173), .CK(CLK), .Q(n9865), .QN(n11748)
         );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n3172), .CK(CLK), .Q(n9864), .QN(n11747)
         );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n3171), .CK(CLK), .Q(n7963), .QN(n11746)
         );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n3170), .CK(CLK), .Q(n7961), .QN(n11745)
         );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n3169), .CK(CLK), .Q(n7959), .QN(n11744)
         );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n3168), .CK(CLK), .Q(n7957), .QN(n11637)
         );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n3167), .CK(CLK), .Q(n7955), .QN(n11636)
         );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n3166), .CK(CLK), .Q(n7953), .QN(n11635)
         );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n3165), .CK(CLK), .Q(n7951), .QN(n11634)
         );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n3164), .CK(CLK), .Q(n7949), .QN(n11633)
         );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n3163), .CK(CLK), .Q(n7947), .QN(n11632)
         );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n3162), .CK(CLK), .Q(n7945), .QN(n11631)
         );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n3161), .CK(CLK), .Q(n7943), .QN(n11630)
         );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n3160), .CK(CLK), .Q(n7941), .QN(n11629)
         );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n3159), .CK(CLK), .Q(n7939), .QN(n11628)
         );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n3158), .CK(CLK), .Q(n7937), .QN(n11627)
         );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n3157), .CK(CLK), .Q(n7935), .QN(n11626)
         );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n3156), .CK(CLK), .Q(n7933), .QN(n11625)
         );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n3155), .CK(CLK), .Q(n7931), .QN(n11624)
         );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n3154), .CK(CLK), .Q(n7929), .QN(n11623)
         );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n3153), .CK(CLK), .Q(n7927), .QN(n11622)
         );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n3152), .CK(CLK), .Q(n7925), .QN(n11621)
         );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n3151), .CK(CLK), .Q(n7923), .QN(n11620)
         );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n3150), .CK(CLK), .Q(n7921), .QN(n11619)
         );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n3149), .CK(CLK), .Q(n7919), .QN(n11618)
         );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n3148), .CK(CLK), .Q(n7917), .QN(n11617)
         );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n3147), .CK(CLK), .Q(n7915), .QN(n11616)
         );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n3146), .CK(CLK), .Q(n9558), .QN(n11823)
         );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n3145), .CK(CLK), .Q(n9557), .QN(n11822)
         );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n3144), .CK(CLK), .Q(n9556), .QN(n11821)
         );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n3143), .CK(CLK), .Q(n9555), .QN(n11820)
         );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n3142), .CK(CLK), .Q(n9554), .QN(n11819)
         );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n3141), .CK(CLK), .Q(n9553), .QN(n11818)
         );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n3140), .CK(CLK), .Q(n9552), .QN(n11817)
         );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n3139), .CK(CLK), .Q(n8419), .QN(n11816)
         );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n3138), .CK(CLK), .Q(n8417), .QN(n11923)
         );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n3137), .CK(CLK), .Q(n8415), .QN(n11922)
         );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n3136), .CK(CLK), .Q(n8413), .QN(n11921)
         );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n3135), .CK(CLK), .Q(n8411), .QN(n11920)
         );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n3134), .CK(CLK), .Q(n8409), .QN(n11919)
         );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n3133), .CK(CLK), .Q(n8407), .QN(n11918)
         );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n3132), .CK(CLK), .Q(n8405), .QN(n11917)
         );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n3131), .CK(CLK), .Q(n8403), .QN(n11916)
         );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n3130), .CK(CLK), .Q(n8401), .QN(n11915)
         );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n3129), .CK(CLK), .Q(n8399), .QN(n11914)
         );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n3128), .CK(CLK), .Q(n8397), .QN(n11913)
         );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n3127), .CK(CLK), .Q(n8395), .QN(n11912)
         );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n3126), .CK(CLK), .Q(n8393), .QN(n11854)
         );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n3125), .CK(CLK), .Q(n8391), .QN(n11853)
         );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n3124), .CK(CLK), .Q(n8389), .QN(n11852)
         );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n3123), .CK(CLK), .Q(n8387), .QN(n11851)
         );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n3122), .CK(CLK), .Q(n11455), .QN(n9959)
         );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n3121), .CK(CLK), .Q(n11454), .QN(n9958)
         );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n3120), .CK(CLK), .Q(n11453), .QN(n9957)
         );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n3119), .CK(CLK), .Q(n11452), .QN(n9956)
         );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n3118), .CK(CLK), .Q(n11451), .QN(n9955)
         );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n3117), .CK(CLK), .Q(n11450), .QN(n9954)
         );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n3116), .CK(CLK), .Q(n11449), .QN(n9953)
         );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n3115), .CK(CLK), .Q(n11448), .QN(n9952)
         );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n3114), .CK(CLK), .QN(n11308) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n3113), .CK(CLK), .QN(n11306) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n3112), .CK(CLK), .QN(n11304) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n3111), .CK(CLK), .QN(n11302) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n3110), .CK(CLK), .QN(n11300) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n3109), .CK(CLK), .QN(n11298) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n3108), .CK(CLK), .QN(n11296) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n3107), .CK(CLK), .QN(n11294) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n3106), .CK(CLK), .QN(n11446) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n3105), .CK(CLK), .QN(n11442) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n3104), .CK(CLK), .QN(n11438) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n3103), .CK(CLK), .QN(n11434) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n3102), .CK(CLK), .QN(n11430) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n3101), .CK(CLK), .QN(n11425) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n3100), .CK(CLK), .QN(n11420) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n3099), .CK(CLK), .QN(n11415) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n3098), .CK(CLK), .QN(n11410) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n3097), .CK(CLK), .QN(n11405) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n3096), .CK(CLK), .QN(n11400) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n3095), .CK(CLK), .QN(n11395) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n3094), .CK(CLK), .QN(n11390) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n3093), .CK(CLK), .QN(n11385) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n3092), .CK(CLK), .QN(n11380) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n3091), .CK(CLK), .QN(n11374) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n3090), .CK(CLK), .QN(n11371) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n3089), .CK(CLK), .QN(n11367) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n3088), .CK(CLK), .QN(n11363) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n3087), .CK(CLK), .QN(n11359) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n3086), .CK(CLK), .QN(n11355) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n3085), .CK(CLK), .QN(n11351) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n3084), .CK(CLK), .QN(n11347) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n3083), .CK(CLK), .QN(n11343) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n3082), .CK(CLK), .QN(n11052) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n3081), .CK(CLK), .QN(n11050) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n3080), .CK(CLK), .QN(n11048) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n3079), .CK(CLK), .QN(n11046) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n3078), .CK(CLK), .QN(n11044) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n3077), .CK(CLK), .QN(n11042) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n3076), .CK(CLK), .QN(n11040) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n3075), .CK(CLK), .QN(n11038) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n3074), .CK(CLK), .QN(n11190) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n3073), .CK(CLK), .QN(n11186) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n3072), .CK(CLK), .QN(n11182) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n3071), .CK(CLK), .QN(n11178) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n3070), .CK(CLK), .QN(n11174) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n3069), .CK(CLK), .QN(n11169) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n3068), .CK(CLK), .QN(n11164) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n3067), .CK(CLK), .QN(n11159) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n3066), .CK(CLK), .QN(n11154) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n3065), .CK(CLK), .QN(n11149) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n3064), .CK(CLK), .QN(n11144) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n3063), .CK(CLK), .QN(n11139) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n3062), .CK(CLK), .QN(n11134) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n3061), .CK(CLK), .QN(n11129) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n3060), .CK(CLK), .QN(n11124) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n3059), .CK(CLK), .QN(n11118) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n3058), .CK(CLK), .QN(n11115) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n3057), .CK(CLK), .QN(n11111) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n3056), .CK(CLK), .QN(n11107) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n3055), .CK(CLK), .QN(n11103) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n3054), .CK(CLK), .QN(n11099) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n3053), .CK(CLK), .QN(n11095) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n3052), .CK(CLK), .QN(n11091) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n3051), .CK(CLK), .QN(n11087) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n3050), .CK(CLK), .Q(n9910), .QN(n11743)
         );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n3049), .CK(CLK), .Q(n9907), .QN(n11742)
         );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n3048), .CK(CLK), .Q(n9904), .QN(n11741)
         );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n3047), .CK(CLK), .Q(n9901), .QN(n11740)
         );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n3046), .CK(CLK), .Q(n9898), .QN(n11739)
         );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n3045), .CK(CLK), .Q(n9895), .QN(n11738)
         );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n3044), .CK(CLK), .Q(n9892), .QN(n11737)
         );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n3043), .CK(CLK), .Q(n8063), .QN(n11736)
         );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n3042), .CK(CLK), .Q(n8113), .QN(n11735)
         );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n3041), .CK(CLK), .Q(n8111), .QN(n11734)
         );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n3040), .CK(CLK), .Q(n8109), .QN(n11615)
         );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n3039), .CK(CLK), .Q(n8107), .QN(n11614)
         );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n3038), .CK(CLK), .Q(n8105), .QN(n11613)
         );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n3037), .CK(CLK), .Q(n8103), .QN(n11612)
         );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n3036), .CK(CLK), .Q(n8101), .QN(n11611)
         );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n3035), .CK(CLK), .Q(n8099), .QN(n11610)
         );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n3034), .CK(CLK), .Q(n8097), .QN(n11609)
         );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n3033), .CK(CLK), .Q(n8095), .QN(n11608)
         );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n3032), .CK(CLK), .Q(n8093), .QN(n11607)
         );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n3031), .CK(CLK), .Q(n8091), .QN(n11606)
         );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n3030), .CK(CLK), .Q(n8089), .QN(n11605)
         );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n3029), .CK(CLK), .Q(n8087), .QN(n11604)
         );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n3028), .CK(CLK), .Q(n8085), .QN(n11603)
         );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n3027), .CK(CLK), .Q(n8083), .QN(n11602)
         );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n3026), .CK(CLK), .Q(n8081), .QN(n11601)
         );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n3025), .CK(CLK), .Q(n8079), .QN(n11600)
         );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n3024), .CK(CLK), .Q(n8077), .QN(n11599)
         );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n3023), .CK(CLK), .Q(n8075), .QN(n11598)
         );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n3022), .CK(CLK), .Q(n8073), .QN(n11597)
         );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n3021), .CK(CLK), .Q(n8071), .QN(n11596)
         );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n3020), .CK(CLK), .Q(n8069), .QN(n11595)
         );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n3019), .CK(CLK), .Q(n8067), .QN(n11594)
         );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n3018), .CK(CLK), .Q(n9598), .QN(n11911)
         );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n3017), .CK(CLK), .Q(n9595), .QN(n11850)
         );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n3016), .CK(CLK), .Q(n9592), .QN(n11849)
         );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n3015), .CK(CLK), .Q(n9589), .QN(n11910)
         );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n3014), .CK(CLK), .Q(n9586), .QN(n11909)
         );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n3013), .CK(CLK), .Q(n9583), .QN(n11908)
         );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n3012), .CK(CLK), .Q(n9580), .QN(n11907)
         );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n3011), .CK(CLK), .Q(n8519), .QN(n11906)
         );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n3010), .CK(CLK), .Q(n8569), .QN(n11905)
         );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n3009), .CK(CLK), .Q(n8567), .QN(n11904)
         );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n3008), .CK(CLK), .Q(n8565), .QN(n11903)
         );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n3007), .CK(CLK), .Q(n11521), .QN(n9999)
         );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n3006), .CK(CLK), .Q(n8561), .QN(n11902)
         );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n3005), .CK(CLK), .Q(n8559), .QN(n11901)
         );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n3004), .CK(CLK), .Q(n8557), .QN(n11900)
         );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n3003), .CK(CLK), .Q(n8555), .QN(n11815)
         );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n3002), .CK(CLK), .Q(n8553), .QN(n11814)
         );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n3001), .CK(CLK), .Q(n8551), .QN(n11813)
         );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n3000), .CK(CLK), .Q(n8549), .QN(n11812)
         );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n2999), .CK(CLK), .Q(n8547), .QN(n11811)
         );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n2998), .CK(CLK), .Q(n8545), .QN(n11810)
         );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n2997), .CK(CLK), .Q(n8543), .QN(n11809)
         );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n2996), .CK(CLK), .Q(n8541), .QN(n11808)
         );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n2995), .CK(CLK), .Q(n8539), .QN(n11848)
         );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n2994), .CK(CLK), .Q(n11517), .QN(n9951)
         );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n2993), .CK(CLK), .Q(n11513), .QN(n9950)
         );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n2992), .CK(CLK), .Q(n11509), .QN(n9949)
         );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n2991), .CK(CLK), .Q(n11505), .QN(n9948)
         );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n2990), .CK(CLK), .Q(n11501), .QN(n9947)
         );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n2989), .CK(CLK), .Q(n11497), .QN(n9946)
         );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n2988), .CK(CLK), .Q(n11493), .QN(n9945)
         );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n2987), .CK(CLK), .Q(n11489), .QN(n9944)
         );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n2986), .CK(CLK), .QN(n11275) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n2985), .CK(CLK), .QN(n11274) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n2984), .CK(CLK), .QN(n11273) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n2983), .CK(CLK), .QN(n11272) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n2982), .CK(CLK), .QN(n11271) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n2981), .CK(CLK), .QN(n11270) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n2980), .CK(CLK), .QN(n11269) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n2979), .CK(CLK), .QN(n11292) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n2978), .CK(CLK), .QN(n11444) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n2977), .CK(CLK), .QN(n11440) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n2976), .CK(CLK), .QN(n11436) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n2975), .CK(CLK), .QN(n11432) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n2974), .CK(CLK), .QN(n11427) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n2973), .CK(CLK), .QN(n11422) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n2972), .CK(CLK), .QN(n11417) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n2971), .CK(CLK), .QN(n11412) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n2970), .CK(CLK), .QN(n11407) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n2969), .CK(CLK), .QN(n11402) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n2968), .CK(CLK), .QN(n11397) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n2967), .CK(CLK), .QN(n11392) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n2966), .CK(CLK), .QN(n11387) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n2965), .CK(CLK), .QN(n11382) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n2964), .CK(CLK), .QN(n11377) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n2963), .CK(CLK), .QN(n11252) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n2962), .CK(CLK), .QN(n11290) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n2961), .CK(CLK), .QN(n11288) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n2960), .CK(CLK), .QN(n11286) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n2959), .CK(CLK), .QN(n11284) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n2958), .CK(CLK), .QN(n11282) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n2957), .CK(CLK), .QN(n11280) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n2956), .CK(CLK), .QN(n11278) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n2955), .CK(CLK), .QN(n11276) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n2954), .CK(CLK), .QN(n11019) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n2953), .CK(CLK), .QN(n11018) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n2952), .CK(CLK), .QN(n11017) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n2951), .CK(CLK), .QN(n11016) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n2950), .CK(CLK), .QN(n11015) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n2949), .CK(CLK), .QN(n11014) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n2948), .CK(CLK), .QN(n11013) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n2947), .CK(CLK), .QN(n11036) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n2946), .CK(CLK), .QN(n11188) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n2945), .CK(CLK), .QN(n11184) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n2944), .CK(CLK), .QN(n11180) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n2943), .CK(CLK), .QN(n11176) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n2942), .CK(CLK), .QN(n11171) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n2941), .CK(CLK), .QN(n11166) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n2940), .CK(CLK), .QN(n11161) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n2939), .CK(CLK), .QN(n11156) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n2938), .CK(CLK), .QN(n11151) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n2937), .CK(CLK), .QN(n11146) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n2936), .CK(CLK), .QN(n11141) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n2935), .CK(CLK), .QN(n11136) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n2934), .CK(CLK), .QN(n11131) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n2933), .CK(CLK), .QN(n11126) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n2932), .CK(CLK), .QN(n11121) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n2931), .CK(CLK), .QN(n10996) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n2930), .CK(CLK), .QN(n11034) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n2929), .CK(CLK), .QN(n11032) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n2928), .CK(CLK), .QN(n11030) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n2927), .CK(CLK), .QN(n11028) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n2926), .CK(CLK), .QN(n11026) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n2925), .CK(CLK), .QN(n11024) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n2924), .CK(CLK), .QN(n11022) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n2923), .CK(CLK), .QN(n11020) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n2922), .CK(CLK), .Q(n9883), .QN(n11733)
         );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n2921), .CK(CLK), .Q(n9881), .QN(n11732)
         );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n2920), .CK(CLK), .Q(n9879), .QN(n11731)
         );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n2919), .CK(CLK), .Q(n9877), .QN(n11730)
         );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n2918), .CK(CLK), .Q(n9875), .QN(n11729)
         );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n2917), .CK(CLK), .Q(n9873), .QN(n11728)
         );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n2916), .CK(CLK), .Q(n9871), .QN(n11727)
         );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n2915), .CK(CLK), .Q(n8038), .QN(n11726)
         );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n2914), .CK(CLK), .Q(n8112), .QN(n11725)
         );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n2913), .CK(CLK), .Q(n8110), .QN(n11724)
         );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n2912), .CK(CLK), .Q(n8108), .QN(n11593)
         );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n2911), .CK(CLK), .Q(n8106), .QN(n11592)
         );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n2910), .CK(CLK), .Q(n8104), .QN(n11591)
         );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n2909), .CK(CLK), .Q(n8102), .QN(n11590)
         );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n2908), .CK(CLK), .Q(n8100), .QN(n11589)
         );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n2907), .CK(CLK), .Q(n8098), .QN(n11588)
         );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n2906), .CK(CLK), .Q(n8096), .QN(n11587)
         );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n2905), .CK(CLK), .Q(n8094), .QN(n11586)
         );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n2904), .CK(CLK), .Q(n8092), .QN(n11585)
         );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n2903), .CK(CLK), .Q(n8090), .QN(n11584)
         );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n2902), .CK(CLK), .Q(n8088), .QN(n11583)
         );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n2901), .CK(CLK), .Q(n8086), .QN(n11582)
         );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n2900), .CK(CLK), .Q(n8084), .QN(n11581)
         );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n2899), .CK(CLK), .Q(n8082), .QN(n11580)
         );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n2898), .CK(CLK), .Q(n8080), .QN(n11579)
         );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n2897), .CK(CLK), .Q(n8078), .QN(n11578)
         );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n2896), .CK(CLK), .Q(n8076), .QN(n11577)
         );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n2895), .CK(CLK), .Q(n8074), .QN(n11576)
         );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n2894), .CK(CLK), .Q(n8072), .QN(n11575)
         );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n2893), .CK(CLK), .Q(n8070), .QN(n11574)
         );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n2892), .CK(CLK), .Q(n8068), .QN(n11573)
         );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n2891), .CK(CLK), .Q(n8066), .QN(n11572)
         );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n2890), .CK(CLK), .Q(n9571), .QN(n11899)
         );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n2889), .CK(CLK), .Q(n9569), .QN(n11898)
         );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n2888), .CK(CLK), .Q(n9567), .QN(n11897)
         );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n2887), .CK(CLK), .Q(n9565), .QN(n11896)
         );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n2886), .CK(CLK), .Q(n9563), .QN(n11895)
         );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n2885), .CK(CLK), .Q(n9561), .QN(n11894)
         );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n2884), .CK(CLK), .Q(n9559), .QN(n11893)
         );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n2883), .CK(CLK), .Q(n11485), .QN(n9998)
         );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n2882), .CK(CLK), .Q(n11526), .QN(n9997)
         );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n2881), .CK(CLK), .Q(n11524), .QN(n9996)
         );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n2880), .CK(CLK), .Q(n11522), .QN(n9995)
         );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n2879), .CK(CLK), .Q(n11519), .QN(n9994)
         );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n2878), .CK(CLK), .Q(n8560), .QN(n11892)
         );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n2877), .CK(CLK), .Q(n8558), .QN(n11891)
         );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n2876), .CK(CLK), .Q(n8556), .QN(n11890)
         );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n2875), .CK(CLK), .Q(n8554), .QN(n11807)
         );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n2874), .CK(CLK), .Q(n8552), .QN(n11806)
         );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n2873), .CK(CLK), .Q(n8550), .QN(n11805)
         );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n2872), .CK(CLK), .Q(n8548), .QN(n11804)
         );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n2871), .CK(CLK), .Q(n8546), .QN(n11803)
         );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n2870), .CK(CLK), .Q(n8544), .QN(n11802)
         );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n2869), .CK(CLK), .Q(n8542), .QN(n11801)
         );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n2868), .CK(CLK), .Q(n8540), .QN(n11800)
         );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n2867), .CK(CLK), .Q(n8538), .QN(n11889)
         );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n2866), .CK(CLK), .Q(n11483), .QN(n9943)
         );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n2865), .CK(CLK), .Q(n11481), .QN(n9942)
         );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n2864), .CK(CLK), .Q(n11479), .QN(n9941)
         );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n2863), .CK(CLK), .Q(n11477), .QN(n9940)
         );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n2862), .CK(CLK), .Q(n11475), .QN(n9939)
         );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n2861), .CK(CLK), .Q(n11473), .QN(n9938)
         );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n2860), .CK(CLK), .Q(n11471), .QN(n9937)
         );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n2859), .CK(CLK), .Q(n11469), .QN(n9936)
         );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n4401), .CK(CLK), .QN(n11238) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n4402), .CK(CLK), .QN(n11237) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n4403), .CK(CLK), .QN(n11236) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n4404), .CK(CLK), .QN(n11235) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n4405), .CK(CLK), .QN(n11234) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n4406), .CK(CLK), .QN(n11233) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n4407), .CK(CLK), .QN(n11232) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n4408), .CK(CLK), .QN(n11251) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n4409), .CK(CLK), .QN(n11250) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n4410), .CK(CLK), .QN(n11249) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n4411), .CK(CLK), .QN(n11248) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n4412), .CK(CLK), .QN(n11247) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n4413), .CK(CLK), .QN(n11429) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n4414), .CK(CLK), .QN(n11424) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n4415), .CK(CLK), .QN(n11419) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n4416), .CK(CLK), .QN(n11414) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n4417), .CK(CLK), .QN(n11409) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n4418), .CK(CLK), .QN(n11404) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n4419), .CK(CLK), .QN(n11399) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n4420), .CK(CLK), .QN(n11394) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n4421), .CK(CLK), .QN(n11389) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n4422), .CK(CLK), .QN(n11384) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n4423), .CK(CLK), .QN(n11379) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n4424), .CK(CLK), .QN(n11215) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n4425), .CK(CLK), .QN(n11370) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n4426), .CK(CLK), .QN(n11366) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n4427), .CK(CLK), .QN(n11362) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n4428), .CK(CLK), .QN(n11358) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n4429), .CK(CLK), .QN(n11354) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n4430), .CK(CLK), .QN(n11350) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n4431), .CK(CLK), .QN(n11346) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n4432), .CK(CLK), .QN(n11342) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n4433), .CK(CLK), .QN(n10982) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n4434), .CK(CLK), .QN(n10981) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n4435), .CK(CLK), .QN(n10980) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n4436), .CK(CLK), .QN(n10979) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n4437), .CK(CLK), .QN(n10978) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n4438), .CK(CLK), .QN(n10977) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n4439), .CK(CLK), .QN(n10976) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n4440), .CK(CLK), .QN(n10995) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n4441), .CK(CLK), .QN(n10994) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n4442), .CK(CLK), .QN(n10993) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n4443), .CK(CLK), .QN(n10992) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n4444), .CK(CLK), .QN(n10991) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n4445), .CK(CLK), .QN(n11173) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n4446), .CK(CLK), .QN(n11168) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n4447), .CK(CLK), .QN(n11163) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n4448), .CK(CLK), .QN(n11158) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n4449), .CK(CLK), .QN(n11153) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n4450), .CK(CLK), .QN(n11148) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n4451), .CK(CLK), .QN(n11143) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n4452), .CK(CLK), .QN(n11138) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n4453), .CK(CLK), .QN(n11133) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n4454), .CK(CLK), .QN(n11128) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n4455), .CK(CLK), .QN(n11123) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n4456), .CK(CLK), .QN(n10959) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n4457), .CK(CLK), .QN(n11114) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n4458), .CK(CLK), .QN(n11110) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n4459), .CK(CLK), .QN(n11106) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n4460), .CK(CLK), .QN(n11102) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n4461), .CK(CLK), .QN(n11098) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n4462), .CK(CLK), .QN(n11094) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n4463), .CK(CLK), .QN(n11090) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n4464), .CK(CLK), .QN(n11086) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n2794), .CK(CLK), .Q(n9891), .QN(n11723)
         );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n2793), .CK(CLK), .Q(n9890), .QN(n11722)
         );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n2792), .CK(CLK), .Q(n9889), .QN(n11721)
         );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n2791), .CK(CLK), .Q(n9888), .QN(n11720)
         );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n2790), .CK(CLK), .Q(n9887), .QN(n11719)
         );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n2789), .CK(CLK), .Q(n9886), .QN(n11718)
         );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n2788), .CK(CLK), .Q(n9885), .QN(n11717)
         );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n2787), .CK(CLK), .Q(n8012), .QN(n11716)
         );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n2786), .CK(CLK), .Q(n8010), .QN(n11715)
         );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n2785), .CK(CLK), .Q(n8008), .QN(n11714)
         );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n2784), .CK(CLK), .Q(n8006), .QN(n11571)
         );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n2783), .CK(CLK), .Q(n8004), .QN(n11570)
         );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n2782), .CK(CLK), .Q(n8002), .QN(n11569)
         );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n2781), .CK(CLK), .Q(n8000), .QN(n11568)
         );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n2780), .CK(CLK), .Q(n7998), .QN(n11567)
         );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n2779), .CK(CLK), .Q(n7996), .QN(n11566)
         );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n2778), .CK(CLK), .Q(n7994), .QN(n11565)
         );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n2777), .CK(CLK), .Q(n7992), .QN(n11564)
         );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n2776), .CK(CLK), .Q(n7990), .QN(n11563)
         );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n2775), .CK(CLK), .Q(n7988), .QN(n11562)
         );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n2774), .CK(CLK), .Q(n7986), .QN(n11561)
         );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n2773), .CK(CLK), .Q(n7984), .QN(n11560)
         );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n2772), .CK(CLK), .Q(n7982), .QN(n11559)
         );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n2771), .CK(CLK), .Q(n7980), .QN(n11558)
         );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n2770), .CK(CLK), .Q(n7978), .QN(n11557)
         );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n2769), .CK(CLK), .Q(n7976), .QN(n11556)
         );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n2768), .CK(CLK), .Q(n7974), .QN(n11555)
         );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n2767), .CK(CLK), .Q(n7972), .QN(n11554)
         );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n2766), .CK(CLK), .Q(n7970), .QN(n11553)
         );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n2765), .CK(CLK), .Q(n7968), .QN(n11552)
         );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n2764), .CK(CLK), .Q(n7966), .QN(n11551)
         );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n2763), .CK(CLK), .Q(n7964), .QN(n11550)
         );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n2762), .CK(CLK), .Q(n9579), .QN(n11888)
         );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n2761), .CK(CLK), .Q(n9578), .QN(n11887)
         );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n2760), .CK(CLK), .Q(n9577), .QN(n11886)
         );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n2759), .CK(CLK), .Q(n9576), .QN(n11885)
         );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n2758), .CK(CLK), .Q(n9575), .QN(n11884)
         );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n2757), .CK(CLK), .Q(n9574), .QN(n11883)
         );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n2756), .CK(CLK), .Q(n9573), .QN(n11882)
         );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n2755), .CK(CLK), .Q(n11468), .QN(n9993)
         );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n2754), .CK(CLK), .Q(n11467), .QN(n9992)
         );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n2753), .CK(CLK), .Q(n11466), .QN(n9991)
         );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n2752), .CK(CLK), .Q(n11465), .QN(n9990)
         );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n2751), .CK(CLK), .Q(n11464), .QN(n9989)
         );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n2750), .CK(CLK), .Q(n8458), .QN(n11881)
         );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n2749), .CK(CLK), .Q(n8456), .QN(n11880)
         );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n2748), .CK(CLK), .Q(n8454), .QN(n11879)
         );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n2747), .CK(CLK), .Q(n8452), .QN(n11799)
         );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n2746), .CK(CLK), .Q(n8450), .QN(n11798)
         );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n2745), .CK(CLK), .Q(n8448), .QN(n11797)
         );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n2744), .CK(CLK), .Q(n8446), .QN(n11796)
         );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n2743), .CK(CLK), .Q(n8444), .QN(n11795)
         );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n2742), .CK(CLK), .Q(n8442), .QN(n11794)
         );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n2741), .CK(CLK), .Q(n8440), .QN(n11793)
         );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n2740), .CK(CLK), .Q(n8438), .QN(n11792)
         );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n2739), .CK(CLK), .Q(n8436), .QN(n11878)
         );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n2738), .CK(CLK), .Q(n11516), .QN(n9935)
         );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n2737), .CK(CLK), .Q(n11512), .QN(n9934)
         );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n2736), .CK(CLK), .Q(n11508), .QN(n9933)
         );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n2735), .CK(CLK), .Q(n11504), .QN(n9932)
         );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n2734), .CK(CLK), .Q(n11500), .QN(n9931)
         );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n2733), .CK(CLK), .Q(n11496), .QN(n9930)
         );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n2732), .CK(CLK), .Q(n11492), .QN(n9929)
         );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n2731), .CK(CLK), .Q(n11488), .QN(n9928)
         );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n4465), .CK(CLK), .QN(n11340) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n4466), .CK(CLK), .QN(n11338) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n4467), .CK(CLK), .QN(n11336) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n4468), .CK(CLK), .QN(n11334) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n4469), .CK(CLK), .QN(n11332) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n4470), .CK(CLK), .QN(n11330) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n4471), .CK(CLK), .QN(n11328) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n4472), .CK(CLK), .QN(n11326) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n4473), .CK(CLK), .QN(n11445) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n4474), .CK(CLK), .QN(n11441) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n4475), .CK(CLK), .QN(n11437) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n4476), .CK(CLK), .QN(n11433) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n4477), .CK(CLK), .QN(n11428) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n4478), .CK(CLK), .QN(n11423) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n4479), .CK(CLK), .QN(n11418) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n4480), .CK(CLK), .QN(n11413) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n4481), .CK(CLK), .QN(n11408) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n4482), .CK(CLK), .QN(n11403) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n4483), .CK(CLK), .QN(n11398) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n4484), .CK(CLK), .QN(n11393) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n4485), .CK(CLK), .QN(n11388) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n4486), .CK(CLK), .QN(n11383) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n4487), .CK(CLK), .QN(n11378) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n4488), .CK(CLK), .QN(n11373) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n4489), .CK(CLK), .QN(n11369) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n4490), .CK(CLK), .QN(n11365) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n4491), .CK(CLK), .QN(n11361) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n4492), .CK(CLK), .QN(n11357) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n4493), .CK(CLK), .QN(n11353) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n4494), .CK(CLK), .QN(n11349) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n4495), .CK(CLK), .QN(n11345) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n4496), .CK(CLK), .QN(n11341) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n4497), .CK(CLK), .QN(n11084) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n4498), .CK(CLK), .QN(n11082) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n4499), .CK(CLK), .QN(n11080) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n4500), .CK(CLK), .QN(n11078) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n4501), .CK(CLK), .QN(n11076) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n4502), .CK(CLK), .QN(n11074) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n4503), .CK(CLK), .QN(n11072) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n4504), .CK(CLK), .QN(n11070) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n4505), .CK(CLK), .QN(n11189) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n4506), .CK(CLK), .QN(n11185) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n4507), .CK(CLK), .QN(n11181) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n4508), .CK(CLK), .QN(n11177) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n4509), .CK(CLK), .QN(n11172) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n4510), .CK(CLK), .QN(n11167) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n4511), .CK(CLK), .QN(n11162) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n4512), .CK(CLK), .QN(n11157) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n4513), .CK(CLK), .QN(n11152) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n4514), .CK(CLK), .QN(n11147) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n4515), .CK(CLK), .QN(n11142) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n4516), .CK(CLK), .QN(n11137) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n4517), .CK(CLK), .QN(n11132) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n4518), .CK(CLK), .QN(n11127) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n4519), .CK(CLK), .QN(n11122) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n4520), .CK(CLK), .QN(n11117) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n4521), .CK(CLK), .QN(n11113) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n4522), .CK(CLK), .QN(n11109) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n4523), .CK(CLK), .QN(n11105) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n4524), .CK(CLK), .QN(n11101) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n4525), .CK(CLK), .QN(n11097) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n4526), .CK(CLK), .QN(n11093) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n4527), .CK(CLK), .QN(n11089) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n4528), .CK(CLK), .QN(n11085) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n2666), .CK(CLK), .Q(n9919), .QN(n11713)
         );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n2665), .CK(CLK), .Q(n9918), .QN(n11712)
         );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n2664), .CK(CLK), .Q(n9917), .QN(n11711)
         );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n2663), .CK(CLK), .Q(n9916), .QN(n11710)
         );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n2662), .CK(CLK), .Q(n9915), .QN(n11709)
         );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n2661), .CK(CLK), .Q(n9914), .QN(n11708)
         );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n2660), .CK(CLK), .Q(n9913), .QN(n11707)
         );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n2659), .CK(CLK), .Q(n7962), .QN(n11706)
         );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n2658), .CK(CLK), .Q(n7960), .QN(n11705)
         );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n2657), .CK(CLK), .Q(n7958), .QN(n11704)
         );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n2656), .CK(CLK), .Q(n7956), .QN(n11549)
         );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n2655), .CK(CLK), .Q(n7954), .QN(n11548)
         );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n2654), .CK(CLK), .Q(n7952), .QN(n11547)
         );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n2653), .CK(CLK), .Q(n7950), .QN(n11546)
         );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n2652), .CK(CLK), .Q(n7948), .QN(n11545)
         );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n2651), .CK(CLK), .Q(n7946), .QN(n11544)
         );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n2650), .CK(CLK), .Q(n7944), .QN(n11543)
         );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n2649), .CK(CLK), .Q(n7942), .QN(n11542)
         );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n2648), .CK(CLK), .Q(n7940), .QN(n11541)
         );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n2647), .CK(CLK), .Q(n7938), .QN(n11540)
         );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n2646), .CK(CLK), .Q(n7936), .QN(n11539)
         );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n2645), .CK(CLK), .Q(n7934), .QN(n11538)
         );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n2644), .CK(CLK), .Q(n7932), .QN(n11537)
         );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n2643), .CK(CLK), .Q(n7930), .QN(n11536)
         );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n2642), .CK(CLK), .Q(n7928), .QN(n11535)
         );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n2641), .CK(CLK), .Q(n7926), .QN(n11534)
         );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n2640), .CK(CLK), .Q(n7924), .QN(n11533)
         );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n2639), .CK(CLK), .Q(n7922), .QN(n11532)
         );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n2638), .CK(CLK), .Q(n7920), .QN(n11531)
         );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n2637), .CK(CLK), .Q(n7918), .QN(n11530)
         );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n2636), .CK(CLK), .Q(n7916), .QN(n11529)
         );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n2635), .CK(CLK), .Q(n7914), .QN(n11528)
         );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n2634), .CK(CLK), .Q(n9607), .QN(n11877)
         );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n2633), .CK(CLK), .Q(n9606), .QN(n11876)
         );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n2632), .CK(CLK), .Q(n9605), .QN(n11875)
         );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n2631), .CK(CLK), .Q(n9604), .QN(n11874)
         );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n2630), .CK(CLK), .Q(n9603), .QN(n11873)
         );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n2629), .CK(CLK), .Q(n9602), .QN(n11872)
         );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n2628), .CK(CLK), .Q(n9601), .QN(n11871)
         );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n2627), .CK(CLK), .Q(n11486), .QN(n9988)
         );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n2626), .CK(CLK), .Q(n11527), .QN(n9987)
         );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n2625), .CK(CLK), .Q(n11525), .QN(n9986)
         );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n2624), .CK(CLK), .Q(n11523), .QN(n9985)
         );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n2623), .CK(CLK), .Q(n11520), .QN(n9984)
         );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n2622), .CK(CLK), .Q(n8408), .QN(n11870)
         );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n2621), .CK(CLK), .Q(n8406), .QN(n11869)
         );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n2620), .CK(CLK), .Q(n8404), .QN(n11868)
         );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n2619), .CK(CLK), .Q(n8402), .QN(n11791)
         );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n2618), .CK(CLK), .Q(n8400), .QN(n11790)
         );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n2617), .CK(CLK), .Q(n8398), .QN(n11789)
         );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n2616), .CK(CLK), .Q(n8396), .QN(n11788)
         );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n2615), .CK(CLK), .Q(n8394), .QN(n11787)
         );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n2614), .CK(CLK), .Q(n8392), .QN(n11786)
         );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n2613), .CK(CLK), .Q(n8390), .QN(n11785)
         );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n2612), .CK(CLK), .Q(n8388), .QN(n11784)
         );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n2611), .CK(CLK), .Q(n8386), .QN(n11867)
         );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n2610), .CK(CLK), .Q(n11515), .QN(n9927)
         );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n2609), .CK(CLK), .Q(n11511), .QN(n9926)
         );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n2608), .CK(CLK), .Q(n11507), .QN(n9925)
         );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n2607), .CK(CLK), .Q(n11503), .QN(n9924)
         );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n2606), .CK(CLK), .Q(n11499), .QN(n9923)
         );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n2605), .CK(CLK), .Q(n11495), .QN(n9922)
         );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n2604), .CK(CLK), .Q(n11491), .QN(n9921)
         );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n2603), .CK(CLK), .Q(n11487), .QN(n9920)
         );
  DFF_X1 \OUT1_reg[31]  ( .D(n2602), .CK(CLK), .Q(OUT1[31]), .QN(n4203) );
  DFF_X1 \OUT1_reg[30]  ( .D(n2601), .CK(CLK), .Q(OUT1[30]), .QN(n4202) );
  DFF_X1 \OUT1_reg[29]  ( .D(n2600), .CK(CLK), .Q(OUT1[29]), .QN(n4201) );
  DFF_X1 \OUT1_reg[28]  ( .D(n2599), .CK(CLK), .Q(OUT1[28]), .QN(n4200) );
  DFF_X1 \OUT1_reg[27]  ( .D(n2598), .CK(CLK), .Q(OUT1[27]), .QN(n4199) );
  DFF_X1 \OUT1_reg[26]  ( .D(n2597), .CK(CLK), .Q(OUT1[26]), .QN(n4198) );
  DFF_X1 \OUT1_reg[25]  ( .D(n2596), .CK(CLK), .Q(OUT1[25]), .QN(n4197) );
  DFF_X1 \OUT1_reg[24]  ( .D(n2595), .CK(CLK), .Q(OUT1[24]), .QN(n4196) );
  DFF_X1 \OUT1_reg[23]  ( .D(n2594), .CK(CLK), .Q(OUT1[23]), .QN(n4195) );
  DFF_X1 \OUT1_reg[22]  ( .D(n2593), .CK(CLK), .Q(OUT1[22]), .QN(n4194) );
  DFF_X1 \OUT1_reg[21]  ( .D(n2592), .CK(CLK), .Q(OUT1[21]), .QN(n4193) );
  DFF_X1 \OUT1_reg[20]  ( .D(n2591), .CK(CLK), .Q(OUT1[20]), .QN(n4192) );
  DFF_X1 \OUT1_reg[19]  ( .D(n2590), .CK(CLK), .Q(OUT1[19]), .QN(n4191) );
  DFF_X1 \OUT1_reg[18]  ( .D(n2589), .CK(CLK), .Q(OUT1[18]), .QN(n4190) );
  DFF_X1 \OUT1_reg[17]  ( .D(n2588), .CK(CLK), .Q(OUT1[17]), .QN(n4189) );
  DFF_X1 \OUT1_reg[16]  ( .D(n2587), .CK(CLK), .Q(OUT1[16]), .QN(n4188) );
  DFF_X1 \OUT1_reg[15]  ( .D(n2586), .CK(CLK), .Q(OUT1[15]), .QN(n4187) );
  DFF_X1 \OUT1_reg[14]  ( .D(n2585), .CK(CLK), .Q(OUT1[14]), .QN(n4186) );
  DFF_X1 \OUT1_reg[13]  ( .D(n2584), .CK(CLK), .Q(OUT1[13]), .QN(n4185) );
  DFF_X1 \OUT1_reg[12]  ( .D(n2583), .CK(CLK), .Q(OUT1[12]), .QN(n4184) );
  DFF_X1 \OUT1_reg[11]  ( .D(n2582), .CK(CLK), .Q(OUT1[11]), .QN(n4183) );
  DFF_X1 \OUT1_reg[10]  ( .D(n2581), .CK(CLK), .Q(OUT1[10]), .QN(n4182) );
  DFF_X1 \OUT1_reg[9]  ( .D(n2580), .CK(CLK), .Q(OUT1[9]), .QN(n4181) );
  DFF_X1 \OUT1_reg[8]  ( .D(n2579), .CK(CLK), .Q(OUT1[8]), .QN(n4180) );
  DFF_X1 \OUT1_reg[7]  ( .D(n2578), .CK(CLK), .Q(OUT1[7]), .QN(n4179) );
  DFF_X1 \OUT1_reg[6]  ( .D(n2577), .CK(CLK), .Q(OUT1[6]), .QN(n4178) );
  DFF_X1 \OUT1_reg[5]  ( .D(n2576), .CK(CLK), .Q(OUT1[5]), .QN(n4177) );
  DFF_X1 \OUT1_reg[4]  ( .D(n2575), .CK(CLK), .Q(OUT1[4]), .QN(n4176) );
  DFF_X1 \OUT1_reg[3]  ( .D(n2574), .CK(CLK), .Q(OUT1[3]), .QN(n4175) );
  DFF_X1 \OUT1_reg[2]  ( .D(n2573), .CK(CLK), .Q(OUT1[2]), .QN(n4174) );
  DFF_X1 \OUT1_reg[1]  ( .D(n2572), .CK(CLK), .Q(OUT1[1]), .QN(n4173) );
  DFF_X1 \OUT1_reg[0]  ( .D(n2571), .CK(CLK), .Q(OUT1[0]), .QN(n4172) );
  DFF_X1 \OUT2_reg[31]  ( .D(n2570), .CK(CLK), .Q(OUT2[31]), .QN(n4171) );
  DFF_X1 \OUT2_reg[30]  ( .D(n2569), .CK(CLK), .Q(OUT2[30]), .QN(n4170) );
  DFF_X1 \OUT2_reg[29]  ( .D(n2568), .CK(CLK), .Q(OUT2[29]), .QN(n4169) );
  DFF_X1 \OUT2_reg[28]  ( .D(n2567), .CK(CLK), .Q(OUT2[28]), .QN(n4168) );
  DFF_X1 \OUT2_reg[27]  ( .D(n2566), .CK(CLK), .Q(OUT2[27]), .QN(n4167) );
  DFF_X1 \OUT2_reg[26]  ( .D(n2565), .CK(CLK), .Q(OUT2[26]), .QN(n4166) );
  DFF_X1 \OUT2_reg[25]  ( .D(n2564), .CK(CLK), .Q(OUT2[25]), .QN(n4165) );
  DFF_X1 \OUT2_reg[24]  ( .D(n2563), .CK(CLK), .Q(OUT2[24]), .QN(n4164) );
  DFF_X1 \OUT2_reg[23]  ( .D(n2562), .CK(CLK), .Q(OUT2[23]), .QN(n4163) );
  DFF_X1 \OUT2_reg[22]  ( .D(n2561), .CK(CLK), .Q(OUT2[22]), .QN(n4162) );
  DFF_X1 \OUT2_reg[21]  ( .D(n2560), .CK(CLK), .Q(OUT2[21]), .QN(n4161) );
  DFF_X1 \OUT2_reg[20]  ( .D(n2559), .CK(CLK), .Q(OUT2[20]), .QN(n4160) );
  DFF_X1 \OUT2_reg[19]  ( .D(n2558), .CK(CLK), .Q(OUT2[19]), .QN(n4159) );
  DFF_X1 \OUT2_reg[18]  ( .D(n2557), .CK(CLK), .Q(OUT2[18]), .QN(n4158) );
  DFF_X1 \OUT2_reg[17]  ( .D(n2556), .CK(CLK), .Q(OUT2[17]), .QN(n4157) );
  DFF_X1 \OUT2_reg[16]  ( .D(n2555), .CK(CLK), .Q(OUT2[16]), .QN(n4156) );
  DFF_X1 \OUT2_reg[15]  ( .D(n2554), .CK(CLK), .Q(OUT2[15]), .QN(n4155) );
  DFF_X1 \OUT2_reg[14]  ( .D(n2553), .CK(CLK), .Q(OUT2[14]), .QN(n4154) );
  DFF_X1 \OUT2_reg[13]  ( .D(n2552), .CK(CLK), .Q(OUT2[13]), .QN(n4153) );
  DFF_X1 \OUT2_reg[12]  ( .D(n2551), .CK(CLK), .Q(OUT2[12]), .QN(n4152) );
  DFF_X1 \OUT2_reg[11]  ( .D(n2550), .CK(CLK), .Q(OUT2[11]), .QN(n4151) );
  DFF_X1 \OUT2_reg[10]  ( .D(n2549), .CK(CLK), .Q(OUT2[10]), .QN(n4150) );
  DFF_X1 \OUT2_reg[9]  ( .D(n2548), .CK(CLK), .Q(OUT2[9]), .QN(n4149) );
  DFF_X1 \OUT2_reg[8]  ( .D(n2547), .CK(CLK), .Q(OUT2[8]), .QN(n4148) );
  DFF_X1 \OUT2_reg[7]  ( .D(n2546), .CK(CLK), .Q(OUT2[7]), .QN(n4147) );
  DFF_X1 \OUT2_reg[6]  ( .D(n2545), .CK(CLK), .Q(OUT2[6]), .QN(n4146) );
  DFF_X1 \OUT2_reg[5]  ( .D(n2544), .CK(CLK), .Q(OUT2[5]), .QN(n4145) );
  DFF_X1 \OUT2_reg[4]  ( .D(n2543), .CK(CLK), .Q(OUT2[4]), .QN(n4144) );
  DFF_X1 \OUT2_reg[3]  ( .D(n2542), .CK(CLK), .Q(OUT2[3]), .QN(n4143) );
  DFF_X1 \OUT2_reg[2]  ( .D(n2541), .CK(CLK), .Q(OUT2[2]), .QN(n4142) );
  DFF_X1 \OUT2_reg[1]  ( .D(n2540), .CK(CLK), .Q(OUT2[1]), .QN(n4141) );
  DFF_X1 \OUT2_reg[0]  ( .D(n2539), .CK(CLK), .Q(OUT2[0]), .QN(n4140) );
  NAND3_X1 U3555 ( .A1(n12563), .A2(n12565), .A3(n12564), .ZN(n1111) );
  NAND3_X1 U3556 ( .A1(n12563), .A2(n12565), .A3(ADD_WR[0]), .ZN(n1109) );
  NAND3_X1 U3557 ( .A1(n12564), .A2(n12563), .A3(ADD_WR[2]), .ZN(n1107) );
  NAND3_X1 U3558 ( .A1(ADD_WR[0]), .A2(n12563), .A3(ADD_WR[2]), .ZN(n1104) );
  NAND3_X1 U3559 ( .A1(n12564), .A2(n12565), .A3(ADD_WR[1]), .ZN(n1120) );
  NAND3_X1 U3560 ( .A1(ADD_WR[0]), .A2(n12565), .A3(ADD_WR[1]), .ZN(n1118) );
  NAND3_X1 U3561 ( .A1(ADD_WR[2]), .A2(n12564), .A3(ADD_WR[1]), .ZN(n1116) );
  NAND3_X1 U3562 ( .A1(ADD_WR[2]), .A2(ADD_WR[0]), .A3(ADD_WR[1]), .ZN(n1114)
         );
  NOR2_X1 U3 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n2448) );
  NOR2_X1 U4 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n1785) );
  BUF_X1 U5 ( .A(n1820), .Z(n12053) );
  BUF_X1 U6 ( .A(n1825), .Z(n12041) );
  BUF_X1 U7 ( .A(n1830), .Z(n12029) );
  BUF_X1 U8 ( .A(n1835), .Z(n12017) );
  BUF_X1 U9 ( .A(n1844), .Z(n12005) );
  BUF_X1 U10 ( .A(n1849), .Z(n11993) );
  BUF_X1 U11 ( .A(n1854), .Z(n11981) );
  BUF_X1 U12 ( .A(n1859), .Z(n11969) );
  BUF_X1 U13 ( .A(n1820), .Z(n12054) );
  BUF_X1 U14 ( .A(n1825), .Z(n12042) );
  BUF_X1 U15 ( .A(n1830), .Z(n12030) );
  BUF_X1 U16 ( .A(n1835), .Z(n12018) );
  BUF_X1 U17 ( .A(n1844), .Z(n12006) );
  BUF_X1 U18 ( .A(n1849), .Z(n11994) );
  BUF_X1 U19 ( .A(n1854), .Z(n11982) );
  BUF_X1 U20 ( .A(n1859), .Z(n11970) );
  BUF_X1 U21 ( .A(n1821), .Z(n12050) );
  BUF_X1 U22 ( .A(n1826), .Z(n12038) );
  BUF_X1 U23 ( .A(n1831), .Z(n12026) );
  BUF_X1 U24 ( .A(n1836), .Z(n12014) );
  BUF_X1 U25 ( .A(n1845), .Z(n12002) );
  BUF_X1 U26 ( .A(n1850), .Z(n11990) );
  BUF_X1 U27 ( .A(n1855), .Z(n11978) );
  BUF_X1 U28 ( .A(n1860), .Z(n11966) );
  BUF_X1 U29 ( .A(n1821), .Z(n12051) );
  BUF_X1 U30 ( .A(n1826), .Z(n12039) );
  BUF_X1 U31 ( .A(n1831), .Z(n12027) );
  BUF_X1 U32 ( .A(n1836), .Z(n12015) );
  BUF_X1 U33 ( .A(n1845), .Z(n12003) );
  BUF_X1 U34 ( .A(n1850), .Z(n11991) );
  BUF_X1 U35 ( .A(n1855), .Z(n11979) );
  BUF_X1 U36 ( .A(n1860), .Z(n11967) );
  BUF_X1 U37 ( .A(n1820), .Z(n12055) );
  BUF_X1 U38 ( .A(n1825), .Z(n12043) );
  BUF_X1 U39 ( .A(n1830), .Z(n12031) );
  BUF_X1 U40 ( .A(n1835), .Z(n12019) );
  BUF_X1 U41 ( .A(n1844), .Z(n12007) );
  BUF_X1 U42 ( .A(n1849), .Z(n11995) );
  BUF_X1 U43 ( .A(n1854), .Z(n11983) );
  BUF_X1 U44 ( .A(n1859), .Z(n11971) );
  BUF_X1 U45 ( .A(n1821), .Z(n12052) );
  BUF_X1 U46 ( .A(n1826), .Z(n12040) );
  BUF_X1 U47 ( .A(n1831), .Z(n12028) );
  BUF_X1 U48 ( .A(n1836), .Z(n12016) );
  BUF_X1 U49 ( .A(n1845), .Z(n12004) );
  BUF_X1 U50 ( .A(n1850), .Z(n11992) );
  BUF_X1 U51 ( .A(n1855), .Z(n11980) );
  BUF_X1 U52 ( .A(n1860), .Z(n11968) );
  BUF_X1 U53 ( .A(n1828), .Z(n12035) );
  BUF_X1 U54 ( .A(n1838), .Z(n12011) );
  BUF_X1 U55 ( .A(n1852), .Z(n11987) );
  BUF_X1 U56 ( .A(n1828), .Z(n12036) );
  BUF_X1 U57 ( .A(n1838), .Z(n12012) );
  BUF_X1 U58 ( .A(n1852), .Z(n11988) );
  BUF_X1 U59 ( .A(n1862), .Z(n11963) );
  BUF_X1 U60 ( .A(n1862), .Z(n11964) );
  BUF_X1 U61 ( .A(n1823), .Z(n12047) );
  BUF_X1 U62 ( .A(n1833), .Z(n12023) );
  BUF_X1 U63 ( .A(n1847), .Z(n11999) );
  BUF_X1 U64 ( .A(n1857), .Z(n11975) );
  BUF_X1 U65 ( .A(n1823), .Z(n12048) );
  BUF_X1 U66 ( .A(n1833), .Z(n12024) );
  BUF_X1 U67 ( .A(n1847), .Z(n12000) );
  BUF_X1 U68 ( .A(n1857), .Z(n11976) );
  BUF_X1 U69 ( .A(n1829), .Z(n12032) );
  BUF_X1 U70 ( .A(n1839), .Z(n12008) );
  BUF_X1 U71 ( .A(n1848), .Z(n11996) );
  BUF_X1 U72 ( .A(n1853), .Z(n11984) );
  BUF_X1 U73 ( .A(n1829), .Z(n12033) );
  BUF_X1 U74 ( .A(n1839), .Z(n12009) );
  BUF_X1 U75 ( .A(n1848), .Z(n11997) );
  BUF_X1 U76 ( .A(n1853), .Z(n11985) );
  BUF_X1 U77 ( .A(n1863), .Z(n11960) );
  BUF_X1 U78 ( .A(n1863), .Z(n11961) );
  BUF_X1 U79 ( .A(n1824), .Z(n12044) );
  BUF_X1 U80 ( .A(n1834), .Z(n12020) );
  BUF_X1 U81 ( .A(n1858), .Z(n11972) );
  BUF_X1 U82 ( .A(n1824), .Z(n12045) );
  BUF_X1 U83 ( .A(n1834), .Z(n12021) );
  BUF_X1 U84 ( .A(n1858), .Z(n11973) );
  BUF_X1 U85 ( .A(n1828), .Z(n12037) );
  BUF_X1 U86 ( .A(n1838), .Z(n12013) );
  BUF_X1 U87 ( .A(n1852), .Z(n11989) );
  BUF_X1 U88 ( .A(n1862), .Z(n11965) );
  BUF_X1 U89 ( .A(n1823), .Z(n12049) );
  BUF_X1 U90 ( .A(n1833), .Z(n12025) );
  BUF_X1 U91 ( .A(n1847), .Z(n12001) );
  BUF_X1 U92 ( .A(n1857), .Z(n11977) );
  BUF_X1 U93 ( .A(n1829), .Z(n12034) );
  BUF_X1 U94 ( .A(n1839), .Z(n12010) );
  BUF_X1 U95 ( .A(n1848), .Z(n11998) );
  BUF_X1 U96 ( .A(n1853), .Z(n11986) );
  BUF_X1 U97 ( .A(n1863), .Z(n11962) );
  BUF_X1 U98 ( .A(n1824), .Z(n12046) );
  BUF_X1 U99 ( .A(n1834), .Z(n12022) );
  BUF_X1 U100 ( .A(n1858), .Z(n11974) );
  INV_X1 U101 ( .A(n12213), .ZN(n12206) );
  INV_X1 U102 ( .A(n12249), .ZN(n12242) );
  INV_X1 U103 ( .A(n12285), .ZN(n12278) );
  INV_X1 U104 ( .A(n12321), .ZN(n12314) );
  INV_X1 U105 ( .A(n12366), .ZN(n12359) );
  INV_X1 U106 ( .A(n12384), .ZN(n12377) );
  INV_X1 U107 ( .A(n12186), .ZN(n12179) );
  INV_X1 U108 ( .A(n12549), .ZN(n12542) );
  INV_X1 U109 ( .A(n12447), .ZN(n12440) );
  INV_X1 U110 ( .A(n12204), .ZN(n12197) );
  INV_X1 U111 ( .A(n12438), .ZN(n12431) );
  INV_X1 U112 ( .A(n12429), .ZN(n12422) );
  INV_X1 U113 ( .A(n12222), .ZN(n12215) );
  INV_X1 U114 ( .A(n12231), .ZN(n12224) );
  INV_X1 U115 ( .A(n12240), .ZN(n12233) );
  INV_X1 U116 ( .A(n12258), .ZN(n12251) );
  INV_X1 U117 ( .A(n12267), .ZN(n12260) );
  INV_X1 U118 ( .A(n12276), .ZN(n12269) );
  INV_X1 U119 ( .A(n12294), .ZN(n12287) );
  INV_X1 U120 ( .A(n12303), .ZN(n12296) );
  INV_X1 U121 ( .A(n12312), .ZN(n12305) );
  INV_X1 U122 ( .A(n12330), .ZN(n12323) );
  INV_X1 U123 ( .A(n12339), .ZN(n12332) );
  INV_X1 U124 ( .A(n12348), .ZN(n12341) );
  INV_X1 U125 ( .A(n12420), .ZN(n12413) );
  INV_X1 U126 ( .A(n12411), .ZN(n12404) );
  INV_X1 U127 ( .A(n12357), .ZN(n12350) );
  INV_X1 U128 ( .A(n12402), .ZN(n12395) );
  INV_X1 U129 ( .A(n12393), .ZN(n12386) );
  INV_X1 U130 ( .A(n12375), .ZN(n12368) );
  NAND2_X1 U131 ( .A1(n2448), .A2(n2459), .ZN(n1853) );
  NAND2_X1 U132 ( .A1(n2448), .A2(n2460), .ZN(n1852) );
  NAND2_X1 U133 ( .A1(n2460), .A2(n2444), .ZN(n1847) );
  NAND2_X1 U134 ( .A1(n2463), .A2(n2446), .ZN(n1858) );
  NAND2_X1 U135 ( .A1(n2464), .A2(n2446), .ZN(n1857) );
  NAND2_X1 U136 ( .A1(n2463), .A2(n2449), .ZN(n1863) );
  NAND2_X1 U137 ( .A1(n2464), .A2(n2449), .ZN(n1862) );
  NAND2_X1 U138 ( .A1(n2443), .A2(n2448), .ZN(n1829) );
  NAND2_X1 U139 ( .A1(n2445), .A2(n2448), .ZN(n1828) );
  NAND2_X1 U140 ( .A1(n2451), .A2(n2448), .ZN(n1839) );
  NAND2_X1 U141 ( .A1(n2452), .A2(n2448), .ZN(n1838) );
  NAND2_X1 U142 ( .A1(n2444), .A2(n2459), .ZN(n1848) );
  NAND2_X1 U143 ( .A1(n2443), .A2(n2444), .ZN(n1824) );
  NAND2_X1 U144 ( .A1(n2445), .A2(n2444), .ZN(n1823) );
  NAND2_X1 U145 ( .A1(n2451), .A2(n2444), .ZN(n1834) );
  NAND2_X1 U146 ( .A1(n2452), .A2(n2444), .ZN(n1833) );
  AND2_X1 U147 ( .A1(n2449), .A2(n2460), .ZN(n1849) );
  AND2_X1 U148 ( .A1(n2449), .A2(n2459), .ZN(n1850) );
  AND2_X1 U149 ( .A1(n2464), .A2(n2444), .ZN(n1854) );
  AND2_X1 U150 ( .A1(n2463), .A2(n2444), .ZN(n1855) );
  AND2_X1 U151 ( .A1(n2464), .A2(n2448), .ZN(n1859) );
  AND2_X1 U152 ( .A1(n2463), .A2(n2448), .ZN(n1860) );
  AND2_X1 U153 ( .A1(n2443), .A2(n2449), .ZN(n1826) );
  AND2_X1 U154 ( .A1(n2445), .A2(n2449), .ZN(n1825) );
  AND2_X1 U155 ( .A1(n2452), .A2(n2449), .ZN(n1835) );
  AND2_X1 U156 ( .A1(n2451), .A2(n2449), .ZN(n1836) );
  AND2_X1 U157 ( .A1(n2446), .A2(n2459), .ZN(n1845) );
  AND2_X1 U158 ( .A1(n2446), .A2(n2460), .ZN(n1844) );
  AND2_X1 U159 ( .A1(n2443), .A2(n2446), .ZN(n1821) );
  AND2_X1 U160 ( .A1(n2445), .A2(n2446), .ZN(n1820) );
  AND2_X1 U161 ( .A1(n2452), .A2(n2446), .ZN(n1830) );
  AND2_X1 U162 ( .A1(n2451), .A2(n2446), .ZN(n1831) );
  NOR2_X1 U163 ( .A1(n12569), .A2(ADD_RD2[2]), .ZN(n2449) );
  NOR3_X1 U164 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n12570), .ZN(n2459) );
  NOR3_X1 U165 ( .A1(n12568), .A2(ADD_RD2[4]), .A3(n12570), .ZN(n2460) );
  NOR3_X1 U166 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(n2464)
         );
  NOR3_X1 U167 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n12568), .ZN(n2463) );
  AND2_X1 U168 ( .A1(ADD_RD2[2]), .A2(n12569), .ZN(n2444) );
  BUF_X1 U169 ( .A(n1815), .Z(n12056) );
  BUF_X1 U170 ( .A(n1815), .Z(n12057) );
  BUF_X1 U171 ( .A(n1810), .Z(n12062) );
  BUF_X1 U172 ( .A(n1085), .Z(n12505) );
  BUF_X1 U173 ( .A(n1086), .Z(n12502) );
  BUF_X1 U174 ( .A(n1087), .Z(n12499) );
  BUF_X1 U175 ( .A(n1099), .Z(n12463) );
  BUF_X1 U176 ( .A(n1100), .Z(n12460) );
  BUF_X1 U177 ( .A(n1103), .Z(n12451) );
  BUF_X1 U178 ( .A(n1815), .Z(n12058) );
  BUF_X1 U179 ( .A(n1810), .Z(n12064) );
  BUF_X1 U180 ( .A(n1085), .Z(n12503) );
  BUF_X1 U181 ( .A(n1086), .Z(n12500) );
  BUF_X1 U182 ( .A(n1087), .Z(n12497) );
  BUF_X1 U183 ( .A(n1099), .Z(n12461) );
  BUF_X1 U184 ( .A(n1100), .Z(n12458) );
  BUF_X1 U185 ( .A(n1103), .Z(n12449) );
  BUF_X1 U186 ( .A(n1086), .Z(n12501) );
  BUF_X1 U187 ( .A(n1087), .Z(n12498) );
  BUF_X1 U188 ( .A(n1099), .Z(n12462) );
  BUF_X1 U189 ( .A(n1100), .Z(n12459) );
  BUF_X1 U190 ( .A(n1103), .Z(n12450) );
  AND2_X1 U191 ( .A1(ADD_RD2[2]), .A2(ADD_RD2[1]), .ZN(n2446) );
  BUF_X1 U192 ( .A(n1810), .Z(n12063) );
  AND3_X1 U193 ( .A1(ADD_RD2[4]), .A2(n12568), .A3(ADD_RD2[3]), .ZN(n2443) );
  AND3_X1 U194 ( .A1(ADD_RD2[4]), .A2(n12570), .A3(ADD_RD2[0]), .ZN(n2452) );
  AND3_X1 U195 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(ADD_RD2[3]), .ZN(n2445)
         );
  AND3_X1 U196 ( .A1(n12568), .A2(n12570), .A3(ADD_RD2[4]), .ZN(n2451) );
  INV_X1 U197 ( .A(ADD_RD2[3]), .ZN(n12570) );
  INV_X1 U198 ( .A(ADD_RD2[0]), .ZN(n12568) );
  BUF_X1 U199 ( .A(n12187), .Z(n12186) );
  BUF_X1 U200 ( .A(n12205), .Z(n12204) );
  BUF_X1 U201 ( .A(n12223), .Z(n12222) );
  BUF_X1 U202 ( .A(n12232), .Z(n12231) );
  BUF_X1 U203 ( .A(n12241), .Z(n12240) );
  BUF_X1 U204 ( .A(n12259), .Z(n12258) );
  BUF_X1 U205 ( .A(n12268), .Z(n12267) );
  BUF_X1 U206 ( .A(n12277), .Z(n12276) );
  BUF_X1 U207 ( .A(n12295), .Z(n12294) );
  BUF_X1 U208 ( .A(n12304), .Z(n12303) );
  BUF_X1 U209 ( .A(n12313), .Z(n12312) );
  BUF_X1 U210 ( .A(n12331), .Z(n12330) );
  BUF_X1 U211 ( .A(n12340), .Z(n12339) );
  BUF_X1 U212 ( .A(n12349), .Z(n12348) );
  BUF_X1 U213 ( .A(n12421), .Z(n12420) );
  BUF_X1 U214 ( .A(n12412), .Z(n12411) );
  BUF_X1 U215 ( .A(n12358), .Z(n12357) );
  BUF_X1 U216 ( .A(n12403), .Z(n12402) );
  BUF_X1 U217 ( .A(n12394), .Z(n12393) );
  BUF_X1 U218 ( .A(n12376), .Z(n12375) );
  BUF_X1 U219 ( .A(n12550), .Z(n12549) );
  BUF_X1 U220 ( .A(n12448), .Z(n12447) );
  BUF_X1 U221 ( .A(n12439), .Z(n12438) );
  BUF_X1 U222 ( .A(n12430), .Z(n12429) );
  BUF_X1 U223 ( .A(n12178), .Z(n12177) );
  BUF_X1 U224 ( .A(n12196), .Z(n12195) );
  BUF_X1 U225 ( .A(n12214), .Z(n12213) );
  BUF_X1 U226 ( .A(n12250), .Z(n12249) );
  BUF_X1 U227 ( .A(n12286), .Z(n12285) );
  BUF_X1 U228 ( .A(n12322), .Z(n12321) );
  BUF_X1 U229 ( .A(n12367), .Z(n12366) );
  BUF_X1 U230 ( .A(n12385), .Z(n12384) );
  INV_X1 U231 ( .A(ADD_RD2[1]), .ZN(n12569) );
  BUF_X1 U232 ( .A(n1167), .Z(n12134) );
  BUF_X1 U233 ( .A(n1157), .Z(n12158) );
  BUF_X1 U234 ( .A(n1162), .Z(n12146) );
  BUF_X1 U235 ( .A(n1172), .Z(n12122) );
  BUF_X1 U236 ( .A(n1181), .Z(n12110) );
  BUF_X1 U237 ( .A(n1186), .Z(n12098) );
  BUF_X1 U238 ( .A(n1191), .Z(n12086) );
  BUF_X1 U239 ( .A(n1196), .Z(n12074) );
  BUF_X1 U240 ( .A(n1167), .Z(n12135) );
  BUF_X1 U241 ( .A(n1157), .Z(n12159) );
  BUF_X1 U242 ( .A(n1162), .Z(n12147) );
  BUF_X1 U243 ( .A(n1172), .Z(n12123) );
  BUF_X1 U244 ( .A(n1181), .Z(n12111) );
  BUF_X1 U245 ( .A(n1186), .Z(n12099) );
  BUF_X1 U246 ( .A(n1191), .Z(n12087) );
  BUF_X1 U247 ( .A(n1196), .Z(n12075) );
  BUF_X1 U248 ( .A(n1152), .Z(n12161) );
  BUF_X1 U249 ( .A(n1152), .Z(n12162) );
  BUF_X1 U250 ( .A(n1168), .Z(n12131) );
  BUF_X1 U251 ( .A(n1158), .Z(n12155) );
  BUF_X1 U252 ( .A(n1163), .Z(n12143) );
  BUF_X1 U253 ( .A(n1173), .Z(n12119) );
  BUF_X1 U254 ( .A(n1182), .Z(n12107) );
  BUF_X1 U255 ( .A(n1187), .Z(n12095) );
  BUF_X1 U256 ( .A(n1192), .Z(n12083) );
  BUF_X1 U257 ( .A(n1197), .Z(n12071) );
  BUF_X1 U258 ( .A(n1168), .Z(n12132) );
  BUF_X1 U259 ( .A(n1158), .Z(n12156) );
  BUF_X1 U260 ( .A(n1163), .Z(n12144) );
  BUF_X1 U261 ( .A(n1173), .Z(n12120) );
  BUF_X1 U262 ( .A(n1182), .Z(n12108) );
  BUF_X1 U263 ( .A(n1187), .Z(n12096) );
  BUF_X1 U264 ( .A(n1192), .Z(n12084) );
  BUF_X1 U265 ( .A(n1197), .Z(n12072) );
  BUF_X1 U266 ( .A(n1147), .Z(n12167) );
  BUF_X1 U267 ( .A(n1083), .Z(n12511) );
  BUF_X1 U268 ( .A(n1084), .Z(n12508) );
  BUF_X1 U269 ( .A(n1088), .Z(n12496) );
  BUF_X1 U270 ( .A(n1090), .Z(n12490) );
  BUF_X1 U271 ( .A(n1091), .Z(n12487) );
  BUF_X1 U272 ( .A(n1093), .Z(n12481) );
  BUF_X1 U273 ( .A(n1094), .Z(n12478) );
  BUF_X1 U274 ( .A(n1074), .Z(n12538) );
  BUF_X1 U275 ( .A(n1076), .Z(n12532) );
  BUF_X1 U276 ( .A(n1077), .Z(n12529) );
  BUF_X1 U277 ( .A(n1078), .Z(n12526) );
  BUF_X1 U278 ( .A(n1079), .Z(n12523) );
  BUF_X1 U279 ( .A(n1080), .Z(n12520) );
  BUF_X1 U280 ( .A(n1181), .Z(n12112) );
  BUF_X1 U281 ( .A(n1186), .Z(n12100) );
  BUF_X1 U282 ( .A(n1191), .Z(n12088) );
  BUF_X1 U283 ( .A(n1196), .Z(n12076) );
  BUF_X1 U284 ( .A(n1167), .Z(n12136) );
  BUF_X1 U285 ( .A(n1157), .Z(n12160) );
  BUF_X1 U286 ( .A(n1162), .Z(n12148) );
  BUF_X1 U287 ( .A(n1172), .Z(n12124) );
  BUF_X1 U288 ( .A(n1152), .Z(n12163) );
  BUF_X1 U289 ( .A(n1182), .Z(n12109) );
  BUF_X1 U290 ( .A(n1187), .Z(n12097) );
  BUF_X1 U291 ( .A(n1192), .Z(n12085) );
  BUF_X1 U292 ( .A(n1197), .Z(n12073) );
  BUF_X1 U293 ( .A(n1168), .Z(n12133) );
  BUF_X1 U294 ( .A(n1158), .Z(n12157) );
  BUF_X1 U295 ( .A(n1163), .Z(n12145) );
  BUF_X1 U296 ( .A(n1173), .Z(n12121) );
  BUF_X1 U297 ( .A(n1147), .Z(n12169) );
  BUF_X1 U298 ( .A(n1083), .Z(n12509) );
  BUF_X1 U299 ( .A(n1084), .Z(n12506) );
  BUF_X1 U300 ( .A(n1088), .Z(n12494) );
  BUF_X1 U301 ( .A(n1090), .Z(n12488) );
  BUF_X1 U302 ( .A(n1091), .Z(n12485) );
  BUF_X1 U303 ( .A(n1093), .Z(n12479) );
  BUF_X1 U304 ( .A(n1094), .Z(n12476) );
  BUF_X1 U305 ( .A(n1074), .Z(n12536) );
  BUF_X1 U306 ( .A(n1076), .Z(n12530) );
  BUF_X1 U307 ( .A(n1077), .Z(n12527) );
  BUF_X1 U308 ( .A(n1078), .Z(n12524) );
  BUF_X1 U309 ( .A(n1079), .Z(n12521) );
  BUF_X1 U310 ( .A(n1080), .Z(n12518) );
  BUF_X1 U311 ( .A(n1083), .Z(n12510) );
  BUF_X1 U312 ( .A(n1084), .Z(n12507) );
  BUF_X1 U313 ( .A(n1085), .Z(n12504) );
  BUF_X1 U314 ( .A(n1088), .Z(n12495) );
  BUF_X1 U315 ( .A(n1090), .Z(n12489) );
  BUF_X1 U316 ( .A(n1091), .Z(n12486) );
  BUF_X1 U317 ( .A(n1093), .Z(n12480) );
  BUF_X1 U318 ( .A(n1094), .Z(n12477) );
  BUF_X1 U319 ( .A(n1074), .Z(n12537) );
  BUF_X1 U320 ( .A(n1076), .Z(n12531) );
  BUF_X1 U321 ( .A(n1077), .Z(n12528) );
  BUF_X1 U322 ( .A(n1078), .Z(n12525) );
  BUF_X1 U323 ( .A(n1079), .Z(n12522) );
  BUF_X1 U324 ( .A(n1080), .Z(n12519) );
  BUF_X1 U325 ( .A(n1165), .Z(n12140) );
  BUF_X1 U326 ( .A(n1175), .Z(n12116) );
  BUF_X1 U327 ( .A(n1165), .Z(n12141) );
  BUF_X1 U328 ( .A(n1175), .Z(n12117) );
  BUF_X1 U329 ( .A(n1189), .Z(n12092) );
  BUF_X1 U330 ( .A(n1199), .Z(n12068) );
  BUF_X1 U331 ( .A(n1189), .Z(n12093) );
  BUF_X1 U332 ( .A(n1199), .Z(n12069) );
  BUF_X1 U333 ( .A(n1184), .Z(n12104) );
  BUF_X1 U334 ( .A(n1194), .Z(n12080) );
  BUF_X1 U335 ( .A(n1184), .Z(n12105) );
  BUF_X1 U336 ( .A(n1194), .Z(n12081) );
  BUF_X1 U337 ( .A(n1170), .Z(n12128) );
  BUF_X1 U338 ( .A(n1160), .Z(n12152) );
  BUF_X1 U339 ( .A(n1170), .Z(n12129) );
  BUF_X1 U340 ( .A(n1160), .Z(n12153) );
  BUF_X1 U341 ( .A(n1166), .Z(n12137) );
  BUF_X1 U342 ( .A(n1176), .Z(n12113) );
  BUF_X1 U343 ( .A(n1166), .Z(n12138) );
  BUF_X1 U344 ( .A(n1176), .Z(n12114) );
  BUF_X1 U345 ( .A(n1185), .Z(n12101) );
  BUF_X1 U346 ( .A(n1190), .Z(n12089) );
  BUF_X1 U347 ( .A(n1185), .Z(n12102) );
  BUF_X1 U348 ( .A(n1190), .Z(n12090) );
  BUF_X1 U349 ( .A(n1200), .Z(n12065) );
  BUF_X1 U350 ( .A(n1200), .Z(n12066) );
  BUF_X1 U351 ( .A(n1195), .Z(n12077) );
  BUF_X1 U352 ( .A(n1195), .Z(n12078) );
  BUF_X1 U353 ( .A(n1171), .Z(n12125) );
  BUF_X1 U354 ( .A(n1161), .Z(n12149) );
  BUF_X1 U355 ( .A(n1171), .Z(n12126) );
  BUF_X1 U356 ( .A(n1161), .Z(n12150) );
  BUF_X1 U357 ( .A(n1165), .Z(n12142) );
  BUF_X1 U358 ( .A(n1175), .Z(n12118) );
  BUF_X1 U359 ( .A(n1189), .Z(n12094) );
  BUF_X1 U360 ( .A(n1199), .Z(n12070) );
  BUF_X1 U361 ( .A(n1184), .Z(n12106) );
  BUF_X1 U362 ( .A(n1194), .Z(n12082) );
  BUF_X1 U363 ( .A(n1170), .Z(n12130) );
  BUF_X1 U364 ( .A(n1160), .Z(n12154) );
  BUF_X1 U365 ( .A(n1166), .Z(n12139) );
  BUF_X1 U366 ( .A(n1176), .Z(n12115) );
  BUF_X1 U367 ( .A(n1185), .Z(n12103) );
  BUF_X1 U368 ( .A(n1190), .Z(n12091) );
  BUF_X1 U369 ( .A(n1200), .Z(n12067) );
  BUF_X1 U370 ( .A(n1195), .Z(n12079) );
  BUF_X1 U371 ( .A(n1171), .Z(n12127) );
  BUF_X1 U372 ( .A(n1161), .Z(n12151) );
  BUF_X1 U373 ( .A(n1147), .Z(n12168) );
  BUF_X1 U374 ( .A(n12178), .Z(n12176) );
  BUF_X1 U375 ( .A(n12178), .Z(n12175) );
  BUF_X1 U376 ( .A(n12178), .Z(n12174) );
  BUF_X1 U377 ( .A(n12178), .Z(n12173) );
  BUF_X1 U378 ( .A(n12178), .Z(n12172) );
  BUF_X1 U379 ( .A(n12178), .Z(n12171) );
  BUF_X1 U380 ( .A(n12187), .Z(n12185) );
  BUF_X1 U381 ( .A(n12187), .Z(n12184) );
  BUF_X1 U382 ( .A(n12187), .Z(n12183) );
  BUF_X1 U383 ( .A(n12187), .Z(n12182) );
  BUF_X1 U384 ( .A(n12187), .Z(n12181) );
  BUF_X1 U385 ( .A(n12187), .Z(n12180) );
  BUF_X1 U386 ( .A(n12196), .Z(n12194) );
  BUF_X1 U387 ( .A(n12196), .Z(n12193) );
  BUF_X1 U388 ( .A(n12196), .Z(n12192) );
  BUF_X1 U389 ( .A(n12196), .Z(n12191) );
  BUF_X1 U390 ( .A(n12196), .Z(n12190) );
  BUF_X1 U391 ( .A(n12196), .Z(n12189) );
  BUF_X1 U392 ( .A(n12205), .Z(n12203) );
  BUF_X1 U393 ( .A(n12205), .Z(n12202) );
  BUF_X1 U394 ( .A(n12205), .Z(n12201) );
  BUF_X1 U395 ( .A(n12205), .Z(n12200) );
  BUF_X1 U396 ( .A(n12205), .Z(n12199) );
  BUF_X1 U397 ( .A(n12205), .Z(n12198) );
  BUF_X1 U398 ( .A(n12214), .Z(n12212) );
  BUF_X1 U399 ( .A(n12214), .Z(n12211) );
  BUF_X1 U400 ( .A(n12214), .Z(n12210) );
  BUF_X1 U401 ( .A(n12214), .Z(n12209) );
  BUF_X1 U402 ( .A(n12214), .Z(n12208) );
  BUF_X1 U403 ( .A(n12214), .Z(n12207) );
  BUF_X1 U404 ( .A(n12223), .Z(n12221) );
  BUF_X1 U405 ( .A(n12223), .Z(n12220) );
  BUF_X1 U406 ( .A(n12223), .Z(n12219) );
  BUF_X1 U407 ( .A(n12223), .Z(n12218) );
  BUF_X1 U408 ( .A(n12223), .Z(n12217) );
  BUF_X1 U409 ( .A(n12223), .Z(n12216) );
  BUF_X1 U410 ( .A(n12232), .Z(n12230) );
  BUF_X1 U411 ( .A(n12232), .Z(n12229) );
  BUF_X1 U412 ( .A(n12232), .Z(n12228) );
  BUF_X1 U413 ( .A(n12232), .Z(n12227) );
  BUF_X1 U414 ( .A(n12232), .Z(n12226) );
  BUF_X1 U415 ( .A(n12232), .Z(n12225) );
  BUF_X1 U416 ( .A(n12241), .Z(n12239) );
  BUF_X1 U417 ( .A(n12241), .Z(n12238) );
  BUF_X1 U418 ( .A(n12241), .Z(n12237) );
  BUF_X1 U419 ( .A(n12241), .Z(n12236) );
  BUF_X1 U420 ( .A(n12241), .Z(n12235) );
  BUF_X1 U421 ( .A(n12241), .Z(n12234) );
  BUF_X1 U422 ( .A(n12250), .Z(n12248) );
  BUF_X1 U423 ( .A(n12250), .Z(n12247) );
  BUF_X1 U424 ( .A(n12250), .Z(n12246) );
  BUF_X1 U425 ( .A(n12250), .Z(n12245) );
  BUF_X1 U426 ( .A(n12250), .Z(n12244) );
  BUF_X1 U427 ( .A(n12250), .Z(n12243) );
  BUF_X1 U428 ( .A(n12259), .Z(n12257) );
  BUF_X1 U429 ( .A(n12259), .Z(n12256) );
  BUF_X1 U430 ( .A(n12259), .Z(n12255) );
  BUF_X1 U431 ( .A(n12259), .Z(n12254) );
  BUF_X1 U432 ( .A(n12259), .Z(n12253) );
  BUF_X1 U433 ( .A(n12259), .Z(n12252) );
  BUF_X1 U434 ( .A(n12268), .Z(n12266) );
  BUF_X1 U435 ( .A(n12268), .Z(n12265) );
  BUF_X1 U436 ( .A(n12268), .Z(n12264) );
  BUF_X1 U437 ( .A(n12268), .Z(n12263) );
  BUF_X1 U438 ( .A(n12268), .Z(n12262) );
  BUF_X1 U439 ( .A(n12268), .Z(n12261) );
  BUF_X1 U440 ( .A(n12277), .Z(n12275) );
  BUF_X1 U441 ( .A(n12277), .Z(n12274) );
  BUF_X1 U442 ( .A(n12277), .Z(n12273) );
  BUF_X1 U443 ( .A(n12277), .Z(n12272) );
  BUF_X1 U444 ( .A(n12277), .Z(n12271) );
  BUF_X1 U445 ( .A(n12277), .Z(n12270) );
  BUF_X1 U446 ( .A(n12286), .Z(n12284) );
  BUF_X1 U447 ( .A(n12286), .Z(n12283) );
  BUF_X1 U448 ( .A(n12286), .Z(n12282) );
  BUF_X1 U449 ( .A(n12286), .Z(n12281) );
  BUF_X1 U450 ( .A(n12286), .Z(n12280) );
  BUF_X1 U451 ( .A(n12286), .Z(n12279) );
  BUF_X1 U452 ( .A(n12295), .Z(n12293) );
  BUF_X1 U453 ( .A(n12295), .Z(n12292) );
  BUF_X1 U454 ( .A(n12295), .Z(n12291) );
  BUF_X1 U455 ( .A(n12295), .Z(n12290) );
  BUF_X1 U456 ( .A(n12295), .Z(n12289) );
  BUF_X1 U457 ( .A(n12295), .Z(n12288) );
  BUF_X1 U458 ( .A(n12304), .Z(n12302) );
  BUF_X1 U459 ( .A(n12304), .Z(n12301) );
  BUF_X1 U460 ( .A(n12304), .Z(n12300) );
  BUF_X1 U461 ( .A(n12304), .Z(n12299) );
  BUF_X1 U462 ( .A(n12304), .Z(n12298) );
  BUF_X1 U463 ( .A(n12304), .Z(n12297) );
  BUF_X1 U464 ( .A(n12313), .Z(n12311) );
  BUF_X1 U465 ( .A(n12313), .Z(n12310) );
  BUF_X1 U466 ( .A(n12313), .Z(n12309) );
  BUF_X1 U467 ( .A(n12313), .Z(n12308) );
  BUF_X1 U468 ( .A(n12313), .Z(n12307) );
  BUF_X1 U469 ( .A(n12313), .Z(n12306) );
  BUF_X1 U470 ( .A(n12322), .Z(n12320) );
  BUF_X1 U471 ( .A(n12322), .Z(n12319) );
  BUF_X1 U472 ( .A(n12322), .Z(n12318) );
  BUF_X1 U473 ( .A(n12322), .Z(n12317) );
  BUF_X1 U474 ( .A(n12322), .Z(n12316) );
  BUF_X1 U475 ( .A(n12322), .Z(n12315) );
  BUF_X1 U476 ( .A(n12331), .Z(n12329) );
  BUF_X1 U477 ( .A(n12331), .Z(n12328) );
  BUF_X1 U478 ( .A(n12331), .Z(n12327) );
  BUF_X1 U479 ( .A(n12331), .Z(n12326) );
  BUF_X1 U480 ( .A(n12331), .Z(n12325) );
  BUF_X1 U481 ( .A(n12331), .Z(n12324) );
  BUF_X1 U482 ( .A(n12340), .Z(n12338) );
  BUF_X1 U483 ( .A(n12340), .Z(n12337) );
  BUF_X1 U484 ( .A(n12340), .Z(n12336) );
  BUF_X1 U485 ( .A(n12340), .Z(n12335) );
  BUF_X1 U486 ( .A(n12340), .Z(n12334) );
  BUF_X1 U487 ( .A(n12340), .Z(n12333) );
  BUF_X1 U488 ( .A(n12349), .Z(n12347) );
  BUF_X1 U489 ( .A(n12349), .Z(n12346) );
  BUF_X1 U490 ( .A(n12349), .Z(n12345) );
  BUF_X1 U491 ( .A(n12349), .Z(n12344) );
  BUF_X1 U492 ( .A(n12349), .Z(n12343) );
  BUF_X1 U493 ( .A(n12349), .Z(n12342) );
  BUF_X1 U494 ( .A(n12421), .Z(n12414) );
  BUF_X1 U495 ( .A(n12421), .Z(n12415) );
  BUF_X1 U496 ( .A(n12421), .Z(n12416) );
  BUF_X1 U497 ( .A(n12421), .Z(n12417) );
  BUF_X1 U498 ( .A(n12421), .Z(n12418) );
  BUF_X1 U499 ( .A(n12421), .Z(n12419) );
  BUF_X1 U500 ( .A(n12412), .Z(n12405) );
  BUF_X1 U501 ( .A(n12412), .Z(n12406) );
  BUF_X1 U502 ( .A(n12412), .Z(n12407) );
  BUF_X1 U503 ( .A(n12412), .Z(n12408) );
  BUF_X1 U504 ( .A(n12412), .Z(n12409) );
  BUF_X1 U505 ( .A(n12412), .Z(n12410) );
  BUF_X1 U506 ( .A(n12358), .Z(n12356) );
  BUF_X1 U507 ( .A(n12358), .Z(n12355) );
  BUF_X1 U508 ( .A(n12358), .Z(n12354) );
  BUF_X1 U509 ( .A(n12358), .Z(n12353) );
  BUF_X1 U510 ( .A(n12358), .Z(n12352) );
  BUF_X1 U511 ( .A(n12358), .Z(n12351) );
  BUF_X1 U512 ( .A(n12367), .Z(n12365) );
  BUF_X1 U513 ( .A(n12367), .Z(n12364) );
  BUF_X1 U514 ( .A(n12367), .Z(n12363) );
  BUF_X1 U515 ( .A(n12367), .Z(n12362) );
  BUF_X1 U516 ( .A(n12367), .Z(n12361) );
  BUF_X1 U517 ( .A(n12367), .Z(n12360) );
  BUF_X1 U518 ( .A(n12403), .Z(n12396) );
  BUF_X1 U519 ( .A(n12403), .Z(n12397) );
  BUF_X1 U520 ( .A(n12403), .Z(n12398) );
  BUF_X1 U521 ( .A(n12403), .Z(n12399) );
  BUF_X1 U522 ( .A(n12403), .Z(n12400) );
  BUF_X1 U523 ( .A(n12403), .Z(n12401) );
  BUF_X1 U524 ( .A(n12394), .Z(n12387) );
  BUF_X1 U525 ( .A(n12394), .Z(n12388) );
  BUF_X1 U526 ( .A(n12394), .Z(n12389) );
  BUF_X1 U527 ( .A(n12394), .Z(n12390) );
  BUF_X1 U528 ( .A(n12394), .Z(n12391) );
  BUF_X1 U529 ( .A(n12394), .Z(n12392) );
  BUF_X1 U530 ( .A(n12376), .Z(n12374) );
  BUF_X1 U531 ( .A(n12376), .Z(n12373) );
  BUF_X1 U532 ( .A(n12376), .Z(n12372) );
  BUF_X1 U533 ( .A(n12376), .Z(n12371) );
  BUF_X1 U534 ( .A(n12376), .Z(n12370) );
  BUF_X1 U535 ( .A(n12376), .Z(n12369) );
  BUF_X1 U536 ( .A(n12385), .Z(n12383) );
  BUF_X1 U537 ( .A(n12385), .Z(n12382) );
  BUF_X1 U538 ( .A(n12385), .Z(n12381) );
  BUF_X1 U539 ( .A(n12385), .Z(n12380) );
  BUF_X1 U540 ( .A(n12385), .Z(n12379) );
  BUF_X1 U541 ( .A(n12385), .Z(n12378) );
  BUF_X1 U542 ( .A(n12550), .Z(n12543) );
  BUF_X1 U543 ( .A(n12550), .Z(n12544) );
  BUF_X1 U544 ( .A(n12550), .Z(n12545) );
  BUF_X1 U545 ( .A(n12550), .Z(n12546) );
  BUF_X1 U546 ( .A(n12550), .Z(n12547) );
  BUF_X1 U547 ( .A(n12550), .Z(n12548) );
  BUF_X1 U548 ( .A(n12448), .Z(n12441) );
  BUF_X1 U549 ( .A(n12448), .Z(n12442) );
  BUF_X1 U550 ( .A(n12448), .Z(n12443) );
  BUF_X1 U551 ( .A(n12448), .Z(n12444) );
  BUF_X1 U552 ( .A(n12448), .Z(n12445) );
  BUF_X1 U553 ( .A(n12448), .Z(n12446) );
  BUF_X1 U554 ( .A(n12439), .Z(n12432) );
  BUF_X1 U555 ( .A(n12439), .Z(n12433) );
  BUF_X1 U556 ( .A(n12439), .Z(n12434) );
  BUF_X1 U557 ( .A(n12439), .Z(n12435) );
  BUF_X1 U558 ( .A(n12439), .Z(n12436) );
  BUF_X1 U559 ( .A(n12439), .Z(n12437) );
  BUF_X1 U560 ( .A(n12430), .Z(n12423) );
  BUF_X1 U561 ( .A(n12430), .Z(n12424) );
  BUF_X1 U562 ( .A(n12430), .Z(n12425) );
  BUF_X1 U563 ( .A(n12430), .Z(n12426) );
  BUF_X1 U564 ( .A(n12430), .Z(n12427) );
  BUF_X1 U565 ( .A(n12430), .Z(n12428) );
  INV_X1 U566 ( .A(n1142), .ZN(n12214) );
  OAI21_X1 U567 ( .B1(n1114), .B2(n1135), .A(n12557), .ZN(n1142) );
  INV_X1 U568 ( .A(n1141), .ZN(n12223) );
  OAI21_X1 U569 ( .B1(n1116), .B2(n1135), .A(n12557), .ZN(n1141) );
  INV_X1 U570 ( .A(n1140), .ZN(n12232) );
  OAI21_X1 U571 ( .B1(n1104), .B2(n1135), .A(n12557), .ZN(n1140) );
  INV_X1 U572 ( .A(n1139), .ZN(n12241) );
  OAI21_X1 U573 ( .B1(n1107), .B2(n1135), .A(n12557), .ZN(n1139) );
  INV_X1 U574 ( .A(n1138), .ZN(n12250) );
  OAI21_X1 U575 ( .B1(n1118), .B2(n1135), .A(n12557), .ZN(n1138) );
  INV_X1 U576 ( .A(n1137), .ZN(n12259) );
  OAI21_X1 U577 ( .B1(n1120), .B2(n1135), .A(n12557), .ZN(n1137) );
  INV_X1 U578 ( .A(n1136), .ZN(n12268) );
  OAI21_X1 U579 ( .B1(n1109), .B2(n1135), .A(n12557), .ZN(n1136) );
  INV_X1 U580 ( .A(n1134), .ZN(n12277) );
  OAI21_X1 U581 ( .B1(n1111), .B2(n1135), .A(n12557), .ZN(n1134) );
  INV_X1 U582 ( .A(n1133), .ZN(n12286) );
  OAI21_X1 U583 ( .B1(n1114), .B2(n1126), .A(n12557), .ZN(n1133) );
  INV_X1 U584 ( .A(n1132), .ZN(n12295) );
  OAI21_X1 U585 ( .B1(n1116), .B2(n1126), .A(n12557), .ZN(n1132) );
  INV_X1 U586 ( .A(n1131), .ZN(n12304) );
  OAI21_X1 U587 ( .B1(n1104), .B2(n1126), .A(n12557), .ZN(n1131) );
  INV_X1 U588 ( .A(n1130), .ZN(n12313) );
  OAI21_X1 U589 ( .B1(n1107), .B2(n1126), .A(n12557), .ZN(n1130) );
  INV_X1 U590 ( .A(n1129), .ZN(n12322) );
  OAI21_X1 U591 ( .B1(n1118), .B2(n1126), .A(n12558), .ZN(n1129) );
  INV_X1 U592 ( .A(n1128), .ZN(n12331) );
  OAI21_X1 U593 ( .B1(n1120), .B2(n1126), .A(n12558), .ZN(n1128) );
  INV_X1 U594 ( .A(n1127), .ZN(n12340) );
  OAI21_X1 U595 ( .B1(n1109), .B2(n1126), .A(n12558), .ZN(n1127) );
  INV_X1 U596 ( .A(n1125), .ZN(n12349) );
  OAI21_X1 U597 ( .B1(n1111), .B2(n1126), .A(n12558), .ZN(n1125) );
  NAND2_X1 U598 ( .A1(DATAIN[14]), .A2(n12555), .ZN(n1086) );
  BUF_X1 U599 ( .A(n1095), .Z(n12475) );
  BUF_X1 U600 ( .A(n1097), .Z(n12469) );
  BUF_X1 U601 ( .A(n1098), .Z(n12466) );
  BUF_X1 U602 ( .A(n1101), .Z(n12457) );
  BUF_X1 U603 ( .A(n1102), .Z(n12454) );
  BUF_X1 U604 ( .A(n1095), .Z(n12473) );
  BUF_X1 U605 ( .A(n1097), .Z(n12467) );
  BUF_X1 U606 ( .A(n1098), .Z(n12464) );
  BUF_X1 U607 ( .A(n1101), .Z(n12455) );
  BUF_X1 U608 ( .A(n1102), .Z(n12452) );
  BUF_X1 U609 ( .A(n1095), .Z(n12474) );
  BUF_X1 U610 ( .A(n1097), .Z(n12468) );
  BUF_X1 U611 ( .A(n1098), .Z(n12465) );
  BUF_X1 U612 ( .A(n1101), .Z(n12456) );
  BUF_X1 U613 ( .A(n1102), .Z(n12453) );
  NOR3_X1 U614 ( .A1(n2471), .A2(n12567), .A3(n2472), .ZN(n2470) );
  XNOR2_X1 U615 ( .A(n12564), .B(ADD_RD2[0]), .ZN(n2471) );
  XNOR2_X1 U616 ( .A(n12566), .B(ADD_RD2[4]), .ZN(n2472) );
  OAI22_X1 U617 ( .A1(n12545), .A2(n12514), .B1(n12542), .B2(n11127), .ZN(
        n4518) );
  OAI22_X1 U618 ( .A1(n12545), .A2(n12511), .B1(n12542), .B2(n11132), .ZN(
        n4517) );
  OAI22_X1 U619 ( .A1(n12545), .A2(n12508), .B1(n12542), .B2(n11137), .ZN(
        n4516) );
  OAI22_X1 U620 ( .A1(n12545), .A2(n12505), .B1(n12542), .B2(n11142), .ZN(
        n4515) );
  OAI22_X1 U621 ( .A1(n12545), .A2(n12502), .B1(n12542), .B2(n11147), .ZN(
        n4514) );
  OAI22_X1 U622 ( .A1(n12546), .A2(n12499), .B1(n12542), .B2(n11152), .ZN(
        n4513) );
  OAI22_X1 U623 ( .A1(n12546), .A2(n12496), .B1(n12542), .B2(n11157), .ZN(
        n4512) );
  OAI22_X1 U624 ( .A1(n12546), .A2(n12493), .B1(n12542), .B2(n11162), .ZN(
        n4511) );
  OAI22_X1 U625 ( .A1(n12546), .A2(n12490), .B1(n12542), .B2(n11167), .ZN(
        n4510) );
  OAI22_X1 U626 ( .A1(n12546), .A2(n12487), .B1(n12542), .B2(n11172), .ZN(
        n4509) );
  OAI22_X1 U627 ( .A1(n12547), .A2(n12484), .B1(n12542), .B2(n11177), .ZN(
        n4508) );
  OAI22_X1 U628 ( .A1(n12547), .A2(n12481), .B1(n12542), .B2(n11181), .ZN(
        n4507) );
  OAI22_X1 U629 ( .A1(n12547), .A2(n12478), .B1(n1072), .B2(n11185), .ZN(n4506) );
  OAI22_X1 U630 ( .A1(n12547), .A2(n12475), .B1(n1072), .B2(n11189), .ZN(n4505) );
  OAI22_X1 U631 ( .A1(n12547), .A2(n12472), .B1(n1072), .B2(n11070), .ZN(n4504) );
  OAI22_X1 U632 ( .A1(n12548), .A2(n12469), .B1(n1072), .B2(n11072), .ZN(n4503) );
  OAI22_X1 U633 ( .A1(n12548), .A2(n12466), .B1(n12542), .B2(n11074), .ZN(
        n4502) );
  OAI22_X1 U634 ( .A1(n12548), .A2(n12463), .B1(n12542), .B2(n11076), .ZN(
        n4501) );
  OAI22_X1 U635 ( .A1(n12548), .A2(n12460), .B1(n12542), .B2(n11078), .ZN(
        n4500) );
  OAI22_X1 U636 ( .A1(n12548), .A2(n12457), .B1(n12542), .B2(n11080), .ZN(
        n4499) );
  OAI22_X1 U637 ( .A1(n12549), .A2(n12454), .B1(n12542), .B2(n11082), .ZN(
        n4498) );
  OAI22_X1 U638 ( .A1(n12549), .A2(n12451), .B1(n12542), .B2(n11084), .ZN(
        n4497) );
  OAI22_X1 U639 ( .A1(n12443), .A2(n12514), .B1(n12440), .B2(n11383), .ZN(
        n4486) );
  OAI22_X1 U640 ( .A1(n12443), .A2(n12511), .B1(n12440), .B2(n11388), .ZN(
        n4485) );
  OAI22_X1 U641 ( .A1(n12443), .A2(n12508), .B1(n12440), .B2(n11393), .ZN(
        n4484) );
  OAI22_X1 U642 ( .A1(n12443), .A2(n12505), .B1(n12440), .B2(n11398), .ZN(
        n4483) );
  OAI22_X1 U643 ( .A1(n12443), .A2(n12502), .B1(n12440), .B2(n11403), .ZN(
        n4482) );
  OAI22_X1 U644 ( .A1(n12444), .A2(n12499), .B1(n12440), .B2(n11408), .ZN(
        n4481) );
  OAI22_X1 U645 ( .A1(n12444), .A2(n12496), .B1(n12440), .B2(n11413), .ZN(
        n4480) );
  OAI22_X1 U646 ( .A1(n12444), .A2(n12493), .B1(n12440), .B2(n11418), .ZN(
        n4479) );
  OAI22_X1 U647 ( .A1(n12444), .A2(n12490), .B1(n12440), .B2(n11423), .ZN(
        n4478) );
  OAI22_X1 U648 ( .A1(n12444), .A2(n12487), .B1(n12440), .B2(n11428), .ZN(
        n4477) );
  OAI22_X1 U649 ( .A1(n12445), .A2(n12484), .B1(n12440), .B2(n11433), .ZN(
        n4476) );
  OAI22_X1 U650 ( .A1(n12445), .A2(n12481), .B1(n12440), .B2(n11437), .ZN(
        n4475) );
  OAI22_X1 U651 ( .A1(n12445), .A2(n12478), .B1(n1106), .B2(n11441), .ZN(n4474) );
  OAI22_X1 U652 ( .A1(n12445), .A2(n12475), .B1(n1106), .B2(n11445), .ZN(n4473) );
  OAI22_X1 U653 ( .A1(n12445), .A2(n12472), .B1(n1106), .B2(n11326), .ZN(n4472) );
  OAI22_X1 U654 ( .A1(n12446), .A2(n12469), .B1(n1106), .B2(n11328), .ZN(n4471) );
  OAI22_X1 U655 ( .A1(n12446), .A2(n12466), .B1(n12440), .B2(n11330), .ZN(
        n4470) );
  OAI22_X1 U656 ( .A1(n12446), .A2(n12463), .B1(n12440), .B2(n11332), .ZN(
        n4469) );
  OAI22_X1 U657 ( .A1(n12446), .A2(n12460), .B1(n12440), .B2(n11334), .ZN(
        n4468) );
  OAI22_X1 U658 ( .A1(n12446), .A2(n12457), .B1(n12440), .B2(n11336), .ZN(
        n4467) );
  OAI22_X1 U659 ( .A1(n12447), .A2(n12454), .B1(n12440), .B2(n11338), .ZN(
        n4466) );
  OAI22_X1 U660 ( .A1(n12447), .A2(n12451), .B1(n12440), .B2(n11340), .ZN(
        n4465) );
  OAI22_X1 U661 ( .A1(n12434), .A2(n12514), .B1(n12431), .B2(n11128), .ZN(
        n4454) );
  OAI22_X1 U662 ( .A1(n12434), .A2(n12511), .B1(n12431), .B2(n11133), .ZN(
        n4453) );
  OAI22_X1 U663 ( .A1(n12434), .A2(n12508), .B1(n12431), .B2(n11138), .ZN(
        n4452) );
  OAI22_X1 U664 ( .A1(n12434), .A2(n12505), .B1(n12431), .B2(n11143), .ZN(
        n4451) );
  OAI22_X1 U665 ( .A1(n12434), .A2(n12502), .B1(n12431), .B2(n11148), .ZN(
        n4450) );
  OAI22_X1 U666 ( .A1(n12435), .A2(n12499), .B1(n12431), .B2(n11153), .ZN(
        n4449) );
  OAI22_X1 U667 ( .A1(n12435), .A2(n12496), .B1(n12431), .B2(n11158), .ZN(
        n4448) );
  OAI22_X1 U668 ( .A1(n12435), .A2(n12493), .B1(n12431), .B2(n11163), .ZN(
        n4447) );
  OAI22_X1 U669 ( .A1(n12435), .A2(n12490), .B1(n12431), .B2(n11168), .ZN(
        n4446) );
  OAI22_X1 U670 ( .A1(n12435), .A2(n12487), .B1(n12431), .B2(n11173), .ZN(
        n4445) );
  OAI22_X1 U671 ( .A1(n12436), .A2(n12484), .B1(n12431), .B2(n10991), .ZN(
        n4444) );
  OAI22_X1 U672 ( .A1(n12436), .A2(n12481), .B1(n12431), .B2(n10992), .ZN(
        n4443) );
  OAI22_X1 U673 ( .A1(n12436), .A2(n12478), .B1(n1108), .B2(n10993), .ZN(n4442) );
  OAI22_X1 U674 ( .A1(n12436), .A2(n12475), .B1(n1108), .B2(n10994), .ZN(n4441) );
  OAI22_X1 U675 ( .A1(n12436), .A2(n12472), .B1(n1108), .B2(n10995), .ZN(n4440) );
  OAI22_X1 U676 ( .A1(n12437), .A2(n12469), .B1(n1108), .B2(n10976), .ZN(n4439) );
  OAI22_X1 U677 ( .A1(n12437), .A2(n12466), .B1(n12431), .B2(n10977), .ZN(
        n4438) );
  OAI22_X1 U678 ( .A1(n12437), .A2(n12463), .B1(n12431), .B2(n10978), .ZN(
        n4437) );
  OAI22_X1 U679 ( .A1(n12437), .A2(n12460), .B1(n12431), .B2(n10979), .ZN(
        n4436) );
  OAI22_X1 U680 ( .A1(n12437), .A2(n12457), .B1(n12431), .B2(n10980), .ZN(
        n4435) );
  OAI22_X1 U681 ( .A1(n12438), .A2(n12454), .B1(n12431), .B2(n10981), .ZN(
        n4434) );
  OAI22_X1 U682 ( .A1(n12438), .A2(n12451), .B1(n12431), .B2(n10982), .ZN(
        n4433) );
  OAI22_X1 U683 ( .A1(n12425), .A2(n12514), .B1(n12422), .B2(n11384), .ZN(
        n4422) );
  OAI22_X1 U684 ( .A1(n12425), .A2(n12511), .B1(n12422), .B2(n11389), .ZN(
        n4421) );
  OAI22_X1 U685 ( .A1(n12425), .A2(n12508), .B1(n12422), .B2(n11394), .ZN(
        n4420) );
  OAI22_X1 U686 ( .A1(n12425), .A2(n12505), .B1(n12422), .B2(n11399), .ZN(
        n4419) );
  OAI22_X1 U687 ( .A1(n12425), .A2(n12502), .B1(n12422), .B2(n11404), .ZN(
        n4418) );
  OAI22_X1 U688 ( .A1(n12426), .A2(n12499), .B1(n12422), .B2(n11409), .ZN(
        n4417) );
  OAI22_X1 U689 ( .A1(n12426), .A2(n12496), .B1(n12422), .B2(n11414), .ZN(
        n4416) );
  OAI22_X1 U690 ( .A1(n12426), .A2(n12493), .B1(n12422), .B2(n11419), .ZN(
        n4415) );
  OAI22_X1 U691 ( .A1(n12426), .A2(n12490), .B1(n12422), .B2(n11424), .ZN(
        n4414) );
  OAI22_X1 U692 ( .A1(n12426), .A2(n12487), .B1(n12422), .B2(n11429), .ZN(
        n4413) );
  OAI22_X1 U693 ( .A1(n12427), .A2(n12484), .B1(n12422), .B2(n11247), .ZN(
        n4412) );
  OAI22_X1 U694 ( .A1(n12427), .A2(n12481), .B1(n12422), .B2(n11248), .ZN(
        n4411) );
  OAI22_X1 U695 ( .A1(n12427), .A2(n12478), .B1(n1110), .B2(n11249), .ZN(n4410) );
  OAI22_X1 U696 ( .A1(n12427), .A2(n12475), .B1(n1110), .B2(n11250), .ZN(n4409) );
  OAI22_X1 U697 ( .A1(n12427), .A2(n12472), .B1(n1110), .B2(n11251), .ZN(n4408) );
  OAI22_X1 U698 ( .A1(n12428), .A2(n12469), .B1(n1110), .B2(n11232), .ZN(n4407) );
  OAI22_X1 U699 ( .A1(n12428), .A2(n12466), .B1(n12422), .B2(n11233), .ZN(
        n4406) );
  OAI22_X1 U700 ( .A1(n12428), .A2(n12463), .B1(n12422), .B2(n11234), .ZN(
        n4405) );
  OAI22_X1 U701 ( .A1(n12428), .A2(n12460), .B1(n12422), .B2(n11235), .ZN(
        n4404) );
  OAI22_X1 U702 ( .A1(n12428), .A2(n12457), .B1(n12422), .B2(n11236), .ZN(
        n4403) );
  OAI22_X1 U703 ( .A1(n12429), .A2(n12454), .B1(n12422), .B2(n11237), .ZN(
        n4402) );
  OAI22_X1 U704 ( .A1(n12429), .A2(n12451), .B1(n12422), .B2(n11238), .ZN(
        n4401) );
  OAI22_X1 U705 ( .A1(n12231), .A2(n12551), .B1(n12224), .B2(n11020), .ZN(
        n2923) );
  OAI22_X1 U706 ( .A1(n12231), .A2(n12539), .B1(n12224), .B2(n11022), .ZN(
        n2924) );
  OAI22_X1 U707 ( .A1(n12230), .A2(n12536), .B1(n12224), .B2(n11024), .ZN(
        n2925) );
  OAI22_X1 U708 ( .A1(n12230), .A2(n12533), .B1(n12224), .B2(n11026), .ZN(
        n2926) );
  OAI22_X1 U709 ( .A1(n12230), .A2(n12530), .B1(n12224), .B2(n11028), .ZN(
        n2927) );
  OAI22_X1 U710 ( .A1(n12230), .A2(n12527), .B1(n12224), .B2(n11030), .ZN(
        n2928) );
  OAI22_X1 U711 ( .A1(n12230), .A2(n12524), .B1(n12224), .B2(n11032), .ZN(
        n2929) );
  OAI22_X1 U712 ( .A1(n12229), .A2(n12521), .B1(n12224), .B2(n11034), .ZN(
        n2930) );
  OAI22_X1 U713 ( .A1(n12229), .A2(n12518), .B1(n12224), .B2(n10996), .ZN(
        n2931) );
  OAI22_X1 U714 ( .A1(n12229), .A2(n12515), .B1(n12224), .B2(n11121), .ZN(
        n2932) );
  OAI22_X1 U715 ( .A1(n12229), .A2(n12512), .B1(n12224), .B2(n11126), .ZN(
        n2933) );
  OAI22_X1 U716 ( .A1(n12229), .A2(n12509), .B1(n12224), .B2(n11131), .ZN(
        n2934) );
  OAI22_X1 U717 ( .A1(n12228), .A2(n12506), .B1(n1140), .B2(n11136), .ZN(n2935) );
  OAI22_X1 U718 ( .A1(n12228), .A2(n12503), .B1(n1140), .B2(n11141), .ZN(n2936) );
  OAI22_X1 U719 ( .A1(n12228), .A2(n12500), .B1(n1140), .B2(n11146), .ZN(n2937) );
  OAI22_X1 U720 ( .A1(n12228), .A2(n12497), .B1(n1140), .B2(n11151), .ZN(n2938) );
  OAI22_X1 U721 ( .A1(n12228), .A2(n12494), .B1(n12224), .B2(n11156), .ZN(
        n2939) );
  OAI22_X1 U722 ( .A1(n12227), .A2(n12491), .B1(n12224), .B2(n11161), .ZN(
        n2940) );
  OAI22_X1 U723 ( .A1(n12227), .A2(n12488), .B1(n12224), .B2(n11166), .ZN(
        n2941) );
  OAI22_X1 U724 ( .A1(n12227), .A2(n12485), .B1(n12224), .B2(n11171), .ZN(
        n2942) );
  OAI22_X1 U725 ( .A1(n12227), .A2(n12482), .B1(n12224), .B2(n11176), .ZN(
        n2943) );
  OAI22_X1 U726 ( .A1(n12227), .A2(n12479), .B1(n12224), .B2(n11180), .ZN(
        n2944) );
  OAI22_X1 U727 ( .A1(n12240), .A2(n12551), .B1(n12233), .B2(n11276), .ZN(
        n2955) );
  OAI22_X1 U728 ( .A1(n12240), .A2(n12539), .B1(n12233), .B2(n11278), .ZN(
        n2956) );
  OAI22_X1 U729 ( .A1(n12239), .A2(n12536), .B1(n12233), .B2(n11280), .ZN(
        n2957) );
  OAI22_X1 U730 ( .A1(n12239), .A2(n12533), .B1(n12233), .B2(n11282), .ZN(
        n2958) );
  OAI22_X1 U731 ( .A1(n12239), .A2(n12530), .B1(n12233), .B2(n11284), .ZN(
        n2959) );
  OAI22_X1 U732 ( .A1(n12239), .A2(n12527), .B1(n12233), .B2(n11286), .ZN(
        n2960) );
  OAI22_X1 U733 ( .A1(n12239), .A2(n12524), .B1(n12233), .B2(n11288), .ZN(
        n2961) );
  OAI22_X1 U734 ( .A1(n12238), .A2(n12521), .B1(n12233), .B2(n11290), .ZN(
        n2962) );
  OAI22_X1 U735 ( .A1(n12238), .A2(n12518), .B1(n12233), .B2(n11252), .ZN(
        n2963) );
  OAI22_X1 U736 ( .A1(n12238), .A2(n12515), .B1(n12233), .B2(n11377), .ZN(
        n2964) );
  OAI22_X1 U737 ( .A1(n12238), .A2(n12512), .B1(n12233), .B2(n11382), .ZN(
        n2965) );
  OAI22_X1 U738 ( .A1(n12238), .A2(n12509), .B1(n12233), .B2(n11387), .ZN(
        n2966) );
  OAI22_X1 U739 ( .A1(n12237), .A2(n12506), .B1(n1139), .B2(n11392), .ZN(n2967) );
  OAI22_X1 U740 ( .A1(n12237), .A2(n12503), .B1(n1139), .B2(n11397), .ZN(n2968) );
  OAI22_X1 U741 ( .A1(n12237), .A2(n12500), .B1(n1139), .B2(n11402), .ZN(n2969) );
  OAI22_X1 U742 ( .A1(n12237), .A2(n12497), .B1(n1139), .B2(n11407), .ZN(n2970) );
  OAI22_X1 U743 ( .A1(n12237), .A2(n12494), .B1(n12233), .B2(n11412), .ZN(
        n2971) );
  OAI22_X1 U744 ( .A1(n12236), .A2(n12491), .B1(n12233), .B2(n11417), .ZN(
        n2972) );
  OAI22_X1 U745 ( .A1(n12236), .A2(n12488), .B1(n12233), .B2(n11422), .ZN(
        n2973) );
  OAI22_X1 U746 ( .A1(n12236), .A2(n12485), .B1(n12233), .B2(n11427), .ZN(
        n2974) );
  OAI22_X1 U747 ( .A1(n12236), .A2(n12482), .B1(n12233), .B2(n11432), .ZN(
        n2975) );
  OAI22_X1 U748 ( .A1(n12236), .A2(n12479), .B1(n12233), .B2(n11436), .ZN(
        n2976) );
  OAI22_X1 U749 ( .A1(n12267), .A2(n12552), .B1(n12260), .B2(n11087), .ZN(
        n3051) );
  OAI22_X1 U750 ( .A1(n12267), .A2(n12540), .B1(n12260), .B2(n11091), .ZN(
        n3052) );
  OAI22_X1 U751 ( .A1(n12266), .A2(n12537), .B1(n12260), .B2(n11095), .ZN(
        n3053) );
  OAI22_X1 U752 ( .A1(n12266), .A2(n12534), .B1(n12260), .B2(n11099), .ZN(
        n3054) );
  OAI22_X1 U753 ( .A1(n12266), .A2(n12531), .B1(n12260), .B2(n11103), .ZN(
        n3055) );
  OAI22_X1 U754 ( .A1(n12266), .A2(n12528), .B1(n12260), .B2(n11107), .ZN(
        n3056) );
  OAI22_X1 U755 ( .A1(n12266), .A2(n12525), .B1(n12260), .B2(n11111), .ZN(
        n3057) );
  OAI22_X1 U756 ( .A1(n12265), .A2(n12522), .B1(n12260), .B2(n11115), .ZN(
        n3058) );
  OAI22_X1 U757 ( .A1(n12265), .A2(n12519), .B1(n12260), .B2(n11118), .ZN(
        n3059) );
  OAI22_X1 U758 ( .A1(n12265), .A2(n12516), .B1(n12260), .B2(n11124), .ZN(
        n3060) );
  OAI22_X1 U759 ( .A1(n12265), .A2(n12513), .B1(n12260), .B2(n11129), .ZN(
        n3061) );
  OAI22_X1 U760 ( .A1(n12265), .A2(n12510), .B1(n12260), .B2(n11134), .ZN(
        n3062) );
  OAI22_X1 U761 ( .A1(n12264), .A2(n12507), .B1(n1136), .B2(n11139), .ZN(n3063) );
  OAI22_X1 U762 ( .A1(n12264), .A2(n12504), .B1(n1136), .B2(n11144), .ZN(n3064) );
  OAI22_X1 U763 ( .A1(n12264), .A2(n12501), .B1(n1136), .B2(n11149), .ZN(n3065) );
  OAI22_X1 U764 ( .A1(n12264), .A2(n12498), .B1(n1136), .B2(n11154), .ZN(n3066) );
  OAI22_X1 U765 ( .A1(n12264), .A2(n12495), .B1(n12260), .B2(n11159), .ZN(
        n3067) );
  OAI22_X1 U766 ( .A1(n12263), .A2(n12492), .B1(n12260), .B2(n11164), .ZN(
        n3068) );
  OAI22_X1 U767 ( .A1(n12263), .A2(n12489), .B1(n12260), .B2(n11169), .ZN(
        n3069) );
  OAI22_X1 U768 ( .A1(n12263), .A2(n12486), .B1(n12260), .B2(n11174), .ZN(
        n3070) );
  OAI22_X1 U769 ( .A1(n12263), .A2(n12483), .B1(n12260), .B2(n11178), .ZN(
        n3071) );
  OAI22_X1 U770 ( .A1(n12263), .A2(n12480), .B1(n12260), .B2(n11182), .ZN(
        n3072) );
  OAI22_X1 U771 ( .A1(n12276), .A2(n12552), .B1(n12269), .B2(n11343), .ZN(
        n3083) );
  OAI22_X1 U772 ( .A1(n12276), .A2(n12540), .B1(n12269), .B2(n11347), .ZN(
        n3084) );
  OAI22_X1 U773 ( .A1(n12275), .A2(n12537), .B1(n12269), .B2(n11351), .ZN(
        n3085) );
  OAI22_X1 U774 ( .A1(n12275), .A2(n12534), .B1(n12269), .B2(n11355), .ZN(
        n3086) );
  OAI22_X1 U775 ( .A1(n12275), .A2(n12531), .B1(n12269), .B2(n11359), .ZN(
        n3087) );
  OAI22_X1 U776 ( .A1(n12275), .A2(n12528), .B1(n12269), .B2(n11363), .ZN(
        n3088) );
  OAI22_X1 U777 ( .A1(n12275), .A2(n12525), .B1(n12269), .B2(n11367), .ZN(
        n3089) );
  OAI22_X1 U778 ( .A1(n12274), .A2(n12522), .B1(n12269), .B2(n11371), .ZN(
        n3090) );
  OAI22_X1 U779 ( .A1(n12274), .A2(n12519), .B1(n12269), .B2(n11374), .ZN(
        n3091) );
  OAI22_X1 U780 ( .A1(n12274), .A2(n12516), .B1(n12269), .B2(n11380), .ZN(
        n3092) );
  OAI22_X1 U781 ( .A1(n12274), .A2(n12513), .B1(n12269), .B2(n11385), .ZN(
        n3093) );
  OAI22_X1 U782 ( .A1(n12274), .A2(n12510), .B1(n12269), .B2(n11390), .ZN(
        n3094) );
  OAI22_X1 U783 ( .A1(n12273), .A2(n12507), .B1(n1134), .B2(n11395), .ZN(n3095) );
  OAI22_X1 U784 ( .A1(n12273), .A2(n12504), .B1(n1134), .B2(n11400), .ZN(n3096) );
  OAI22_X1 U785 ( .A1(n12273), .A2(n12501), .B1(n1134), .B2(n11405), .ZN(n3097) );
  OAI22_X1 U786 ( .A1(n12273), .A2(n12498), .B1(n1134), .B2(n11410), .ZN(n3098) );
  OAI22_X1 U787 ( .A1(n12273), .A2(n12495), .B1(n12269), .B2(n11415), .ZN(
        n3099) );
  OAI22_X1 U788 ( .A1(n12272), .A2(n12492), .B1(n12269), .B2(n11420), .ZN(
        n3100) );
  OAI22_X1 U789 ( .A1(n12272), .A2(n12489), .B1(n12269), .B2(n11425), .ZN(
        n3101) );
  OAI22_X1 U790 ( .A1(n12272), .A2(n12486), .B1(n12269), .B2(n11430), .ZN(
        n3102) );
  OAI22_X1 U791 ( .A1(n12272), .A2(n12483), .B1(n12269), .B2(n11434), .ZN(
        n3103) );
  OAI22_X1 U792 ( .A1(n12272), .A2(n12480), .B1(n12269), .B2(n11438), .ZN(
        n3104) );
  OAI22_X1 U793 ( .A1(n12303), .A2(n12552), .B1(n12296), .B2(n10951), .ZN(
        n3179) );
  OAI22_X1 U794 ( .A1(n12303), .A2(n12540), .B1(n12296), .B2(n10952), .ZN(
        n3180) );
  OAI22_X1 U795 ( .A1(n12302), .A2(n12537), .B1(n12296), .B2(n10953), .ZN(
        n3181) );
  OAI22_X1 U796 ( .A1(n12302), .A2(n12534), .B1(n12296), .B2(n10954), .ZN(
        n3182) );
  OAI22_X1 U797 ( .A1(n12302), .A2(n12531), .B1(n12296), .B2(n10955), .ZN(
        n3183) );
  OAI22_X1 U798 ( .A1(n12302), .A2(n12528), .B1(n12296), .B2(n10956), .ZN(
        n3184) );
  OAI22_X1 U799 ( .A1(n12302), .A2(n12525), .B1(n12296), .B2(n10957), .ZN(
        n3185) );
  OAI22_X1 U800 ( .A1(n12301), .A2(n12522), .B1(n12296), .B2(n10958), .ZN(
        n3186) );
  OAI22_X1 U801 ( .A1(n12301), .A2(n12519), .B1(n12296), .B2(n11119), .ZN(
        n3187) );
  OAI22_X1 U802 ( .A1(n12301), .A2(n12516), .B1(n12296), .B2(n10936), .ZN(
        n3188) );
  OAI22_X1 U803 ( .A1(n12301), .A2(n12513), .B1(n12296), .B2(n10937), .ZN(
        n3189) );
  OAI22_X1 U804 ( .A1(n12301), .A2(n12510), .B1(n12296), .B2(n10938), .ZN(
        n3190) );
  OAI22_X1 U805 ( .A1(n12300), .A2(n12507), .B1(n1131), .B2(n10939), .ZN(n3191) );
  OAI22_X1 U806 ( .A1(n12300), .A2(n12504), .B1(n1131), .B2(n10940), .ZN(n3192) );
  OAI22_X1 U807 ( .A1(n12300), .A2(n12501), .B1(n1131), .B2(n10941), .ZN(n3193) );
  OAI22_X1 U808 ( .A1(n12300), .A2(n12498), .B1(n1131), .B2(n10942), .ZN(n3194) );
  OAI22_X1 U809 ( .A1(n12300), .A2(n12495), .B1(n12296), .B2(n10943), .ZN(
        n3195) );
  OAI22_X1 U810 ( .A1(n12299), .A2(n12492), .B1(n12296), .B2(n10944), .ZN(
        n3196) );
  OAI22_X1 U811 ( .A1(n12299), .A2(n12489), .B1(n12296), .B2(n10945), .ZN(
        n3197) );
  OAI22_X1 U812 ( .A1(n12299), .A2(n12486), .B1(n12296), .B2(n10946), .ZN(
        n3198) );
  OAI22_X1 U813 ( .A1(n12299), .A2(n12483), .B1(n12296), .B2(n10947), .ZN(
        n3199) );
  OAI22_X1 U814 ( .A1(n12299), .A2(n12480), .B1(n12296), .B2(n10948), .ZN(
        n3200) );
  OAI22_X1 U815 ( .A1(n12312), .A2(n12552), .B1(n12305), .B2(n11207), .ZN(
        n3211) );
  OAI22_X1 U816 ( .A1(n12312), .A2(n12540), .B1(n12305), .B2(n11208), .ZN(
        n3212) );
  OAI22_X1 U817 ( .A1(n12311), .A2(n12537), .B1(n12305), .B2(n11209), .ZN(
        n3213) );
  OAI22_X1 U818 ( .A1(n12311), .A2(n12534), .B1(n12305), .B2(n11210), .ZN(
        n3214) );
  OAI22_X1 U819 ( .A1(n12311), .A2(n12531), .B1(n12305), .B2(n11211), .ZN(
        n3215) );
  OAI22_X1 U820 ( .A1(n12311), .A2(n12528), .B1(n12305), .B2(n11212), .ZN(
        n3216) );
  OAI22_X1 U821 ( .A1(n12311), .A2(n12525), .B1(n12305), .B2(n11213), .ZN(
        n3217) );
  OAI22_X1 U822 ( .A1(n12310), .A2(n12522), .B1(n12305), .B2(n11214), .ZN(
        n3218) );
  OAI22_X1 U823 ( .A1(n12310), .A2(n12519), .B1(n12305), .B2(n11375), .ZN(
        n3219) );
  OAI22_X1 U824 ( .A1(n12310), .A2(n12516), .B1(n12305), .B2(n11192), .ZN(
        n3220) );
  OAI22_X1 U825 ( .A1(n12310), .A2(n12513), .B1(n12305), .B2(n11193), .ZN(
        n3221) );
  OAI22_X1 U826 ( .A1(n12310), .A2(n12510), .B1(n12305), .B2(n11194), .ZN(
        n3222) );
  OAI22_X1 U827 ( .A1(n12309), .A2(n12507), .B1(n1130), .B2(n11195), .ZN(n3223) );
  OAI22_X1 U828 ( .A1(n12309), .A2(n12504), .B1(n1130), .B2(n11196), .ZN(n3224) );
  OAI22_X1 U829 ( .A1(n12309), .A2(n12501), .B1(n1130), .B2(n11197), .ZN(n3225) );
  OAI22_X1 U830 ( .A1(n12309), .A2(n12498), .B1(n1130), .B2(n11198), .ZN(n3226) );
  OAI22_X1 U831 ( .A1(n12309), .A2(n12495), .B1(n12305), .B2(n11199), .ZN(
        n3227) );
  OAI22_X1 U832 ( .A1(n12308), .A2(n12492), .B1(n12305), .B2(n11200), .ZN(
        n3228) );
  OAI22_X1 U833 ( .A1(n12308), .A2(n12489), .B1(n12305), .B2(n11201), .ZN(
        n3229) );
  OAI22_X1 U834 ( .A1(n12308), .A2(n12486), .B1(n12305), .B2(n11202), .ZN(
        n3230) );
  OAI22_X1 U835 ( .A1(n12308), .A2(n12483), .B1(n12305), .B2(n11203), .ZN(
        n3231) );
  OAI22_X1 U836 ( .A1(n12308), .A2(n12480), .B1(n12305), .B2(n11204), .ZN(
        n3232) );
  OAI22_X1 U837 ( .A1(n12339), .A2(n12552), .B1(n12332), .B2(n10983), .ZN(
        n3307) );
  OAI22_X1 U838 ( .A1(n12339), .A2(n12540), .B1(n12332), .B2(n10984), .ZN(
        n3308) );
  OAI22_X1 U839 ( .A1(n12338), .A2(n12537), .B1(n12332), .B2(n10985), .ZN(
        n3309) );
  OAI22_X1 U840 ( .A1(n12338), .A2(n12534), .B1(n12332), .B2(n10986), .ZN(
        n3310) );
  OAI22_X1 U841 ( .A1(n12338), .A2(n12531), .B1(n12332), .B2(n10987), .ZN(
        n3311) );
  OAI22_X1 U842 ( .A1(n12338), .A2(n12528), .B1(n12332), .B2(n10988), .ZN(
        n3312) );
  OAI22_X1 U843 ( .A1(n12338), .A2(n12525), .B1(n12332), .B2(n10989), .ZN(
        n3313) );
  OAI22_X1 U844 ( .A1(n12337), .A2(n12522), .B1(n12332), .B2(n10990), .ZN(
        n3314) );
  OAI22_X1 U845 ( .A1(n12337), .A2(n12519), .B1(n12332), .B2(n10960), .ZN(
        n3315) );
  OAI22_X1 U846 ( .A1(n12337), .A2(n12516), .B1(n12332), .B2(n10961), .ZN(
        n3316) );
  OAI22_X1 U847 ( .A1(n12337), .A2(n12513), .B1(n12332), .B2(n10962), .ZN(
        n3317) );
  OAI22_X1 U848 ( .A1(n12337), .A2(n12510), .B1(n12332), .B2(n10963), .ZN(
        n3318) );
  OAI22_X1 U849 ( .A1(n12336), .A2(n12507), .B1(n1127), .B2(n10964), .ZN(n3319) );
  OAI22_X1 U850 ( .A1(n12336), .A2(n12504), .B1(n1127), .B2(n10965), .ZN(n3320) );
  OAI22_X1 U851 ( .A1(n12336), .A2(n12501), .B1(n1127), .B2(n10966), .ZN(n3321) );
  OAI22_X1 U852 ( .A1(n12336), .A2(n12498), .B1(n1127), .B2(n10967), .ZN(n3322) );
  OAI22_X1 U853 ( .A1(n12336), .A2(n12495), .B1(n12332), .B2(n10968), .ZN(
        n3323) );
  OAI22_X1 U854 ( .A1(n12335), .A2(n12492), .B1(n12332), .B2(n10969), .ZN(
        n3324) );
  OAI22_X1 U855 ( .A1(n12335), .A2(n12489), .B1(n12332), .B2(n10970), .ZN(
        n3325) );
  OAI22_X1 U856 ( .A1(n12335), .A2(n12486), .B1(n12332), .B2(n10971), .ZN(
        n3326) );
  OAI22_X1 U857 ( .A1(n12335), .A2(n12483), .B1(n12332), .B2(n10972), .ZN(
        n3327) );
  OAI22_X1 U858 ( .A1(n12335), .A2(n12480), .B1(n12332), .B2(n10973), .ZN(
        n3328) );
  OAI22_X1 U859 ( .A1(n12348), .A2(n12552), .B1(n12341), .B2(n11239), .ZN(
        n3339) );
  OAI22_X1 U860 ( .A1(n12348), .A2(n12540), .B1(n12341), .B2(n11240), .ZN(
        n3340) );
  OAI22_X1 U861 ( .A1(n12347), .A2(n12537), .B1(n12341), .B2(n11241), .ZN(
        n3341) );
  OAI22_X1 U862 ( .A1(n12347), .A2(n12534), .B1(n12341), .B2(n11242), .ZN(
        n3342) );
  OAI22_X1 U863 ( .A1(n12347), .A2(n12531), .B1(n12341), .B2(n11243), .ZN(
        n3343) );
  OAI22_X1 U864 ( .A1(n12347), .A2(n12528), .B1(n12341), .B2(n11244), .ZN(
        n3344) );
  OAI22_X1 U865 ( .A1(n12347), .A2(n12525), .B1(n12341), .B2(n11245), .ZN(
        n3345) );
  OAI22_X1 U866 ( .A1(n12346), .A2(n12522), .B1(n12341), .B2(n11246), .ZN(
        n3346) );
  OAI22_X1 U867 ( .A1(n12346), .A2(n12519), .B1(n12341), .B2(n11216), .ZN(
        n3347) );
  OAI22_X1 U868 ( .A1(n12346), .A2(n12516), .B1(n12341), .B2(n11217), .ZN(
        n3348) );
  OAI22_X1 U869 ( .A1(n12346), .A2(n12513), .B1(n12341), .B2(n11218), .ZN(
        n3349) );
  OAI22_X1 U870 ( .A1(n12346), .A2(n12510), .B1(n12341), .B2(n11219), .ZN(
        n3350) );
  OAI22_X1 U871 ( .A1(n12345), .A2(n12507), .B1(n1125), .B2(n11220), .ZN(n3351) );
  OAI22_X1 U872 ( .A1(n12345), .A2(n12504), .B1(n1125), .B2(n11221), .ZN(n3352) );
  OAI22_X1 U873 ( .A1(n12345), .A2(n12501), .B1(n1125), .B2(n11222), .ZN(n3353) );
  OAI22_X1 U874 ( .A1(n12345), .A2(n12498), .B1(n1125), .B2(n11223), .ZN(n3354) );
  OAI22_X1 U875 ( .A1(n12345), .A2(n12495), .B1(n12341), .B2(n11224), .ZN(
        n3355) );
  OAI22_X1 U876 ( .A1(n12344), .A2(n12492), .B1(n12341), .B2(n11225), .ZN(
        n3356) );
  OAI22_X1 U877 ( .A1(n12344), .A2(n12489), .B1(n12341), .B2(n11226), .ZN(
        n3357) );
  OAI22_X1 U878 ( .A1(n12344), .A2(n12486), .B1(n12341), .B2(n11227), .ZN(
        n3358) );
  OAI22_X1 U879 ( .A1(n12344), .A2(n12483), .B1(n12341), .B2(n11228), .ZN(
        n3359) );
  OAI22_X1 U880 ( .A1(n12344), .A2(n12480), .B1(n12341), .B2(n11229), .ZN(
        n3360) );
  OAI22_X1 U881 ( .A1(n12416), .A2(n12514), .B1(n12413), .B2(n11255), .ZN(
        n4390) );
  OAI22_X1 U882 ( .A1(n12416), .A2(n12511), .B1(n12413), .B2(n11256), .ZN(
        n4389) );
  OAI22_X1 U883 ( .A1(n12416), .A2(n12508), .B1(n12413), .B2(n11257), .ZN(
        n4388) );
  OAI22_X1 U884 ( .A1(n12416), .A2(n12505), .B1(n12413), .B2(n11258), .ZN(
        n4387) );
  OAI22_X1 U885 ( .A1(n12416), .A2(n12502), .B1(n12413), .B2(n11259), .ZN(
        n4386) );
  OAI22_X1 U886 ( .A1(n12417), .A2(n12499), .B1(n12413), .B2(n11260), .ZN(
        n4385) );
  OAI22_X1 U887 ( .A1(n12417), .A2(n12496), .B1(n12413), .B2(n11261), .ZN(
        n4384) );
  OAI22_X1 U888 ( .A1(n12417), .A2(n12493), .B1(n12413), .B2(n11262), .ZN(
        n4383) );
  OAI22_X1 U889 ( .A1(n12417), .A2(n12490), .B1(n12413), .B2(n11263), .ZN(
        n4382) );
  OAI22_X1 U890 ( .A1(n12417), .A2(n12487), .B1(n12413), .B2(n11264), .ZN(
        n4381) );
  OAI22_X1 U891 ( .A1(n12418), .A2(n12484), .B1(n12413), .B2(n11265), .ZN(
        n4380) );
  OAI22_X1 U892 ( .A1(n12418), .A2(n12481), .B1(n12413), .B2(n11266), .ZN(
        n4379) );
  OAI22_X1 U893 ( .A1(n12418), .A2(n12478), .B1(n1112), .B2(n11267), .ZN(n4378) );
  OAI22_X1 U894 ( .A1(n12418), .A2(n12475), .B1(n1112), .B2(n11268), .ZN(n4377) );
  OAI22_X1 U895 ( .A1(n12418), .A2(n12472), .B1(n1112), .B2(n11317), .ZN(n4376) );
  OAI22_X1 U896 ( .A1(n12419), .A2(n12469), .B1(n1112), .B2(n11318), .ZN(n4375) );
  OAI22_X1 U897 ( .A1(n12419), .A2(n12466), .B1(n12413), .B2(n11319), .ZN(
        n4374) );
  OAI22_X1 U898 ( .A1(n12419), .A2(n12463), .B1(n12413), .B2(n11320), .ZN(
        n4373) );
  OAI22_X1 U899 ( .A1(n12419), .A2(n12460), .B1(n12413), .B2(n11321), .ZN(
        n4372) );
  OAI22_X1 U900 ( .A1(n12419), .A2(n12457), .B1(n12413), .B2(n11322), .ZN(
        n4371) );
  OAI22_X1 U901 ( .A1(n12420), .A2(n12454), .B1(n12413), .B2(n11323), .ZN(
        n4370) );
  OAI22_X1 U902 ( .A1(n12420), .A2(n12451), .B1(n12413), .B2(n11324), .ZN(
        n4369) );
  OAI22_X1 U903 ( .A1(n12407), .A2(n12514), .B1(n12404), .B2(n10999), .ZN(
        n4358) );
  OAI22_X1 U904 ( .A1(n12407), .A2(n12511), .B1(n12404), .B2(n11000), .ZN(
        n4357) );
  OAI22_X1 U905 ( .A1(n12407), .A2(n12508), .B1(n12404), .B2(n11001), .ZN(
        n4356) );
  OAI22_X1 U906 ( .A1(n12407), .A2(n12505), .B1(n12404), .B2(n11002), .ZN(
        n4355) );
  OAI22_X1 U907 ( .A1(n12407), .A2(n12502), .B1(n12404), .B2(n11003), .ZN(
        n4354) );
  OAI22_X1 U908 ( .A1(n12408), .A2(n12499), .B1(n12404), .B2(n11004), .ZN(
        n4353) );
  OAI22_X1 U909 ( .A1(n12408), .A2(n12496), .B1(n12404), .B2(n11005), .ZN(
        n4352) );
  OAI22_X1 U910 ( .A1(n12408), .A2(n12493), .B1(n12404), .B2(n11006), .ZN(
        n4351) );
  OAI22_X1 U911 ( .A1(n12408), .A2(n12490), .B1(n12404), .B2(n11007), .ZN(
        n4350) );
  OAI22_X1 U912 ( .A1(n12408), .A2(n12487), .B1(n12404), .B2(n11008), .ZN(
        n4349) );
  OAI22_X1 U913 ( .A1(n12409), .A2(n12484), .B1(n12404), .B2(n11009), .ZN(
        n4348) );
  OAI22_X1 U914 ( .A1(n12409), .A2(n12481), .B1(n12404), .B2(n11010), .ZN(
        n4347) );
  OAI22_X1 U915 ( .A1(n12409), .A2(n12478), .B1(n1115), .B2(n11011), .ZN(n4346) );
  OAI22_X1 U916 ( .A1(n12409), .A2(n12475), .B1(n1115), .B2(n11012), .ZN(n4345) );
  OAI22_X1 U917 ( .A1(n12409), .A2(n12472), .B1(n1115), .B2(n11061), .ZN(n4344) );
  OAI22_X1 U918 ( .A1(n12410), .A2(n12469), .B1(n1115), .B2(n11062), .ZN(n4343) );
  OAI22_X1 U919 ( .A1(n12410), .A2(n12466), .B1(n12404), .B2(n11063), .ZN(
        n4342) );
  OAI22_X1 U920 ( .A1(n12410), .A2(n12463), .B1(n12404), .B2(n11064), .ZN(
        n4341) );
  OAI22_X1 U921 ( .A1(n12410), .A2(n12460), .B1(n12404), .B2(n11065), .ZN(
        n4340) );
  OAI22_X1 U922 ( .A1(n12410), .A2(n12457), .B1(n12404), .B2(n11066), .ZN(
        n4339) );
  OAI22_X1 U923 ( .A1(n12411), .A2(n12454), .B1(n12404), .B2(n11067), .ZN(
        n4338) );
  OAI22_X1 U924 ( .A1(n12411), .A2(n12451), .B1(n12404), .B2(n11068), .ZN(
        n4337) );
  OAI22_X1 U925 ( .A1(n12398), .A2(n12514), .B1(n12395), .B2(n11386), .ZN(
        n4326) );
  OAI22_X1 U926 ( .A1(n12398), .A2(n12511), .B1(n12395), .B2(n11391), .ZN(
        n4325) );
  OAI22_X1 U927 ( .A1(n12398), .A2(n12508), .B1(n12395), .B2(n11396), .ZN(
        n4324) );
  OAI22_X1 U928 ( .A1(n12398), .A2(n12505), .B1(n12395), .B2(n11401), .ZN(
        n4323) );
  OAI22_X1 U929 ( .A1(n12398), .A2(n12502), .B1(n12395), .B2(n11406), .ZN(
        n4322) );
  OAI22_X1 U930 ( .A1(n12399), .A2(n12499), .B1(n12395), .B2(n11411), .ZN(
        n4321) );
  OAI22_X1 U931 ( .A1(n12399), .A2(n12496), .B1(n12395), .B2(n11416), .ZN(
        n4320) );
  OAI22_X1 U932 ( .A1(n12399), .A2(n12493), .B1(n12395), .B2(n11421), .ZN(
        n4319) );
  OAI22_X1 U933 ( .A1(n12399), .A2(n12490), .B1(n12395), .B2(n11426), .ZN(
        n4318) );
  OAI22_X1 U934 ( .A1(n12399), .A2(n12487), .B1(n12395), .B2(n11431), .ZN(
        n4317) );
  OAI22_X1 U935 ( .A1(n12400), .A2(n12484), .B1(n12395), .B2(n11435), .ZN(
        n4316) );
  OAI22_X1 U936 ( .A1(n12400), .A2(n12481), .B1(n12395), .B2(n11439), .ZN(
        n4315) );
  OAI22_X1 U937 ( .A1(n12400), .A2(n12478), .B1(n1117), .B2(n11443), .ZN(n4314) );
  OAI22_X1 U938 ( .A1(n12400), .A2(n12475), .B1(n1117), .B2(n11447), .ZN(n4313) );
  OAI22_X1 U939 ( .A1(n12400), .A2(n12472), .B1(n1117), .B2(n11293), .ZN(n4312) );
  OAI22_X1 U940 ( .A1(n12401), .A2(n12469), .B1(n1117), .B2(n11295), .ZN(n4311) );
  OAI22_X1 U941 ( .A1(n12401), .A2(n12466), .B1(n12395), .B2(n11297), .ZN(
        n4310) );
  OAI22_X1 U942 ( .A1(n12401), .A2(n12463), .B1(n12395), .B2(n11299), .ZN(
        n4309) );
  OAI22_X1 U943 ( .A1(n12401), .A2(n12460), .B1(n12395), .B2(n11301), .ZN(
        n4308) );
  OAI22_X1 U944 ( .A1(n12401), .A2(n12457), .B1(n12395), .B2(n11303), .ZN(
        n4307) );
  OAI22_X1 U945 ( .A1(n12402), .A2(n12454), .B1(n12395), .B2(n11305), .ZN(
        n4306) );
  OAI22_X1 U946 ( .A1(n12402), .A2(n12451), .B1(n12395), .B2(n11307), .ZN(
        n4305) );
  OAI22_X1 U947 ( .A1(n12389), .A2(n12514), .B1(n12386), .B2(n11130), .ZN(
        n4294) );
  OAI22_X1 U948 ( .A1(n12389), .A2(n12511), .B1(n12386), .B2(n11135), .ZN(
        n4293) );
  OAI22_X1 U949 ( .A1(n12389), .A2(n12508), .B1(n12386), .B2(n11140), .ZN(
        n4292) );
  OAI22_X1 U950 ( .A1(n12389), .A2(n12505), .B1(n12386), .B2(n11145), .ZN(
        n4291) );
  OAI22_X1 U951 ( .A1(n12389), .A2(n12502), .B1(n12386), .B2(n11150), .ZN(
        n4290) );
  OAI22_X1 U952 ( .A1(n12390), .A2(n12499), .B1(n12386), .B2(n11155), .ZN(
        n4289) );
  OAI22_X1 U953 ( .A1(n12390), .A2(n12496), .B1(n12386), .B2(n11160), .ZN(
        n4288) );
  OAI22_X1 U954 ( .A1(n12390), .A2(n12493), .B1(n12386), .B2(n11165), .ZN(
        n4287) );
  OAI22_X1 U955 ( .A1(n12390), .A2(n12490), .B1(n12386), .B2(n11170), .ZN(
        n4286) );
  OAI22_X1 U956 ( .A1(n12390), .A2(n12487), .B1(n12386), .B2(n11175), .ZN(
        n4285) );
  OAI22_X1 U957 ( .A1(n12391), .A2(n12484), .B1(n12386), .B2(n11179), .ZN(
        n4284) );
  OAI22_X1 U958 ( .A1(n12391), .A2(n12481), .B1(n12386), .B2(n11183), .ZN(
        n4283) );
  OAI22_X1 U959 ( .A1(n12391), .A2(n12478), .B1(n1119), .B2(n11187), .ZN(n4282) );
  OAI22_X1 U960 ( .A1(n12391), .A2(n12475), .B1(n1119), .B2(n11191), .ZN(n4281) );
  OAI22_X1 U961 ( .A1(n12391), .A2(n12472), .B1(n1119), .B2(n11037), .ZN(n4280) );
  OAI22_X1 U962 ( .A1(n12392), .A2(n12469), .B1(n1119), .B2(n11039), .ZN(n4279) );
  OAI22_X1 U963 ( .A1(n12392), .A2(n12466), .B1(n12386), .B2(n11041), .ZN(
        n4278) );
  OAI22_X1 U964 ( .A1(n12392), .A2(n12463), .B1(n12386), .B2(n11043), .ZN(
        n4277) );
  OAI22_X1 U965 ( .A1(n12392), .A2(n12460), .B1(n12386), .B2(n11045), .ZN(
        n4276) );
  OAI22_X1 U966 ( .A1(n12392), .A2(n12457), .B1(n12386), .B2(n11047), .ZN(
        n4275) );
  OAI22_X1 U967 ( .A1(n12393), .A2(n12454), .B1(n12386), .B2(n11049), .ZN(
        n4274) );
  OAI22_X1 U968 ( .A1(n12393), .A2(n12451), .B1(n12386), .B2(n11051), .ZN(
        n4273) );
  OAI22_X1 U969 ( .A1(n12543), .A2(n12553), .B1(n12542), .B2(n11085), .ZN(
        n4528) );
  OAI22_X1 U970 ( .A1(n12543), .A2(n12541), .B1(n12542), .B2(n11089), .ZN(
        n4527) );
  OAI22_X1 U971 ( .A1(n12543), .A2(n12538), .B1(n12542), .B2(n11093), .ZN(
        n4526) );
  OAI22_X1 U972 ( .A1(n12543), .A2(n12535), .B1(n12542), .B2(n11097), .ZN(
        n4525) );
  OAI22_X1 U973 ( .A1(n12543), .A2(n12532), .B1(n1072), .B2(n11101), .ZN(n4524) );
  OAI22_X1 U974 ( .A1(n12544), .A2(n12529), .B1(n1072), .B2(n11105), .ZN(n4523) );
  OAI22_X1 U975 ( .A1(n12544), .A2(n12526), .B1(n1072), .B2(n11109), .ZN(n4522) );
  OAI22_X1 U976 ( .A1(n12544), .A2(n12523), .B1(n1072), .B2(n11113), .ZN(n4521) );
  OAI22_X1 U977 ( .A1(n12544), .A2(n12520), .B1(n1072), .B2(n11117), .ZN(n4520) );
  OAI22_X1 U978 ( .A1(n12544), .A2(n12517), .B1(n1072), .B2(n11122), .ZN(n4519) );
  OAI22_X1 U979 ( .A1(n12441), .A2(n12553), .B1(n12440), .B2(n11341), .ZN(
        n4496) );
  OAI22_X1 U980 ( .A1(n12441), .A2(n12541), .B1(n12440), .B2(n11345), .ZN(
        n4495) );
  OAI22_X1 U981 ( .A1(n12441), .A2(n12538), .B1(n12440), .B2(n11349), .ZN(
        n4494) );
  OAI22_X1 U982 ( .A1(n12441), .A2(n12535), .B1(n12440), .B2(n11353), .ZN(
        n4493) );
  OAI22_X1 U983 ( .A1(n12441), .A2(n12532), .B1(n1106), .B2(n11357), .ZN(n4492) );
  OAI22_X1 U984 ( .A1(n12442), .A2(n12529), .B1(n1106), .B2(n11361), .ZN(n4491) );
  OAI22_X1 U985 ( .A1(n12442), .A2(n12526), .B1(n1106), .B2(n11365), .ZN(n4490) );
  OAI22_X1 U986 ( .A1(n12442), .A2(n12523), .B1(n1106), .B2(n11369), .ZN(n4489) );
  OAI22_X1 U987 ( .A1(n12442), .A2(n12520), .B1(n1106), .B2(n11373), .ZN(n4488) );
  OAI22_X1 U988 ( .A1(n12442), .A2(n12517), .B1(n1106), .B2(n11378), .ZN(n4487) );
  OAI22_X1 U989 ( .A1(n12432), .A2(n12553), .B1(n12431), .B2(n11086), .ZN(
        n4464) );
  OAI22_X1 U990 ( .A1(n12432), .A2(n12541), .B1(n12431), .B2(n11090), .ZN(
        n4463) );
  OAI22_X1 U991 ( .A1(n12432), .A2(n12538), .B1(n12431), .B2(n11094), .ZN(
        n4462) );
  OAI22_X1 U992 ( .A1(n12432), .A2(n12535), .B1(n12431), .B2(n11098), .ZN(
        n4461) );
  OAI22_X1 U993 ( .A1(n12432), .A2(n12532), .B1(n1108), .B2(n11102), .ZN(n4460) );
  OAI22_X1 U994 ( .A1(n12433), .A2(n12529), .B1(n1108), .B2(n11106), .ZN(n4459) );
  OAI22_X1 U995 ( .A1(n12433), .A2(n12526), .B1(n1108), .B2(n11110), .ZN(n4458) );
  OAI22_X1 U996 ( .A1(n12433), .A2(n12523), .B1(n1108), .B2(n11114), .ZN(n4457) );
  OAI22_X1 U997 ( .A1(n12433), .A2(n12520), .B1(n1108), .B2(n10959), .ZN(n4456) );
  OAI22_X1 U998 ( .A1(n12433), .A2(n12517), .B1(n1108), .B2(n11123), .ZN(n4455) );
  OAI22_X1 U999 ( .A1(n12423), .A2(n12553), .B1(n12422), .B2(n11342), .ZN(
        n4432) );
  OAI22_X1 U1000 ( .A1(n12423), .A2(n12541), .B1(n12422), .B2(n11346), .ZN(
        n4431) );
  OAI22_X1 U1001 ( .A1(n12423), .A2(n12538), .B1(n12422), .B2(n11350), .ZN(
        n4430) );
  OAI22_X1 U1002 ( .A1(n12423), .A2(n12535), .B1(n12422), .B2(n11354), .ZN(
        n4429) );
  OAI22_X1 U1003 ( .A1(n12423), .A2(n12532), .B1(n1110), .B2(n11358), .ZN(
        n4428) );
  OAI22_X1 U1004 ( .A1(n12424), .A2(n12529), .B1(n1110), .B2(n11362), .ZN(
        n4427) );
  OAI22_X1 U1005 ( .A1(n12424), .A2(n12526), .B1(n1110), .B2(n11366), .ZN(
        n4426) );
  OAI22_X1 U1006 ( .A1(n12424), .A2(n12523), .B1(n1110), .B2(n11370), .ZN(
        n4425) );
  OAI22_X1 U1007 ( .A1(n12424), .A2(n12520), .B1(n1110), .B2(n11215), .ZN(
        n4424) );
  OAI22_X1 U1008 ( .A1(n12424), .A2(n12517), .B1(n1110), .B2(n11379), .ZN(
        n4423) );
  OAI22_X1 U1009 ( .A1(n12226), .A2(n12476), .B1(n12224), .B2(n11184), .ZN(
        n2945) );
  OAI22_X1 U1010 ( .A1(n12226), .A2(n12473), .B1(n12224), .B2(n11188), .ZN(
        n2946) );
  OAI22_X1 U1011 ( .A1(n12226), .A2(n12470), .B1(n12224), .B2(n11036), .ZN(
        n2947) );
  OAI22_X1 U1012 ( .A1(n12226), .A2(n12467), .B1(n12224), .B2(n11013), .ZN(
        n2948) );
  OAI22_X1 U1013 ( .A1(n12226), .A2(n12464), .B1(n1140), .B2(n11014), .ZN(
        n2949) );
  OAI22_X1 U1014 ( .A1(n12225), .A2(n12461), .B1(n1140), .B2(n11015), .ZN(
        n2950) );
  OAI22_X1 U1015 ( .A1(n12225), .A2(n12458), .B1(n1140), .B2(n11016), .ZN(
        n2951) );
  OAI22_X1 U1016 ( .A1(n12225), .A2(n12455), .B1(n1140), .B2(n11017), .ZN(
        n2952) );
  OAI22_X1 U1017 ( .A1(n12225), .A2(n12452), .B1(n1140), .B2(n11018), .ZN(
        n2953) );
  OAI22_X1 U1018 ( .A1(n12225), .A2(n12449), .B1(n1140), .B2(n11019), .ZN(
        n2954) );
  OAI22_X1 U1019 ( .A1(n12235), .A2(n12476), .B1(n12233), .B2(n11440), .ZN(
        n2977) );
  OAI22_X1 U1020 ( .A1(n12235), .A2(n12473), .B1(n12233), .B2(n11444), .ZN(
        n2978) );
  OAI22_X1 U1021 ( .A1(n12235), .A2(n12470), .B1(n12233), .B2(n11292), .ZN(
        n2979) );
  OAI22_X1 U1022 ( .A1(n12235), .A2(n12467), .B1(n12233), .B2(n11269), .ZN(
        n2980) );
  OAI22_X1 U1023 ( .A1(n12235), .A2(n12464), .B1(n1139), .B2(n11270), .ZN(
        n2981) );
  OAI22_X1 U1024 ( .A1(n12234), .A2(n12461), .B1(n1139), .B2(n11271), .ZN(
        n2982) );
  OAI22_X1 U1025 ( .A1(n12234), .A2(n12458), .B1(n1139), .B2(n11272), .ZN(
        n2983) );
  OAI22_X1 U1026 ( .A1(n12234), .A2(n12455), .B1(n1139), .B2(n11273), .ZN(
        n2984) );
  OAI22_X1 U1027 ( .A1(n12234), .A2(n12452), .B1(n1139), .B2(n11274), .ZN(
        n2985) );
  OAI22_X1 U1028 ( .A1(n12234), .A2(n12449), .B1(n1139), .B2(n11275), .ZN(
        n2986) );
  OAI22_X1 U1029 ( .A1(n12262), .A2(n12477), .B1(n12260), .B2(n11186), .ZN(
        n3073) );
  OAI22_X1 U1030 ( .A1(n12262), .A2(n12474), .B1(n12260), .B2(n11190), .ZN(
        n3074) );
  OAI22_X1 U1031 ( .A1(n12262), .A2(n12471), .B1(n12260), .B2(n11038), .ZN(
        n3075) );
  OAI22_X1 U1032 ( .A1(n12262), .A2(n12468), .B1(n12260), .B2(n11040), .ZN(
        n3076) );
  OAI22_X1 U1033 ( .A1(n12262), .A2(n12465), .B1(n1136), .B2(n11042), .ZN(
        n3077) );
  OAI22_X1 U1034 ( .A1(n12261), .A2(n12462), .B1(n1136), .B2(n11044), .ZN(
        n3078) );
  OAI22_X1 U1035 ( .A1(n12261), .A2(n12459), .B1(n1136), .B2(n11046), .ZN(
        n3079) );
  OAI22_X1 U1036 ( .A1(n12261), .A2(n12456), .B1(n1136), .B2(n11048), .ZN(
        n3080) );
  OAI22_X1 U1037 ( .A1(n12261), .A2(n12453), .B1(n1136), .B2(n11050), .ZN(
        n3081) );
  OAI22_X1 U1038 ( .A1(n12261), .A2(n12450), .B1(n1136), .B2(n11052), .ZN(
        n3082) );
  OAI22_X1 U1039 ( .A1(n12271), .A2(n12477), .B1(n12269), .B2(n11442), .ZN(
        n3105) );
  OAI22_X1 U1040 ( .A1(n12271), .A2(n12474), .B1(n12269), .B2(n11446), .ZN(
        n3106) );
  OAI22_X1 U1041 ( .A1(n12271), .A2(n12471), .B1(n12269), .B2(n11294), .ZN(
        n3107) );
  OAI22_X1 U1042 ( .A1(n12271), .A2(n12468), .B1(n12269), .B2(n11296), .ZN(
        n3108) );
  OAI22_X1 U1043 ( .A1(n12271), .A2(n12465), .B1(n1134), .B2(n11298), .ZN(
        n3109) );
  OAI22_X1 U1044 ( .A1(n12270), .A2(n12462), .B1(n1134), .B2(n11300), .ZN(
        n3110) );
  OAI22_X1 U1045 ( .A1(n12270), .A2(n12459), .B1(n1134), .B2(n11302), .ZN(
        n3111) );
  OAI22_X1 U1046 ( .A1(n12270), .A2(n12456), .B1(n1134), .B2(n11304), .ZN(
        n3112) );
  OAI22_X1 U1047 ( .A1(n12270), .A2(n12453), .B1(n1134), .B2(n11306), .ZN(
        n3113) );
  OAI22_X1 U1048 ( .A1(n12270), .A2(n12450), .B1(n1134), .B2(n11308), .ZN(
        n3114) );
  OAI22_X1 U1049 ( .A1(n12298), .A2(n12477), .B1(n12296), .B2(n10949), .ZN(
        n3201) );
  OAI22_X1 U1050 ( .A1(n12298), .A2(n12474), .B1(n12296), .B2(n10950), .ZN(
        n3202) );
  OAI22_X1 U1051 ( .A1(n12298), .A2(n12471), .B1(n12296), .B2(n11069), .ZN(
        n3203) );
  OAI22_X1 U1052 ( .A1(n12298), .A2(n12468), .B1(n12296), .B2(n11071), .ZN(
        n3204) );
  OAI22_X1 U1053 ( .A1(n12298), .A2(n12465), .B1(n1131), .B2(n11073), .ZN(
        n3205) );
  OAI22_X1 U1054 ( .A1(n12297), .A2(n12462), .B1(n1131), .B2(n11075), .ZN(
        n3206) );
  OAI22_X1 U1055 ( .A1(n12297), .A2(n12459), .B1(n1131), .B2(n11077), .ZN(
        n3207) );
  OAI22_X1 U1056 ( .A1(n12297), .A2(n12456), .B1(n1131), .B2(n11079), .ZN(
        n3208) );
  OAI22_X1 U1057 ( .A1(n12297), .A2(n12453), .B1(n1131), .B2(n11081), .ZN(
        n3209) );
  OAI22_X1 U1058 ( .A1(n12297), .A2(n12450), .B1(n1131), .B2(n11083), .ZN(
        n3210) );
  OAI22_X1 U1059 ( .A1(n12307), .A2(n12477), .B1(n12305), .B2(n11205), .ZN(
        n3233) );
  OAI22_X1 U1060 ( .A1(n12307), .A2(n12474), .B1(n12305), .B2(n11206), .ZN(
        n3234) );
  OAI22_X1 U1061 ( .A1(n12307), .A2(n12471), .B1(n12305), .B2(n11325), .ZN(
        n3235) );
  OAI22_X1 U1062 ( .A1(n12307), .A2(n12468), .B1(n12305), .B2(n11327), .ZN(
        n3236) );
  OAI22_X1 U1063 ( .A1(n12307), .A2(n12465), .B1(n1130), .B2(n11329), .ZN(
        n3237) );
  OAI22_X1 U1064 ( .A1(n12306), .A2(n12462), .B1(n1130), .B2(n11331), .ZN(
        n3238) );
  OAI22_X1 U1065 ( .A1(n12306), .A2(n12459), .B1(n1130), .B2(n11333), .ZN(
        n3239) );
  OAI22_X1 U1066 ( .A1(n12306), .A2(n12456), .B1(n1130), .B2(n11335), .ZN(
        n3240) );
  OAI22_X1 U1067 ( .A1(n12306), .A2(n12453), .B1(n1130), .B2(n11337), .ZN(
        n3241) );
  OAI22_X1 U1068 ( .A1(n12306), .A2(n12450), .B1(n1130), .B2(n11339), .ZN(
        n3242) );
  OAI22_X1 U1069 ( .A1(n12334), .A2(n12477), .B1(n12332), .B2(n10974), .ZN(
        n3329) );
  OAI22_X1 U1070 ( .A1(n12334), .A2(n12474), .B1(n12332), .B2(n10975), .ZN(
        n3330) );
  OAI22_X1 U1071 ( .A1(n12334), .A2(n12471), .B1(n12332), .B2(n11053), .ZN(
        n3331) );
  OAI22_X1 U1072 ( .A1(n12334), .A2(n12468), .B1(n12332), .B2(n11054), .ZN(
        n3332) );
  OAI22_X1 U1073 ( .A1(n12334), .A2(n12465), .B1(n1127), .B2(n11055), .ZN(
        n3333) );
  OAI22_X1 U1074 ( .A1(n12333), .A2(n12462), .B1(n1127), .B2(n11056), .ZN(
        n3334) );
  OAI22_X1 U1075 ( .A1(n12333), .A2(n12459), .B1(n1127), .B2(n11057), .ZN(
        n3335) );
  OAI22_X1 U1076 ( .A1(n12333), .A2(n12456), .B1(n1127), .B2(n11058), .ZN(
        n3336) );
  OAI22_X1 U1077 ( .A1(n12333), .A2(n12453), .B1(n1127), .B2(n11059), .ZN(
        n3337) );
  OAI22_X1 U1078 ( .A1(n12333), .A2(n12450), .B1(n1127), .B2(n11060), .ZN(
        n3338) );
  OAI22_X1 U1079 ( .A1(n12343), .A2(n12477), .B1(n12341), .B2(n11230), .ZN(
        n3361) );
  OAI22_X1 U1080 ( .A1(n12343), .A2(n12474), .B1(n12341), .B2(n11231), .ZN(
        n3362) );
  OAI22_X1 U1081 ( .A1(n12343), .A2(n12471), .B1(n12341), .B2(n11309), .ZN(
        n3363) );
  OAI22_X1 U1082 ( .A1(n12343), .A2(n12468), .B1(n12341), .B2(n11310), .ZN(
        n3364) );
  OAI22_X1 U1083 ( .A1(n12343), .A2(n12465), .B1(n1125), .B2(n11311), .ZN(
        n3365) );
  OAI22_X1 U1084 ( .A1(n12342), .A2(n12462), .B1(n1125), .B2(n11312), .ZN(
        n3366) );
  OAI22_X1 U1085 ( .A1(n12342), .A2(n12459), .B1(n1125), .B2(n11313), .ZN(
        n3367) );
  OAI22_X1 U1086 ( .A1(n12342), .A2(n12456), .B1(n1125), .B2(n11314), .ZN(
        n3368) );
  OAI22_X1 U1087 ( .A1(n12342), .A2(n12453), .B1(n1125), .B2(n11315), .ZN(
        n3369) );
  OAI22_X1 U1088 ( .A1(n12342), .A2(n12450), .B1(n1125), .B2(n11316), .ZN(
        n3370) );
  OAI22_X1 U1089 ( .A1(n12414), .A2(n12553), .B1(n12413), .B2(n11277), .ZN(
        n4400) );
  OAI22_X1 U1090 ( .A1(n12414), .A2(n12541), .B1(n12413), .B2(n11279), .ZN(
        n4399) );
  OAI22_X1 U1091 ( .A1(n12414), .A2(n12538), .B1(n12413), .B2(n11281), .ZN(
        n4398) );
  OAI22_X1 U1092 ( .A1(n12414), .A2(n12535), .B1(n12413), .B2(n11283), .ZN(
        n4397) );
  OAI22_X1 U1093 ( .A1(n12414), .A2(n12532), .B1(n1112), .B2(n11285), .ZN(
        n4396) );
  OAI22_X1 U1094 ( .A1(n12415), .A2(n12529), .B1(n1112), .B2(n11287), .ZN(
        n4395) );
  OAI22_X1 U1095 ( .A1(n12415), .A2(n12526), .B1(n1112), .B2(n11289), .ZN(
        n4394) );
  OAI22_X1 U1096 ( .A1(n12415), .A2(n12523), .B1(n1112), .B2(n11291), .ZN(
        n4393) );
  OAI22_X1 U1097 ( .A1(n12415), .A2(n12520), .B1(n1112), .B2(n11253), .ZN(
        n4392) );
  OAI22_X1 U1098 ( .A1(n12415), .A2(n12517), .B1(n1112), .B2(n11254), .ZN(
        n4391) );
  OAI22_X1 U1099 ( .A1(n12405), .A2(n12553), .B1(n12404), .B2(n11021), .ZN(
        n4368) );
  OAI22_X1 U1100 ( .A1(n12405), .A2(n12541), .B1(n12404), .B2(n11023), .ZN(
        n4367) );
  OAI22_X1 U1101 ( .A1(n12405), .A2(n12538), .B1(n12404), .B2(n11025), .ZN(
        n4366) );
  OAI22_X1 U1102 ( .A1(n12405), .A2(n12535), .B1(n12404), .B2(n11027), .ZN(
        n4365) );
  OAI22_X1 U1103 ( .A1(n12405), .A2(n12532), .B1(n1115), .B2(n11029), .ZN(
        n4364) );
  OAI22_X1 U1104 ( .A1(n12406), .A2(n12529), .B1(n1115), .B2(n11031), .ZN(
        n4363) );
  OAI22_X1 U1105 ( .A1(n12406), .A2(n12526), .B1(n1115), .B2(n11033), .ZN(
        n4362) );
  OAI22_X1 U1106 ( .A1(n12406), .A2(n12523), .B1(n1115), .B2(n11035), .ZN(
        n4361) );
  OAI22_X1 U1107 ( .A1(n12406), .A2(n12520), .B1(n1115), .B2(n10997), .ZN(
        n4360) );
  OAI22_X1 U1108 ( .A1(n12406), .A2(n12517), .B1(n1115), .B2(n10998), .ZN(
        n4359) );
  OAI22_X1 U1109 ( .A1(n12396), .A2(n12553), .B1(n12395), .B2(n11344), .ZN(
        n4336) );
  OAI22_X1 U1110 ( .A1(n12396), .A2(n12541), .B1(n12395), .B2(n11348), .ZN(
        n4335) );
  OAI22_X1 U1111 ( .A1(n12396), .A2(n12538), .B1(n12395), .B2(n11352), .ZN(
        n4334) );
  OAI22_X1 U1112 ( .A1(n12396), .A2(n12535), .B1(n12395), .B2(n11356), .ZN(
        n4333) );
  OAI22_X1 U1113 ( .A1(n12396), .A2(n12532), .B1(n1117), .B2(n11360), .ZN(
        n4332) );
  OAI22_X1 U1114 ( .A1(n12397), .A2(n12529), .B1(n1117), .B2(n11364), .ZN(
        n4331) );
  OAI22_X1 U1115 ( .A1(n12397), .A2(n12526), .B1(n1117), .B2(n11368), .ZN(
        n4330) );
  OAI22_X1 U1116 ( .A1(n12397), .A2(n12523), .B1(n1117), .B2(n11372), .ZN(
        n4329) );
  OAI22_X1 U1117 ( .A1(n12397), .A2(n12520), .B1(n1117), .B2(n11376), .ZN(
        n4328) );
  OAI22_X1 U1118 ( .A1(n12397), .A2(n12517), .B1(n1117), .B2(n11381), .ZN(
        n4327) );
  OAI22_X1 U1119 ( .A1(n12387), .A2(n12553), .B1(n12386), .B2(n11088), .ZN(
        n4304) );
  OAI22_X1 U1120 ( .A1(n12387), .A2(n12541), .B1(n12386), .B2(n11092), .ZN(
        n4303) );
  OAI22_X1 U1121 ( .A1(n12387), .A2(n12538), .B1(n12386), .B2(n11096), .ZN(
        n4302) );
  OAI22_X1 U1122 ( .A1(n12387), .A2(n12535), .B1(n12386), .B2(n11100), .ZN(
        n4301) );
  OAI22_X1 U1123 ( .A1(n12387), .A2(n12532), .B1(n1119), .B2(n11104), .ZN(
        n4300) );
  OAI22_X1 U1124 ( .A1(n12388), .A2(n12529), .B1(n1119), .B2(n11108), .ZN(
        n4299) );
  OAI22_X1 U1125 ( .A1(n12388), .A2(n12526), .B1(n1119), .B2(n11112), .ZN(
        n4298) );
  OAI22_X1 U1126 ( .A1(n12388), .A2(n12523), .B1(n1119), .B2(n11116), .ZN(
        n4297) );
  OAI22_X1 U1127 ( .A1(n12388), .A2(n12520), .B1(n1119), .B2(n11120), .ZN(
        n4296) );
  OAI22_X1 U1128 ( .A1(n12388), .A2(n12517), .B1(n1119), .B2(n11125), .ZN(
        n4295) );
  NAND2_X1 U1129 ( .A1(n12561), .A2(n12059), .ZN(n1810) );
  INV_X1 U1130 ( .A(n2437), .ZN(n12561) );
  INV_X1 U1131 ( .A(n1112), .ZN(n12421) );
  OAI21_X1 U1132 ( .B1(n1113), .B2(n1114), .A(n12558), .ZN(n1112) );
  INV_X1 U1133 ( .A(n1115), .ZN(n12412) );
  OAI21_X1 U1134 ( .B1(n1113), .B2(n1116), .A(n12558), .ZN(n1115) );
  INV_X1 U1135 ( .A(n1117), .ZN(n12403) );
  OAI21_X1 U1136 ( .B1(n1113), .B2(n1118), .A(n12558), .ZN(n1117) );
  INV_X1 U1137 ( .A(n1119), .ZN(n12394) );
  OAI21_X1 U1138 ( .B1(n1113), .B2(n1120), .A(n12558), .ZN(n1119) );
  INV_X1 U1139 ( .A(n1146), .ZN(n12178) );
  OAI21_X1 U1140 ( .B1(n1105), .B2(n1114), .A(n12556), .ZN(n1146) );
  INV_X1 U1141 ( .A(n1145), .ZN(n12187) );
  OAI21_X1 U1142 ( .B1(n1105), .B2(n1116), .A(n12556), .ZN(n1145) );
  INV_X1 U1143 ( .A(n1106), .ZN(n12448) );
  OAI21_X1 U1144 ( .B1(n1105), .B2(n1107), .A(n12559), .ZN(n1106) );
  INV_X1 U1145 ( .A(n1144), .ZN(n12196) );
  OAI21_X1 U1146 ( .B1(n1105), .B2(n1118), .A(n12556), .ZN(n1144) );
  INV_X1 U1147 ( .A(n1143), .ZN(n12205) );
  OAI21_X1 U1148 ( .B1(n1105), .B2(n1120), .A(n12556), .ZN(n1143) );
  INV_X1 U1149 ( .A(n1108), .ZN(n12439) );
  OAI21_X1 U1150 ( .B1(n1105), .B2(n1109), .A(n12559), .ZN(n1108) );
  INV_X1 U1151 ( .A(n1110), .ZN(n12430) );
  OAI21_X1 U1152 ( .B1(n1105), .B2(n1111), .A(n12559), .ZN(n1110) );
  INV_X1 U1153 ( .A(n1124), .ZN(n12358) );
  OAI21_X1 U1154 ( .B1(n1104), .B2(n1113), .A(n12558), .ZN(n1124) );
  INV_X1 U1155 ( .A(n1123), .ZN(n12367) );
  OAI21_X1 U1156 ( .B1(n1107), .B2(n1113), .A(n12558), .ZN(n1123) );
  INV_X1 U1157 ( .A(n1122), .ZN(n12376) );
  OAI21_X1 U1158 ( .B1(n1109), .B2(n1113), .A(n12558), .ZN(n1122) );
  INV_X1 U1159 ( .A(n1121), .ZN(n12385) );
  OAI21_X1 U1160 ( .B1(n1111), .B2(n1113), .A(n12558), .ZN(n1121) );
  INV_X1 U1161 ( .A(n1072), .ZN(n12550) );
  OAI21_X1 U1162 ( .B1(n1104), .B2(n1105), .A(n12559), .ZN(n1072) );
  AND3_X1 U1163 ( .A1(n2437), .A2(n12061), .A3(n12559), .ZN(n1815) );
  NAND2_X1 U1164 ( .A1(DATAIN[27]), .A2(n12554), .ZN(n1099) );
  NAND2_X1 U1165 ( .A1(DATAIN[28]), .A2(n12554), .ZN(n1100) );
  NAND2_X1 U1166 ( .A1(DATAIN[31]), .A2(n12554), .ZN(n1103) );
  NAND2_X1 U1167 ( .A1(DATAIN[13]), .A2(n12555), .ZN(n1085) );
  NAND2_X1 U1168 ( .A1(DATAIN[15]), .A2(n12555), .ZN(n1087) );
  BUF_X1 U1169 ( .A(n1071), .Z(n12553) );
  BUF_X1 U1170 ( .A(n1081), .Z(n12517) );
  BUF_X1 U1171 ( .A(n1082), .Z(n12514) );
  BUF_X1 U1172 ( .A(n1089), .Z(n12493) );
  BUF_X1 U1173 ( .A(n1092), .Z(n12484) );
  BUF_X1 U1174 ( .A(n1096), .Z(n12472) );
  BUF_X1 U1175 ( .A(n1073), .Z(n12541) );
  BUF_X1 U1176 ( .A(n1075), .Z(n12535) );
  BUF_X1 U1177 ( .A(n1811), .Z(n12061) );
  BUF_X1 U1178 ( .A(n1148), .Z(n12166) );
  BUF_X1 U1179 ( .A(n1071), .Z(n12551) );
  BUF_X1 U1180 ( .A(n1081), .Z(n12515) );
  BUF_X1 U1181 ( .A(n1082), .Z(n12512) );
  BUF_X1 U1182 ( .A(n1089), .Z(n12491) );
  BUF_X1 U1183 ( .A(n1092), .Z(n12482) );
  BUF_X1 U1184 ( .A(n1096), .Z(n12470) );
  BUF_X1 U1185 ( .A(n1073), .Z(n12539) );
  BUF_X1 U1186 ( .A(n1075), .Z(n12533) );
  BUF_X1 U1187 ( .A(n1071), .Z(n12552) );
  BUF_X1 U1188 ( .A(n1081), .Z(n12516) );
  BUF_X1 U1189 ( .A(n1082), .Z(n12513) );
  BUF_X1 U1190 ( .A(n1089), .Z(n12492) );
  BUF_X1 U1191 ( .A(n1092), .Z(n12483) );
  BUF_X1 U1192 ( .A(n1096), .Z(n12471) );
  BUF_X1 U1193 ( .A(n1073), .Z(n12540) );
  BUF_X1 U1194 ( .A(n1075), .Z(n12534) );
  BUF_X1 U1195 ( .A(n1811), .Z(n12059) );
  BUF_X1 U1196 ( .A(n1148), .Z(n12164) );
  BUF_X1 U1197 ( .A(n1811), .Z(n12060) );
  BUF_X1 U1198 ( .A(n1148), .Z(n12165) );
  NAND2_X1 U1199 ( .A1(n1785), .A2(n1796), .ZN(n1190) );
  NAND2_X1 U1200 ( .A1(n1785), .A2(n1797), .ZN(n1189) );
  NAND2_X1 U1201 ( .A1(n1797), .A2(n1781), .ZN(n1184) );
  NAND2_X1 U1202 ( .A1(n1800), .A2(n1783), .ZN(n1195) );
  NAND2_X1 U1203 ( .A1(n1801), .A2(n1783), .ZN(n1194) );
  NAND2_X1 U1204 ( .A1(n1800), .A2(n1786), .ZN(n1200) );
  NAND2_X1 U1205 ( .A1(n1801), .A2(n1786), .ZN(n1199) );
  NAND2_X1 U1206 ( .A1(n1780), .A2(n1785), .ZN(n1166) );
  NAND2_X1 U1207 ( .A1(n1782), .A2(n1785), .ZN(n1165) );
  NAND2_X1 U1208 ( .A1(n1788), .A2(n1785), .ZN(n1176) );
  NAND2_X1 U1209 ( .A1(n1789), .A2(n1785), .ZN(n1175) );
  NAND2_X1 U1210 ( .A1(n1781), .A2(n1796), .ZN(n1185) );
  NAND2_X1 U1211 ( .A1(n1788), .A2(n1781), .ZN(n1171) );
  NAND2_X1 U1212 ( .A1(n1789), .A2(n1781), .ZN(n1170) );
  NAND2_X1 U1213 ( .A1(n1780), .A2(n1781), .ZN(n1161) );
  NAND2_X1 U1214 ( .A1(n1782), .A2(n1781), .ZN(n1160) );
  NAND2_X1 U1215 ( .A1(n12562), .A2(n12164), .ZN(n1147) );
  INV_X1 U1216 ( .A(n1774), .ZN(n12562) );
  AND3_X1 U1217 ( .A1(n1774), .A2(n12166), .A3(n12559), .ZN(n1152) );
  AND2_X1 U1218 ( .A1(n1786), .A2(n1797), .ZN(n1186) );
  AND2_X1 U1219 ( .A1(n1786), .A2(n1796), .ZN(n1187) );
  AND2_X1 U1220 ( .A1(n1801), .A2(n1781), .ZN(n1191) );
  AND2_X1 U1221 ( .A1(n1800), .A2(n1781), .ZN(n1192) );
  AND2_X1 U1222 ( .A1(n1801), .A2(n1785), .ZN(n1196) );
  AND2_X1 U1223 ( .A1(n1800), .A2(n1785), .ZN(n1197) );
  AND2_X1 U1224 ( .A1(n1780), .A2(n1786), .ZN(n1163) );
  AND2_X1 U1225 ( .A1(n1782), .A2(n1786), .ZN(n1162) );
  AND2_X1 U1226 ( .A1(n1789), .A2(n1786), .ZN(n1172) );
  AND2_X1 U1227 ( .A1(n1788), .A2(n1786), .ZN(n1173) );
  AND2_X1 U1228 ( .A1(n1783), .A2(n1796), .ZN(n1182) );
  AND2_X1 U1229 ( .A1(n1783), .A2(n1797), .ZN(n1181) );
  AND2_X1 U1230 ( .A1(n1789), .A2(n1783), .ZN(n1167) );
  AND2_X1 U1231 ( .A1(n1788), .A2(n1783), .ZN(n1168) );
  AND2_X1 U1232 ( .A1(n1780), .A2(n1783), .ZN(n1158) );
  AND2_X1 U1233 ( .A1(n1782), .A2(n1783), .ZN(n1157) );
  NAND2_X1 U1234 ( .A1(DATAIN[4]), .A2(n12556), .ZN(n1076) );
  NAND2_X1 U1235 ( .A1(DATAIN[5]), .A2(n12556), .ZN(n1077) );
  NAND2_X1 U1236 ( .A1(DATAIN[6]), .A2(n12556), .ZN(n1078) );
  NAND2_X1 U1237 ( .A1(DATAIN[7]), .A2(n12556), .ZN(n1079) );
  NAND2_X1 U1238 ( .A1(DATAIN[8]), .A2(n12556), .ZN(n1080) );
  NAND2_X1 U1239 ( .A1(DATAIN[11]), .A2(n12555), .ZN(n1083) );
  NAND2_X1 U1240 ( .A1(DATAIN[12]), .A2(n12555), .ZN(n1084) );
  NAND2_X1 U1241 ( .A1(DATAIN[16]), .A2(n12555), .ZN(n1088) );
  NAND2_X1 U1242 ( .A1(DATAIN[18]), .A2(n12555), .ZN(n1090) );
  NAND2_X1 U1243 ( .A1(DATAIN[19]), .A2(n12555), .ZN(n1091) );
  NAND2_X1 U1244 ( .A1(DATAIN[21]), .A2(n12554), .ZN(n1093) );
  NAND2_X1 U1245 ( .A1(DATAIN[22]), .A2(n12554), .ZN(n1094) );
  NAND2_X1 U1246 ( .A1(DATAIN[2]), .A2(n12556), .ZN(n1074) );
  NAND4_X1 U1247 ( .A1(WR), .A2(EN), .A3(ADD_WR[4]), .A4(n12560), .ZN(n1135)
         );
  NAND4_X1 U1248 ( .A1(WR), .A2(EN), .A3(ADD_WR[3]), .A4(n12566), .ZN(n1126)
         );
  NAND4_X1 U1249 ( .A1(WR), .A2(EN), .A3(n12560), .A4(n12566), .ZN(n1113) );
  NAND4_X1 U1250 ( .A1(WR), .A2(EN), .A3(ADD_WR[4]), .A4(ADD_WR[3]), .ZN(n1105) );
  AOI221_X1 U1251 ( .B1(n12041), .B2(n8436), .C1(n12038), .C2(n7980), .A(n2290), .ZN(n2287) );
  OAI22_X1 U1252 ( .A1(n10959), .A2(n12035), .B1(n11215), .B2(n12032), .ZN(
        n2290) );
  AOI221_X1 U1253 ( .B1(n12041), .B2(n8438), .C1(n12038), .C2(n7982), .A(n2271), .ZN(n2268) );
  OAI22_X1 U1254 ( .A1(n11123), .A2(n12035), .B1(n11379), .B2(n12032), .ZN(
        n2271) );
  AOI221_X1 U1255 ( .B1(n12041), .B2(n8440), .C1(n12038), .C2(n7984), .A(n2252), .ZN(n2249) );
  OAI22_X1 U1256 ( .A1(n11128), .A2(n12035), .B1(n11384), .B2(n12032), .ZN(
        n2252) );
  AOI221_X1 U1257 ( .B1(n12042), .B2(n8442), .C1(n12039), .C2(n7986), .A(n2233), .ZN(n2230) );
  OAI22_X1 U1258 ( .A1(n11133), .A2(n12035), .B1(n11389), .B2(n12032), .ZN(
        n2233) );
  AOI221_X1 U1259 ( .B1(n12042), .B2(n8444), .C1(n12039), .C2(n7988), .A(n2214), .ZN(n2211) );
  OAI22_X1 U1260 ( .A1(n11138), .A2(n12036), .B1(n11394), .B2(n12033), .ZN(
        n2214) );
  AOI221_X1 U1261 ( .B1(n12042), .B2(n8446), .C1(n12039), .C2(n7990), .A(n2195), .ZN(n2192) );
  OAI22_X1 U1262 ( .A1(n11143), .A2(n12036), .B1(n11399), .B2(n12033), .ZN(
        n2195) );
  AOI221_X1 U1263 ( .B1(n12042), .B2(n8448), .C1(n12039), .C2(n7992), .A(n2176), .ZN(n2173) );
  OAI22_X1 U1264 ( .A1(n11148), .A2(n12036), .B1(n11404), .B2(n12033), .ZN(
        n2176) );
  AOI221_X1 U1265 ( .B1(n12042), .B2(n8450), .C1(n12039), .C2(n7994), .A(n2157), .ZN(n2154) );
  OAI22_X1 U1266 ( .A1(n11153), .A2(n12036), .B1(n11409), .B2(n12033), .ZN(
        n2157) );
  AOI221_X1 U1267 ( .B1(n12042), .B2(n8452), .C1(n12039), .C2(n7996), .A(n2138), .ZN(n2135) );
  OAI22_X1 U1268 ( .A1(n11158), .A2(n12036), .B1(n11414), .B2(n12033), .ZN(
        n2138) );
  AOI221_X1 U1269 ( .B1(n12042), .B2(n8454), .C1(n12039), .C2(n7998), .A(n2119), .ZN(n2116) );
  OAI22_X1 U1270 ( .A1(n11163), .A2(n12036), .B1(n11419), .B2(n12033), .ZN(
        n2119) );
  AOI221_X1 U1271 ( .B1(n12042), .B2(n8456), .C1(n12039), .C2(n8000), .A(n2100), .ZN(n2097) );
  OAI22_X1 U1272 ( .A1(n11168), .A2(n12036), .B1(n11424), .B2(n12033), .ZN(
        n2100) );
  AOI221_X1 U1273 ( .B1(n12042), .B2(n8458), .C1(n12039), .C2(n8002), .A(n2081), .ZN(n2078) );
  OAI22_X1 U1274 ( .A1(n11173), .A2(n12036), .B1(n11429), .B2(n12033), .ZN(
        n2081) );
  AOI221_X1 U1275 ( .B1(n12041), .B2(n11488), .C1(n12038), .C2(n7964), .A(
        n2447), .ZN(n2440) );
  OAI22_X1 U1276 ( .A1(n11086), .A2(n12035), .B1(n11342), .B2(n12032), .ZN(
        n2447) );
  AOI221_X1 U1277 ( .B1(n12041), .B2(n11492), .C1(n12038), .C2(n7966), .A(
        n2423), .ZN(n2420) );
  OAI22_X1 U1278 ( .A1(n11090), .A2(n12035), .B1(n11346), .B2(n12032), .ZN(
        n2423) );
  AOI221_X1 U1279 ( .B1(n12041), .B2(n11496), .C1(n12038), .C2(n7968), .A(
        n2404), .ZN(n2401) );
  OAI22_X1 U1280 ( .A1(n11094), .A2(n12035), .B1(n11350), .B2(n12032), .ZN(
        n2404) );
  AOI221_X1 U1281 ( .B1(n12041), .B2(n11500), .C1(n12038), .C2(n7970), .A(
        n2385), .ZN(n2382) );
  OAI22_X1 U1282 ( .A1(n11098), .A2(n12035), .B1(n11354), .B2(n12032), .ZN(
        n2385) );
  AOI221_X1 U1283 ( .B1(n12041), .B2(n11504), .C1(n12038), .C2(n7972), .A(
        n2366), .ZN(n2363) );
  OAI22_X1 U1284 ( .A1(n11102), .A2(n12035), .B1(n11358), .B2(n12032), .ZN(
        n2366) );
  AOI221_X1 U1285 ( .B1(n12041), .B2(n11508), .C1(n12038), .C2(n7974), .A(
        n2347), .ZN(n2344) );
  OAI22_X1 U1286 ( .A1(n11106), .A2(n12035), .B1(n11362), .B2(n12032), .ZN(
        n2347) );
  AOI221_X1 U1287 ( .B1(n12041), .B2(n11512), .C1(n12038), .C2(n7976), .A(
        n2328), .ZN(n2325) );
  OAI22_X1 U1288 ( .A1(n11110), .A2(n12035), .B1(n11366), .B2(n12032), .ZN(
        n2328) );
  AOI221_X1 U1289 ( .B1(n12041), .B2(n11516), .C1(n12038), .C2(n7978), .A(
        n2309), .ZN(n2306) );
  OAI22_X1 U1290 ( .A1(n11114), .A2(n12035), .B1(n11370), .B2(n12032), .ZN(
        n2309) );
  AOI221_X1 U1291 ( .B1(n12042), .B2(n11464), .C1(n12039), .C2(n8004), .A(
        n2062), .ZN(n2059) );
  OAI22_X1 U1292 ( .A1(n10991), .A2(n12036), .B1(n11247), .B2(n12033), .ZN(
        n2062) );
  AOI221_X1 U1293 ( .B1(n12042), .B2(n11465), .C1(n12039), .C2(n8006), .A(
        n2043), .ZN(n2040) );
  OAI22_X1 U1294 ( .A1(n10992), .A2(n12036), .B1(n11248), .B2(n12033), .ZN(
        n2043) );
  AOI221_X1 U1295 ( .B1(n12043), .B2(n11466), .C1(n12040), .C2(n8008), .A(
        n2024), .ZN(n2021) );
  OAI22_X1 U1296 ( .A1(n10993), .A2(n12036), .B1(n11249), .B2(n12033), .ZN(
        n2024) );
  AOI221_X1 U1297 ( .B1(n12043), .B2(n11467), .C1(n12040), .C2(n8010), .A(
        n2005), .ZN(n2002) );
  OAI22_X1 U1298 ( .A1(n10994), .A2(n12036), .B1(n11250), .B2(n12033), .ZN(
        n2005) );
  AOI221_X1 U1299 ( .B1(n12029), .B2(n8538), .C1(n12026), .C2(n8082), .A(n2291), .ZN(n2286) );
  OAI22_X1 U1300 ( .A1(n10996), .A2(n12023), .B1(n11252), .B2(n12020), .ZN(
        n2291) );
  AOI221_X1 U1301 ( .B1(n11981), .B2(n8478), .C1(n11978), .C2(n8022), .A(n2299), .ZN(n2294) );
  OAI22_X1 U1302 ( .A1(n10997), .A2(n11975), .B1(n11253), .B2(n11972), .ZN(
        n2299) );
  AOI221_X1 U1303 ( .B1(n12029), .B2(n8540), .C1(n12026), .C2(n8084), .A(n2272), .ZN(n2267) );
  OAI22_X1 U1304 ( .A1(n11121), .A2(n12023), .B1(n11377), .B2(n12020), .ZN(
        n2272) );
  AOI221_X1 U1305 ( .B1(n11981), .B2(n8479), .C1(n11978), .C2(n8023), .A(n2280), .ZN(n2275) );
  OAI22_X1 U1306 ( .A1(n10998), .A2(n11975), .B1(n11254), .B2(n11972), .ZN(
        n2280) );
  AOI221_X1 U1307 ( .B1(n12029), .B2(n8542), .C1(n12026), .C2(n8086), .A(n2253), .ZN(n2248) );
  OAI22_X1 U1308 ( .A1(n11126), .A2(n12023), .B1(n11382), .B2(n12020), .ZN(
        n2253) );
  AOI221_X1 U1309 ( .B1(n11981), .B2(n8480), .C1(n11978), .C2(n8024), .A(n2261), .ZN(n2256) );
  OAI22_X1 U1310 ( .A1(n10999), .A2(n11975), .B1(n11255), .B2(n11972), .ZN(
        n2261) );
  AOI221_X1 U1311 ( .B1(n12030), .B2(n8544), .C1(n12027), .C2(n8088), .A(n2234), .ZN(n2229) );
  OAI22_X1 U1312 ( .A1(n11131), .A2(n12023), .B1(n11387), .B2(n12020), .ZN(
        n2234) );
  AOI221_X1 U1313 ( .B1(n11982), .B2(n8481), .C1(n11979), .C2(n8025), .A(n2242), .ZN(n2237) );
  OAI22_X1 U1314 ( .A1(n11000), .A2(n11975), .B1(n11256), .B2(n11972), .ZN(
        n2242) );
  AOI221_X1 U1315 ( .B1(n12030), .B2(n8546), .C1(n12027), .C2(n8090), .A(n2215), .ZN(n2210) );
  OAI22_X1 U1316 ( .A1(n11136), .A2(n12024), .B1(n11392), .B2(n12021), .ZN(
        n2215) );
  AOI221_X1 U1317 ( .B1(n11982), .B2(n8482), .C1(n11979), .C2(n8026), .A(n2223), .ZN(n2218) );
  OAI22_X1 U1318 ( .A1(n11001), .A2(n11976), .B1(n11257), .B2(n11973), .ZN(
        n2223) );
  AOI221_X1 U1319 ( .B1(n12030), .B2(n8548), .C1(n12027), .C2(n8092), .A(n2196), .ZN(n2191) );
  OAI22_X1 U1320 ( .A1(n11141), .A2(n12024), .B1(n11397), .B2(n12021), .ZN(
        n2196) );
  AOI221_X1 U1321 ( .B1(n11982), .B2(n8483), .C1(n11979), .C2(n8027), .A(n2204), .ZN(n2199) );
  OAI22_X1 U1322 ( .A1(n11002), .A2(n11976), .B1(n11258), .B2(n11973), .ZN(
        n2204) );
  AOI221_X1 U1323 ( .B1(n12030), .B2(n8550), .C1(n12027), .C2(n8094), .A(n2177), .ZN(n2172) );
  OAI22_X1 U1324 ( .A1(n11146), .A2(n12024), .B1(n11402), .B2(n12021), .ZN(
        n2177) );
  AOI221_X1 U1325 ( .B1(n11982), .B2(n8484), .C1(n11979), .C2(n8028), .A(n2185), .ZN(n2180) );
  OAI22_X1 U1326 ( .A1(n11003), .A2(n11976), .B1(n11259), .B2(n11973), .ZN(
        n2185) );
  AOI221_X1 U1327 ( .B1(n12030), .B2(n8552), .C1(n12027), .C2(n8096), .A(n2158), .ZN(n2153) );
  OAI22_X1 U1328 ( .A1(n11151), .A2(n12024), .B1(n11407), .B2(n12021), .ZN(
        n2158) );
  AOI221_X1 U1329 ( .B1(n11982), .B2(n8485), .C1(n11979), .C2(n8029), .A(n2166), .ZN(n2161) );
  OAI22_X1 U1330 ( .A1(n11004), .A2(n11976), .B1(n11260), .B2(n11973), .ZN(
        n2166) );
  AOI221_X1 U1331 ( .B1(n12030), .B2(n8554), .C1(n12027), .C2(n8098), .A(n2139), .ZN(n2134) );
  OAI22_X1 U1332 ( .A1(n11156), .A2(n12024), .B1(n11412), .B2(n12021), .ZN(
        n2139) );
  AOI221_X1 U1333 ( .B1(n11982), .B2(n8486), .C1(n11979), .C2(n8030), .A(n2147), .ZN(n2142) );
  OAI22_X1 U1334 ( .A1(n11005), .A2(n11976), .B1(n11261), .B2(n11973), .ZN(
        n2147) );
  AOI221_X1 U1335 ( .B1(n12030), .B2(n8556), .C1(n12027), .C2(n8100), .A(n2120), .ZN(n2115) );
  OAI22_X1 U1336 ( .A1(n11161), .A2(n12024), .B1(n11417), .B2(n12021), .ZN(
        n2120) );
  AOI221_X1 U1337 ( .B1(n11982), .B2(n8487), .C1(n11979), .C2(n8031), .A(n2128), .ZN(n2123) );
  OAI22_X1 U1338 ( .A1(n11006), .A2(n11976), .B1(n11262), .B2(n11973), .ZN(
        n2128) );
  AOI221_X1 U1339 ( .B1(n12030), .B2(n8558), .C1(n12027), .C2(n8102), .A(n2101), .ZN(n2096) );
  OAI22_X1 U1340 ( .A1(n11166), .A2(n12024), .B1(n11422), .B2(n12021), .ZN(
        n2101) );
  AOI221_X1 U1341 ( .B1(n11982), .B2(n8488), .C1(n11979), .C2(n8032), .A(n2109), .ZN(n2104) );
  OAI22_X1 U1342 ( .A1(n11007), .A2(n11976), .B1(n11263), .B2(n11973), .ZN(
        n2109) );
  AOI221_X1 U1343 ( .B1(n12030), .B2(n8560), .C1(n12027), .C2(n8104), .A(n2082), .ZN(n2077) );
  OAI22_X1 U1344 ( .A1(n11171), .A2(n12024), .B1(n11427), .B2(n12021), .ZN(
        n2082) );
  AOI221_X1 U1345 ( .B1(n11982), .B2(n8489), .C1(n11979), .C2(n8033), .A(n2090), .ZN(n2085) );
  OAI22_X1 U1346 ( .A1(n11008), .A2(n11976), .B1(n11264), .B2(n11973), .ZN(
        n2090) );
  AOI221_X1 U1347 ( .B1(n11982), .B2(n8490), .C1(n11979), .C2(n8034), .A(n2071), .ZN(n2066) );
  OAI22_X1 U1348 ( .A1(n11009), .A2(n11976), .B1(n11265), .B2(n11973), .ZN(
        n2071) );
  AOI221_X1 U1349 ( .B1(n11982), .B2(n8491), .C1(n11979), .C2(n8035), .A(n2052), .ZN(n2047) );
  OAI22_X1 U1350 ( .A1(n11010), .A2(n11976), .B1(n11266), .B2(n11973), .ZN(
        n2052) );
  AOI221_X1 U1351 ( .B1(n11983), .B2(n8492), .C1(n11980), .C2(n8036), .A(n2033), .ZN(n2028) );
  OAI22_X1 U1352 ( .A1(n11011), .A2(n11976), .B1(n11267), .B2(n11973), .ZN(
        n2033) );
  AOI221_X1 U1353 ( .B1(n11983), .B2(n8493), .C1(n11980), .C2(n8037), .A(n2014), .ZN(n2009) );
  OAI22_X1 U1354 ( .A1(n11012), .A2(n11976), .B1(n11268), .B2(n11973), .ZN(
        n2014) );
  AOI221_X1 U1355 ( .B1(n11983), .B2(n8520), .C1(n11980), .C2(n8064), .A(n1995), .ZN(n1990) );
  OAI22_X1 U1356 ( .A1(n11061), .A2(n11977), .B1(n11317), .B2(n11974), .ZN(
        n1995) );
  AOI221_X1 U1357 ( .B1(n12031), .B2(n9559), .C1(n12028), .C2(n9871), .A(n1968), .ZN(n1963) );
  OAI22_X1 U1358 ( .A1(n11013), .A2(n12025), .B1(n11269), .B2(n12022), .ZN(
        n1968) );
  AOI221_X1 U1359 ( .B1(n11983), .B2(n9560), .C1(n11980), .C2(n9872), .A(n1976), .ZN(n1971) );
  OAI22_X1 U1360 ( .A1(n11062), .A2(n11977), .B1(n11318), .B2(n11974), .ZN(
        n1976) );
  AOI221_X1 U1361 ( .B1(n12031), .B2(n9561), .C1(n12028), .C2(n9873), .A(n1949), .ZN(n1944) );
  OAI22_X1 U1362 ( .A1(n11014), .A2(n12025), .B1(n11270), .B2(n12022), .ZN(
        n1949) );
  AOI221_X1 U1363 ( .B1(n11983), .B2(n9562), .C1(n11980), .C2(n9874), .A(n1957), .ZN(n1952) );
  OAI22_X1 U1364 ( .A1(n11063), .A2(n11977), .B1(n11319), .B2(n11974), .ZN(
        n1957) );
  AOI221_X1 U1365 ( .B1(n12031), .B2(n9563), .C1(n12028), .C2(n9875), .A(n1930), .ZN(n1925) );
  OAI22_X1 U1366 ( .A1(n11015), .A2(n12025), .B1(n11271), .B2(n12022), .ZN(
        n1930) );
  AOI221_X1 U1367 ( .B1(n11983), .B2(n9564), .C1(n11980), .C2(n9876), .A(n1938), .ZN(n1933) );
  OAI22_X1 U1368 ( .A1(n11064), .A2(n11977), .B1(n11320), .B2(n11974), .ZN(
        n1938) );
  AOI221_X1 U1369 ( .B1(n12031), .B2(n9565), .C1(n12028), .C2(n9877), .A(n1911), .ZN(n1906) );
  OAI22_X1 U1370 ( .A1(n11016), .A2(n12025), .B1(n11272), .B2(n12022), .ZN(
        n1911) );
  AOI221_X1 U1371 ( .B1(n11983), .B2(n9566), .C1(n11980), .C2(n9878), .A(n1919), .ZN(n1914) );
  OAI22_X1 U1372 ( .A1(n11065), .A2(n11977), .B1(n11321), .B2(n11974), .ZN(
        n1919) );
  AOI221_X1 U1373 ( .B1(n12031), .B2(n9567), .C1(n12028), .C2(n9879), .A(n1892), .ZN(n1887) );
  OAI22_X1 U1374 ( .A1(n11017), .A2(n12025), .B1(n11273), .B2(n12022), .ZN(
        n1892) );
  AOI221_X1 U1375 ( .B1(n11983), .B2(n9568), .C1(n11980), .C2(n9880), .A(n1900), .ZN(n1895) );
  OAI22_X1 U1376 ( .A1(n11066), .A2(n11977), .B1(n11322), .B2(n11974), .ZN(
        n1900) );
  AOI221_X1 U1377 ( .B1(n12031), .B2(n9569), .C1(n12028), .C2(n9881), .A(n1873), .ZN(n1868) );
  OAI22_X1 U1378 ( .A1(n11018), .A2(n12025), .B1(n11274), .B2(n12022), .ZN(
        n1873) );
  AOI221_X1 U1379 ( .B1(n11983), .B2(n9570), .C1(n11980), .C2(n9882), .A(n1881), .ZN(n1876) );
  OAI22_X1 U1380 ( .A1(n11067), .A2(n11977), .B1(n11323), .B2(n11974), .ZN(
        n1881) );
  AOI221_X1 U1381 ( .B1(n12031), .B2(n9571), .C1(n12028), .C2(n9883), .A(n1832), .ZN(n1817) );
  OAI22_X1 U1382 ( .A1(n11019), .A2(n12025), .B1(n11275), .B2(n12022), .ZN(
        n1832) );
  AOI221_X1 U1383 ( .B1(n11983), .B2(n9572), .C1(n11980), .C2(n9884), .A(n1856), .ZN(n1841) );
  OAI22_X1 U1384 ( .A1(n11068), .A2(n11977), .B1(n11324), .B2(n11974), .ZN(
        n1856) );
  AOI221_X1 U1385 ( .B1(n12029), .B2(n11469), .C1(n12026), .C2(n8066), .A(
        n2450), .ZN(n2439) );
  OAI22_X1 U1386 ( .A1(n11020), .A2(n12023), .B1(n11276), .B2(n12020), .ZN(
        n2450) );
  AOI221_X1 U1387 ( .B1(n11981), .B2(n11470), .C1(n11978), .C2(n8014), .A(
        n2462), .ZN(n2455) );
  OAI22_X1 U1388 ( .A1(n11021), .A2(n11975), .B1(n11277), .B2(n11972), .ZN(
        n2462) );
  AOI221_X1 U1389 ( .B1(n12029), .B2(n11471), .C1(n12026), .C2(n8068), .A(
        n2424), .ZN(n2419) );
  OAI22_X1 U1390 ( .A1(n11022), .A2(n12023), .B1(n11278), .B2(n12020), .ZN(
        n2424) );
  AOI221_X1 U1391 ( .B1(n11981), .B2(n11472), .C1(n11978), .C2(n8015), .A(
        n2432), .ZN(n2427) );
  OAI22_X1 U1392 ( .A1(n11023), .A2(n11975), .B1(n11279), .B2(n11972), .ZN(
        n2432) );
  AOI221_X1 U1393 ( .B1(n12029), .B2(n11473), .C1(n12026), .C2(n8070), .A(
        n2405), .ZN(n2400) );
  OAI22_X1 U1394 ( .A1(n11024), .A2(n12023), .B1(n11280), .B2(n12020), .ZN(
        n2405) );
  AOI221_X1 U1395 ( .B1(n11981), .B2(n11474), .C1(n11978), .C2(n8016), .A(
        n2413), .ZN(n2408) );
  OAI22_X1 U1396 ( .A1(n11025), .A2(n11975), .B1(n11281), .B2(n11972), .ZN(
        n2413) );
  AOI221_X1 U1397 ( .B1(n12029), .B2(n11475), .C1(n12026), .C2(n8072), .A(
        n2386), .ZN(n2381) );
  OAI22_X1 U1398 ( .A1(n11026), .A2(n12023), .B1(n11282), .B2(n12020), .ZN(
        n2386) );
  AOI221_X1 U1399 ( .B1(n11981), .B2(n11476), .C1(n11978), .C2(n8017), .A(
        n2394), .ZN(n2389) );
  OAI22_X1 U1400 ( .A1(n11027), .A2(n11975), .B1(n11283), .B2(n11972), .ZN(
        n2394) );
  AOI221_X1 U1401 ( .B1(n12029), .B2(n11477), .C1(n12026), .C2(n8074), .A(
        n2367), .ZN(n2362) );
  OAI22_X1 U1402 ( .A1(n11028), .A2(n12023), .B1(n11284), .B2(n12020), .ZN(
        n2367) );
  AOI221_X1 U1403 ( .B1(n11981), .B2(n11478), .C1(n11978), .C2(n8018), .A(
        n2375), .ZN(n2370) );
  OAI22_X1 U1404 ( .A1(n11029), .A2(n11975), .B1(n11285), .B2(n11972), .ZN(
        n2375) );
  AOI221_X1 U1405 ( .B1(n12029), .B2(n11479), .C1(n12026), .C2(n8076), .A(
        n2348), .ZN(n2343) );
  OAI22_X1 U1406 ( .A1(n11030), .A2(n12023), .B1(n11286), .B2(n12020), .ZN(
        n2348) );
  AOI221_X1 U1407 ( .B1(n11981), .B2(n11480), .C1(n11978), .C2(n8019), .A(
        n2356), .ZN(n2351) );
  OAI22_X1 U1408 ( .A1(n11031), .A2(n11975), .B1(n11287), .B2(n11972), .ZN(
        n2356) );
  AOI221_X1 U1409 ( .B1(n12029), .B2(n11481), .C1(n12026), .C2(n8078), .A(
        n2329), .ZN(n2324) );
  OAI22_X1 U1410 ( .A1(n11032), .A2(n12023), .B1(n11288), .B2(n12020), .ZN(
        n2329) );
  AOI221_X1 U1411 ( .B1(n11981), .B2(n11482), .C1(n11978), .C2(n8020), .A(
        n2337), .ZN(n2332) );
  OAI22_X1 U1412 ( .A1(n11033), .A2(n11975), .B1(n11289), .B2(n11972), .ZN(
        n2337) );
  AOI221_X1 U1413 ( .B1(n12029), .B2(n11483), .C1(n12026), .C2(n8080), .A(
        n2310), .ZN(n2305) );
  OAI22_X1 U1414 ( .A1(n11034), .A2(n12023), .B1(n11290), .B2(n12020), .ZN(
        n2310) );
  AOI221_X1 U1415 ( .B1(n11981), .B2(n11484), .C1(n11978), .C2(n8021), .A(
        n2318), .ZN(n2313) );
  OAI22_X1 U1416 ( .A1(n11035), .A2(n11975), .B1(n11291), .B2(n11972), .ZN(
        n2318) );
  AOI221_X1 U1417 ( .B1(n12030), .B2(n11519), .C1(n12027), .C2(n8106), .A(
        n2063), .ZN(n2058) );
  OAI22_X1 U1418 ( .A1(n11176), .A2(n12024), .B1(n11432), .B2(n12021), .ZN(
        n2063) );
  AOI221_X1 U1419 ( .B1(n12030), .B2(n11522), .C1(n12027), .C2(n8108), .A(
        n2044), .ZN(n2039) );
  OAI22_X1 U1420 ( .A1(n11180), .A2(n12024), .B1(n11436), .B2(n12021), .ZN(
        n2044) );
  AOI221_X1 U1421 ( .B1(n12031), .B2(n11524), .C1(n12028), .C2(n8110), .A(
        n2025), .ZN(n2020) );
  OAI22_X1 U1422 ( .A1(n11184), .A2(n12024), .B1(n11440), .B2(n12021), .ZN(
        n2025) );
  AOI221_X1 U1423 ( .B1(n12031), .B2(n11526), .C1(n12028), .C2(n8112), .A(
        n2006), .ZN(n2001) );
  OAI22_X1 U1424 ( .A1(n11188), .A2(n12024), .B1(n11444), .B2(n12021), .ZN(
        n2006) );
  AOI221_X1 U1425 ( .B1(n12031), .B2(n11485), .C1(n12028), .C2(n8038), .A(
        n1987), .ZN(n1982) );
  OAI22_X1 U1426 ( .A1(n11036), .A2(n12025), .B1(n11292), .B2(n12022), .ZN(
        n1987) );
  AOI221_X1 U1427 ( .B1(n12017), .B2(n8539), .C1(n12014), .C2(n8083), .A(n2292), .ZN(n2285) );
  OAI22_X1 U1428 ( .A1(n11118), .A2(n12011), .B1(n11374), .B2(n12008), .ZN(
        n2292) );
  AOI221_X1 U1429 ( .B1(n11969), .B2(n8503), .C1(n11966), .C2(n8047), .A(n2300), .ZN(n2293) );
  OAI22_X1 U1430 ( .A1(n11120), .A2(n11963), .B1(n11376), .B2(n11960), .ZN(
        n2300) );
  AOI221_X1 U1431 ( .B1(n12017), .B2(n8541), .C1(n12014), .C2(n8085), .A(n2273), .ZN(n2266) );
  OAI22_X1 U1432 ( .A1(n11124), .A2(n12011), .B1(n11380), .B2(n12008), .ZN(
        n2273) );
  AOI221_X1 U1433 ( .B1(n11969), .B2(n8504), .C1(n11966), .C2(n8048), .A(n2281), .ZN(n2274) );
  OAI22_X1 U1434 ( .A1(n11125), .A2(n11963), .B1(n11381), .B2(n11960), .ZN(
        n2281) );
  AOI221_X1 U1435 ( .B1(n12017), .B2(n8543), .C1(n12014), .C2(n8087), .A(n2254), .ZN(n2247) );
  OAI22_X1 U1436 ( .A1(n11129), .A2(n12011), .B1(n11385), .B2(n12008), .ZN(
        n2254) );
  AOI221_X1 U1437 ( .B1(n11969), .B2(n8505), .C1(n11966), .C2(n8049), .A(n2262), .ZN(n2255) );
  OAI22_X1 U1438 ( .A1(n11130), .A2(n11963), .B1(n11386), .B2(n11960), .ZN(
        n2262) );
  AOI221_X1 U1439 ( .B1(n12018), .B2(n8545), .C1(n12015), .C2(n8089), .A(n2235), .ZN(n2228) );
  OAI22_X1 U1440 ( .A1(n11134), .A2(n12011), .B1(n11390), .B2(n12008), .ZN(
        n2235) );
  AOI221_X1 U1441 ( .B1(n12018), .B2(n8547), .C1(n12015), .C2(n8091), .A(n2216), .ZN(n2209) );
  OAI22_X1 U1442 ( .A1(n11139), .A2(n12012), .B1(n11395), .B2(n12009), .ZN(
        n2216) );
  AOI221_X1 U1443 ( .B1(n12018), .B2(n8549), .C1(n12015), .C2(n8093), .A(n2197), .ZN(n2190) );
  OAI22_X1 U1444 ( .A1(n11144), .A2(n12012), .B1(n11400), .B2(n12009), .ZN(
        n2197) );
  AOI221_X1 U1445 ( .B1(n12018), .B2(n8551), .C1(n12015), .C2(n8095), .A(n2178), .ZN(n2171) );
  OAI22_X1 U1446 ( .A1(n11149), .A2(n12012), .B1(n11405), .B2(n12009), .ZN(
        n2178) );
  AOI221_X1 U1447 ( .B1(n12018), .B2(n8553), .C1(n12015), .C2(n8097), .A(n2159), .ZN(n2152) );
  OAI22_X1 U1448 ( .A1(n11154), .A2(n12012), .B1(n11410), .B2(n12009), .ZN(
        n2159) );
  AOI221_X1 U1449 ( .B1(n12018), .B2(n8555), .C1(n12015), .C2(n8099), .A(n2140), .ZN(n2133) );
  OAI22_X1 U1450 ( .A1(n11159), .A2(n12012), .B1(n11415), .B2(n12009), .ZN(
        n2140) );
  AOI221_X1 U1451 ( .B1(n12018), .B2(n8557), .C1(n12015), .C2(n8101), .A(n2121), .ZN(n2114) );
  OAI22_X1 U1452 ( .A1(n11164), .A2(n12012), .B1(n11420), .B2(n12009), .ZN(
        n2121) );
  AOI221_X1 U1453 ( .B1(n12018), .B2(n8559), .C1(n12015), .C2(n8103), .A(n2102), .ZN(n2095) );
  OAI22_X1 U1454 ( .A1(n11169), .A2(n12012), .B1(n11425), .B2(n12009), .ZN(
        n2102) );
  AOI221_X1 U1455 ( .B1(n12018), .B2(n8561), .C1(n12015), .C2(n8105), .A(n2083), .ZN(n2076) );
  OAI22_X1 U1456 ( .A1(n11174), .A2(n12012), .B1(n11430), .B2(n12009), .ZN(
        n2083) );
  AOI221_X1 U1457 ( .B1(n12018), .B2(n8565), .C1(n12015), .C2(n8109), .A(n2045), .ZN(n2038) );
  OAI22_X1 U1458 ( .A1(n11182), .A2(n12012), .B1(n11438), .B2(n12009), .ZN(
        n2045) );
  AOI221_X1 U1459 ( .B1(n12019), .B2(n8567), .C1(n12016), .C2(n8111), .A(n2026), .ZN(n2019) );
  OAI22_X1 U1460 ( .A1(n11186), .A2(n12012), .B1(n11442), .B2(n12009), .ZN(
        n2026) );
  AOI221_X1 U1461 ( .B1(n12019), .B2(n8569), .C1(n12016), .C2(n8113), .A(n2007), .ZN(n2000) );
  OAI22_X1 U1462 ( .A1(n11190), .A2(n12012), .B1(n11446), .B2(n12009), .ZN(
        n2007) );
  AOI221_X1 U1463 ( .B1(n12017), .B2(n11489), .C1(n12014), .C2(n8067), .A(
        n2453), .ZN(n2438) );
  OAI22_X1 U1464 ( .A1(n11087), .A2(n12011), .B1(n11343), .B2(n12008), .ZN(
        n2453) );
  AOI221_X1 U1465 ( .B1(n11969), .B2(n11490), .C1(n11966), .C2(n8039), .A(
        n2465), .ZN(n2454) );
  OAI22_X1 U1466 ( .A1(n11088), .A2(n11963), .B1(n11344), .B2(n11960), .ZN(
        n2465) );
  AOI221_X1 U1467 ( .B1(n12017), .B2(n11493), .C1(n12014), .C2(n8069), .A(
        n2425), .ZN(n2418) );
  OAI22_X1 U1468 ( .A1(n11091), .A2(n12011), .B1(n11347), .B2(n12008), .ZN(
        n2425) );
  AOI221_X1 U1469 ( .B1(n11969), .B2(n11494), .C1(n11966), .C2(n8040), .A(
        n2433), .ZN(n2426) );
  OAI22_X1 U1470 ( .A1(n11092), .A2(n11963), .B1(n11348), .B2(n11960), .ZN(
        n2433) );
  AOI221_X1 U1471 ( .B1(n12017), .B2(n11497), .C1(n12014), .C2(n8071), .A(
        n2406), .ZN(n2399) );
  OAI22_X1 U1472 ( .A1(n11095), .A2(n12011), .B1(n11351), .B2(n12008), .ZN(
        n2406) );
  AOI221_X1 U1473 ( .B1(n11969), .B2(n11498), .C1(n11966), .C2(n8041), .A(
        n2414), .ZN(n2407) );
  OAI22_X1 U1474 ( .A1(n11096), .A2(n11963), .B1(n11352), .B2(n11960), .ZN(
        n2414) );
  AOI221_X1 U1475 ( .B1(n12017), .B2(n11501), .C1(n12014), .C2(n8073), .A(
        n2387), .ZN(n2380) );
  OAI22_X1 U1476 ( .A1(n11099), .A2(n12011), .B1(n11355), .B2(n12008), .ZN(
        n2387) );
  AOI221_X1 U1477 ( .B1(n11969), .B2(n11502), .C1(n11966), .C2(n8042), .A(
        n2395), .ZN(n2388) );
  OAI22_X1 U1478 ( .A1(n11100), .A2(n11963), .B1(n11356), .B2(n11960), .ZN(
        n2395) );
  AOI221_X1 U1479 ( .B1(n12017), .B2(n11505), .C1(n12014), .C2(n8075), .A(
        n2368), .ZN(n2361) );
  OAI22_X1 U1480 ( .A1(n11103), .A2(n12011), .B1(n11359), .B2(n12008), .ZN(
        n2368) );
  AOI221_X1 U1481 ( .B1(n11969), .B2(n11506), .C1(n11966), .C2(n8043), .A(
        n2376), .ZN(n2369) );
  OAI22_X1 U1482 ( .A1(n11104), .A2(n11963), .B1(n11360), .B2(n11960), .ZN(
        n2376) );
  AOI221_X1 U1483 ( .B1(n12017), .B2(n11509), .C1(n12014), .C2(n8077), .A(
        n2349), .ZN(n2342) );
  OAI22_X1 U1484 ( .A1(n11107), .A2(n12011), .B1(n11363), .B2(n12008), .ZN(
        n2349) );
  AOI221_X1 U1485 ( .B1(n11969), .B2(n11510), .C1(n11966), .C2(n8044), .A(
        n2357), .ZN(n2350) );
  OAI22_X1 U1486 ( .A1(n11108), .A2(n11963), .B1(n11364), .B2(n11960), .ZN(
        n2357) );
  AOI221_X1 U1487 ( .B1(n12017), .B2(n11513), .C1(n12014), .C2(n8079), .A(
        n2330), .ZN(n2323) );
  OAI22_X1 U1488 ( .A1(n11111), .A2(n12011), .B1(n11367), .B2(n12008), .ZN(
        n2330) );
  AOI221_X1 U1489 ( .B1(n11969), .B2(n11514), .C1(n11966), .C2(n8045), .A(
        n2338), .ZN(n2331) );
  OAI22_X1 U1490 ( .A1(n11112), .A2(n11963), .B1(n11368), .B2(n11960), .ZN(
        n2338) );
  AOI221_X1 U1491 ( .B1(n12017), .B2(n11517), .C1(n12014), .C2(n8081), .A(
        n2311), .ZN(n2304) );
  OAI22_X1 U1492 ( .A1(n11115), .A2(n12011), .B1(n11371), .B2(n12008), .ZN(
        n2311) );
  AOI221_X1 U1493 ( .B1(n11969), .B2(n11518), .C1(n11966), .C2(n8046), .A(
        n2319), .ZN(n2312) );
  OAI22_X1 U1494 ( .A1(n11116), .A2(n11963), .B1(n11372), .B2(n11960), .ZN(
        n2319) );
  AOI221_X1 U1495 ( .B1(n12018), .B2(n11521), .C1(n12015), .C2(n8107), .A(
        n2064), .ZN(n2057) );
  OAI22_X1 U1496 ( .A1(n11178), .A2(n12012), .B1(n11434), .B2(n12009), .ZN(
        n2064) );
  OAI221_X1 U1497 ( .B1(n12551), .B2(n12062), .C1(n4140), .C2(n12061), .A(
        n2434), .ZN(n2539) );
  OAI21_X1 U1498 ( .B1(n2435), .B2(n2436), .A(n12056), .ZN(n2434) );
  NAND4_X1 U1499 ( .A1(n2454), .A2(n2455), .A3(n2456), .A4(n2457), .ZN(n2435)
         );
  NAND4_X1 U1500 ( .A1(n2438), .A2(n2439), .A3(n2440), .A4(n2441), .ZN(n2436)
         );
  OAI221_X1 U1501 ( .B1(n12539), .B2(n12062), .C1(n4141), .C2(n12061), .A(
        n2415), .ZN(n2540) );
  OAI21_X1 U1502 ( .B1(n2416), .B2(n2417), .A(n12056), .ZN(n2415) );
  NAND4_X1 U1503 ( .A1(n2426), .A2(n2427), .A3(n2428), .A4(n2429), .ZN(n2416)
         );
  NAND4_X1 U1504 ( .A1(n2418), .A2(n2419), .A3(n2420), .A4(n2421), .ZN(n2417)
         );
  OAI221_X1 U1505 ( .B1(n12536), .B2(n12062), .C1(n4142), .C2(n12061), .A(
        n2396), .ZN(n2541) );
  OAI21_X1 U1506 ( .B1(n2397), .B2(n2398), .A(n12056), .ZN(n2396) );
  NAND4_X1 U1507 ( .A1(n2407), .A2(n2408), .A3(n2409), .A4(n2410), .ZN(n2397)
         );
  NAND4_X1 U1508 ( .A1(n2399), .A2(n2400), .A3(n2401), .A4(n2402), .ZN(n2398)
         );
  OAI221_X1 U1509 ( .B1(n12533), .B2(n12062), .C1(n4143), .C2(n12061), .A(
        n2377), .ZN(n2542) );
  OAI21_X1 U1510 ( .B1(n2378), .B2(n2379), .A(n12056), .ZN(n2377) );
  NAND4_X1 U1511 ( .A1(n2388), .A2(n2389), .A3(n2390), .A4(n2391), .ZN(n2378)
         );
  NAND4_X1 U1512 ( .A1(n2380), .A2(n2381), .A3(n2382), .A4(n2383), .ZN(n2379)
         );
  OAI221_X1 U1513 ( .B1(n12530), .B2(n12062), .C1(n4144), .C2(n12061), .A(
        n2358), .ZN(n2543) );
  OAI21_X1 U1514 ( .B1(n2359), .B2(n2360), .A(n12056), .ZN(n2358) );
  NAND4_X1 U1515 ( .A1(n2369), .A2(n2370), .A3(n2371), .A4(n2372), .ZN(n2359)
         );
  NAND4_X1 U1516 ( .A1(n2361), .A2(n2362), .A3(n2363), .A4(n2364), .ZN(n2360)
         );
  OAI221_X1 U1517 ( .B1(n12527), .B2(n12062), .C1(n4145), .C2(n12061), .A(
        n2339), .ZN(n2544) );
  OAI21_X1 U1518 ( .B1(n2340), .B2(n2341), .A(n12056), .ZN(n2339) );
  NAND4_X1 U1519 ( .A1(n2350), .A2(n2351), .A3(n2352), .A4(n2353), .ZN(n2340)
         );
  NAND4_X1 U1520 ( .A1(n2342), .A2(n2343), .A3(n2344), .A4(n2345), .ZN(n2341)
         );
  OAI221_X1 U1521 ( .B1(n12524), .B2(n12062), .C1(n4146), .C2(n12061), .A(
        n2320), .ZN(n2545) );
  OAI21_X1 U1522 ( .B1(n2321), .B2(n2322), .A(n12056), .ZN(n2320) );
  NAND4_X1 U1523 ( .A1(n2331), .A2(n2332), .A3(n2333), .A4(n2334), .ZN(n2321)
         );
  NAND4_X1 U1524 ( .A1(n2323), .A2(n2324), .A3(n2325), .A4(n2326), .ZN(n2322)
         );
  OAI221_X1 U1525 ( .B1(n12521), .B2(n12062), .C1(n4147), .C2(n12061), .A(
        n2301), .ZN(n2546) );
  OAI21_X1 U1526 ( .B1(n2302), .B2(n2303), .A(n12056), .ZN(n2301) );
  NAND4_X1 U1527 ( .A1(n2312), .A2(n2313), .A3(n2314), .A4(n2315), .ZN(n2302)
         );
  NAND4_X1 U1528 ( .A1(n2304), .A2(n2305), .A3(n2306), .A4(n2307), .ZN(n2303)
         );
  OAI221_X1 U1529 ( .B1(n12518), .B2(n12062), .C1(n4148), .C2(n12061), .A(
        n2282), .ZN(n2547) );
  OAI21_X1 U1530 ( .B1(n2283), .B2(n2284), .A(n12056), .ZN(n2282) );
  NAND4_X1 U1531 ( .A1(n2293), .A2(n2294), .A3(n2295), .A4(n2296), .ZN(n2283)
         );
  NAND4_X1 U1532 ( .A1(n2285), .A2(n2286), .A3(n2287), .A4(n2288), .ZN(n2284)
         );
  OAI221_X1 U1533 ( .B1(n12515), .B2(n12062), .C1(n4149), .C2(n12060), .A(
        n2263), .ZN(n2548) );
  OAI21_X1 U1534 ( .B1(n2264), .B2(n2265), .A(n12056), .ZN(n2263) );
  NAND4_X1 U1535 ( .A1(n2274), .A2(n2275), .A3(n2276), .A4(n2277), .ZN(n2264)
         );
  NAND4_X1 U1536 ( .A1(n2266), .A2(n2267), .A3(n2268), .A4(n2269), .ZN(n2265)
         );
  OAI221_X1 U1537 ( .B1(n12512), .B2(n12062), .C1(n4150), .C2(n12060), .A(
        n2244), .ZN(n2549) );
  OAI21_X1 U1538 ( .B1(n2245), .B2(n2246), .A(n12056), .ZN(n2244) );
  NAND4_X1 U1539 ( .A1(n2255), .A2(n2256), .A3(n2257), .A4(n2258), .ZN(n2245)
         );
  NAND4_X1 U1540 ( .A1(n2247), .A2(n2248), .A3(n2249), .A4(n2250), .ZN(n2246)
         );
  OAI221_X1 U1541 ( .B1(n12476), .B2(n12064), .C1(n4162), .C2(n12059), .A(
        n2016), .ZN(n2561) );
  OAI21_X1 U1542 ( .B1(n2017), .B2(n2018), .A(n12058), .ZN(n2016) );
  NAND4_X1 U1543 ( .A1(n2027), .A2(n2028), .A3(n2029), .A4(n2030), .ZN(n2017)
         );
  NAND4_X1 U1544 ( .A1(n2019), .A2(n2020), .A3(n2021), .A4(n2022), .ZN(n2018)
         );
  OAI221_X1 U1545 ( .B1(n12473), .B2(n12064), .C1(n4163), .C2(n12059), .A(
        n1997), .ZN(n2562) );
  OAI21_X1 U1546 ( .B1(n1998), .B2(n1999), .A(n12058), .ZN(n1997) );
  NAND4_X1 U1547 ( .A1(n2008), .A2(n2009), .A3(n2010), .A4(n2011), .ZN(n1998)
         );
  NAND4_X1 U1548 ( .A1(n2000), .A2(n2001), .A3(n2002), .A4(n2003), .ZN(n1999)
         );
  OAI221_X1 U1549 ( .B1(n12470), .B2(n12064), .C1(n4164), .C2(n12059), .A(
        n1978), .ZN(n2563) );
  OAI21_X1 U1550 ( .B1(n1979), .B2(n1980), .A(n12058), .ZN(n1978) );
  NAND4_X1 U1551 ( .A1(n1989), .A2(n1990), .A3(n1991), .A4(n1992), .ZN(n1979)
         );
  NAND4_X1 U1552 ( .A1(n1981), .A2(n1982), .A3(n1983), .A4(n1984), .ZN(n1980)
         );
  OAI221_X1 U1553 ( .B1(n12467), .B2(n12064), .C1(n4165), .C2(n12059), .A(
        n1959), .ZN(n2564) );
  OAI21_X1 U1554 ( .B1(n1960), .B2(n1961), .A(n12058), .ZN(n1959) );
  NAND4_X1 U1555 ( .A1(n1970), .A2(n1971), .A3(n1972), .A4(n1973), .ZN(n1960)
         );
  NAND4_X1 U1556 ( .A1(n1962), .A2(n1963), .A3(n1964), .A4(n1965), .ZN(n1961)
         );
  OAI221_X1 U1557 ( .B1(n12464), .B2(n12064), .C1(n4166), .C2(n12059), .A(
        n1940), .ZN(n2565) );
  OAI21_X1 U1558 ( .B1(n1941), .B2(n1942), .A(n12058), .ZN(n1940) );
  NAND4_X1 U1559 ( .A1(n1951), .A2(n1952), .A3(n1953), .A4(n1954), .ZN(n1941)
         );
  NAND4_X1 U1560 ( .A1(n1943), .A2(n1944), .A3(n1945), .A4(n1946), .ZN(n1942)
         );
  OAI221_X1 U1561 ( .B1(n12461), .B2(n12064), .C1(n4167), .C2(n12059), .A(
        n1921), .ZN(n2566) );
  OAI21_X1 U1562 ( .B1(n1922), .B2(n1923), .A(n12058), .ZN(n1921) );
  NAND4_X1 U1563 ( .A1(n1932), .A2(n1933), .A3(n1934), .A4(n1935), .ZN(n1922)
         );
  NAND4_X1 U1564 ( .A1(n1924), .A2(n1925), .A3(n1926), .A4(n1927), .ZN(n1923)
         );
  OAI221_X1 U1565 ( .B1(n12458), .B2(n12064), .C1(n4168), .C2(n12059), .A(
        n1902), .ZN(n2567) );
  OAI21_X1 U1566 ( .B1(n1903), .B2(n1904), .A(n12058), .ZN(n1902) );
  NAND4_X1 U1567 ( .A1(n1913), .A2(n1914), .A3(n1915), .A4(n1916), .ZN(n1903)
         );
  NAND4_X1 U1568 ( .A1(n1905), .A2(n1906), .A3(n1907), .A4(n1908), .ZN(n1904)
         );
  OAI221_X1 U1569 ( .B1(n12455), .B2(n12064), .C1(n4169), .C2(n12059), .A(
        n1883), .ZN(n2568) );
  OAI21_X1 U1570 ( .B1(n1884), .B2(n1885), .A(n12058), .ZN(n1883) );
  NAND4_X1 U1571 ( .A1(n1894), .A2(n1895), .A3(n1896), .A4(n1897), .ZN(n1884)
         );
  NAND4_X1 U1572 ( .A1(n1886), .A2(n1887), .A3(n1888), .A4(n1889), .ZN(n1885)
         );
  OAI221_X1 U1573 ( .B1(n12452), .B2(n12064), .C1(n4170), .C2(n12059), .A(
        n1864), .ZN(n2569) );
  OAI21_X1 U1574 ( .B1(n1865), .B2(n1866), .A(n12058), .ZN(n1864) );
  NAND4_X1 U1575 ( .A1(n1875), .A2(n1876), .A3(n1877), .A4(n1878), .ZN(n1865)
         );
  NAND4_X1 U1576 ( .A1(n1867), .A2(n1868), .A3(n1869), .A4(n1870), .ZN(n1866)
         );
  OAI221_X1 U1577 ( .B1(n12449), .B2(n12064), .C1(n4171), .C2(n12060), .A(
        n1812), .ZN(n2570) );
  OAI21_X1 U1578 ( .B1(n1813), .B2(n1814), .A(n12058), .ZN(n1812) );
  NAND4_X1 U1579 ( .A1(n1840), .A2(n1841), .A3(n1842), .A4(n1843), .ZN(n1813)
         );
  NAND4_X1 U1580 ( .A1(n1816), .A2(n1817), .A3(n1818), .A4(n1819), .ZN(n1814)
         );
  OAI221_X1 U1581 ( .B1(n12473), .B2(n12169), .C1(n4195), .C2(n12164), .A(
        n1334), .ZN(n2594) );
  OAI21_X1 U1582 ( .B1(n1335), .B2(n1336), .A(n12163), .ZN(n1334) );
  NAND4_X1 U1583 ( .A1(n1345), .A2(n1346), .A3(n1347), .A4(n1348), .ZN(n1335)
         );
  NAND4_X1 U1584 ( .A1(n1337), .A2(n1338), .A3(n1339), .A4(n1340), .ZN(n1336)
         );
  OAI221_X1 U1585 ( .B1(n12467), .B2(n12169), .C1(n4197), .C2(n12164), .A(
        n1296), .ZN(n2596) );
  OAI21_X1 U1586 ( .B1(n1297), .B2(n1298), .A(n12163), .ZN(n1296) );
  NAND4_X1 U1587 ( .A1(n1299), .A2(n1300), .A3(n1301), .A4(n1302), .ZN(n1298)
         );
  NAND4_X1 U1588 ( .A1(n1307), .A2(n1308), .A3(n1309), .A4(n1310), .ZN(n1297)
         );
  OAI221_X1 U1589 ( .B1(n12464), .B2(n12169), .C1(n4198), .C2(n12164), .A(
        n1277), .ZN(n2597) );
  OAI21_X1 U1590 ( .B1(n1278), .B2(n1279), .A(n12163), .ZN(n1277) );
  NAND4_X1 U1591 ( .A1(n1280), .A2(n1281), .A3(n1282), .A4(n1283), .ZN(n1279)
         );
  NAND4_X1 U1592 ( .A1(n1288), .A2(n1289), .A3(n1290), .A4(n1291), .ZN(n1278)
         );
  OAI221_X1 U1593 ( .B1(n12461), .B2(n12169), .C1(n4199), .C2(n12164), .A(
        n1258), .ZN(n2598) );
  OAI21_X1 U1594 ( .B1(n1259), .B2(n1260), .A(n12163), .ZN(n1258) );
  NAND4_X1 U1595 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1260)
         );
  NAND4_X1 U1596 ( .A1(n1269), .A2(n1270), .A3(n1271), .A4(n1272), .ZN(n1259)
         );
  OAI221_X1 U1597 ( .B1(n12458), .B2(n12169), .C1(n4200), .C2(n12164), .A(
        n1239), .ZN(n2599) );
  OAI21_X1 U1598 ( .B1(n1240), .B2(n1241), .A(n12163), .ZN(n1239) );
  NAND4_X1 U1599 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1241)
         );
  NAND4_X1 U1600 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1240)
         );
  OAI221_X1 U1601 ( .B1(n12455), .B2(n12169), .C1(n4201), .C2(n12164), .A(
        n1220), .ZN(n2600) );
  OAI21_X1 U1602 ( .B1(n1221), .B2(n1222), .A(n12163), .ZN(n1220) );
  NAND4_X1 U1603 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1222)
         );
  NAND4_X1 U1604 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1221)
         );
  OAI221_X1 U1605 ( .B1(n12452), .B2(n12169), .C1(n4202), .C2(n12164), .A(
        n1201), .ZN(n2601) );
  OAI21_X1 U1606 ( .B1(n1202), .B2(n1203), .A(n12163), .ZN(n1201) );
  NAND4_X1 U1607 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203)
         );
  NAND4_X1 U1608 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1202)
         );
  OAI221_X1 U1609 ( .B1(n12449), .B2(n12169), .C1(n4203), .C2(n12165), .A(
        n1149), .ZN(n2602) );
  OAI21_X1 U1610 ( .B1(n1150), .B2(n1151), .A(n12163), .ZN(n1149) );
  NAND4_X1 U1611 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1151)
         );
  NAND4_X1 U1612 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1150)
         );
  OAI221_X1 U1613 ( .B1(n12509), .B2(n12063), .C1(n4151), .C2(n12060), .A(
        n2225), .ZN(n2550) );
  OAI21_X1 U1614 ( .B1(n2226), .B2(n2227), .A(n12057), .ZN(n2225) );
  NAND4_X1 U1615 ( .A1(n2236), .A2(n2237), .A3(n2238), .A4(n2239), .ZN(n2226)
         );
  NAND4_X1 U1616 ( .A1(n2228), .A2(n2229), .A3(n2230), .A4(n2231), .ZN(n2227)
         );
  OAI221_X1 U1617 ( .B1(n12506), .B2(n12063), .C1(n4152), .C2(n12060), .A(
        n2206), .ZN(n2551) );
  OAI21_X1 U1618 ( .B1(n2207), .B2(n2208), .A(n12057), .ZN(n2206) );
  NAND4_X1 U1619 ( .A1(n2217), .A2(n2218), .A3(n2219), .A4(n2220), .ZN(n2207)
         );
  NAND4_X1 U1620 ( .A1(n2209), .A2(n2210), .A3(n2211), .A4(n2212), .ZN(n2208)
         );
  OAI221_X1 U1621 ( .B1(n12503), .B2(n12063), .C1(n4153), .C2(n12060), .A(
        n2187), .ZN(n2552) );
  OAI21_X1 U1622 ( .B1(n2188), .B2(n2189), .A(n12057), .ZN(n2187) );
  NAND4_X1 U1623 ( .A1(n2198), .A2(n2199), .A3(n2200), .A4(n2201), .ZN(n2188)
         );
  NAND4_X1 U1624 ( .A1(n2190), .A2(n2191), .A3(n2192), .A4(n2193), .ZN(n2189)
         );
  OAI221_X1 U1625 ( .B1(n12500), .B2(n12063), .C1(n4154), .C2(n12060), .A(
        n2168), .ZN(n2553) );
  OAI21_X1 U1626 ( .B1(n2169), .B2(n2170), .A(n12057), .ZN(n2168) );
  NAND4_X1 U1627 ( .A1(n2179), .A2(n2180), .A3(n2181), .A4(n2182), .ZN(n2169)
         );
  NAND4_X1 U1628 ( .A1(n2171), .A2(n2172), .A3(n2173), .A4(n2174), .ZN(n2170)
         );
  OAI221_X1 U1629 ( .B1(n12497), .B2(n12063), .C1(n4155), .C2(n12060), .A(
        n2149), .ZN(n2554) );
  OAI21_X1 U1630 ( .B1(n2150), .B2(n2151), .A(n12057), .ZN(n2149) );
  NAND4_X1 U1631 ( .A1(n2160), .A2(n2161), .A3(n2162), .A4(n2163), .ZN(n2150)
         );
  NAND4_X1 U1632 ( .A1(n2152), .A2(n2153), .A3(n2154), .A4(n2155), .ZN(n2151)
         );
  OAI221_X1 U1633 ( .B1(n12494), .B2(n12063), .C1(n4156), .C2(n12060), .A(
        n2130), .ZN(n2555) );
  OAI21_X1 U1634 ( .B1(n2131), .B2(n2132), .A(n12057), .ZN(n2130) );
  NAND4_X1 U1635 ( .A1(n2141), .A2(n2142), .A3(n2143), .A4(n2144), .ZN(n2131)
         );
  NAND4_X1 U1636 ( .A1(n2133), .A2(n2134), .A3(n2135), .A4(n2136), .ZN(n2132)
         );
  OAI221_X1 U1637 ( .B1(n12491), .B2(n12063), .C1(n4157), .C2(n12060), .A(
        n2111), .ZN(n2556) );
  OAI21_X1 U1638 ( .B1(n2112), .B2(n2113), .A(n12057), .ZN(n2111) );
  NAND4_X1 U1639 ( .A1(n2122), .A2(n2123), .A3(n2124), .A4(n2125), .ZN(n2112)
         );
  NAND4_X1 U1640 ( .A1(n2114), .A2(n2115), .A3(n2116), .A4(n2117), .ZN(n2113)
         );
  OAI221_X1 U1641 ( .B1(n12488), .B2(n12063), .C1(n4158), .C2(n12060), .A(
        n2092), .ZN(n2557) );
  OAI21_X1 U1642 ( .B1(n2093), .B2(n2094), .A(n12057), .ZN(n2092) );
  NAND4_X1 U1643 ( .A1(n2103), .A2(n2104), .A3(n2105), .A4(n2106), .ZN(n2093)
         );
  NAND4_X1 U1644 ( .A1(n2095), .A2(n2096), .A3(n2097), .A4(n2098), .ZN(n2094)
         );
  OAI221_X1 U1645 ( .B1(n12485), .B2(n12063), .C1(n4159), .C2(n12060), .A(
        n2073), .ZN(n2558) );
  OAI21_X1 U1646 ( .B1(n2074), .B2(n2075), .A(n12057), .ZN(n2073) );
  NAND4_X1 U1647 ( .A1(n2084), .A2(n2085), .A3(n2086), .A4(n2087), .ZN(n2074)
         );
  NAND4_X1 U1648 ( .A1(n2076), .A2(n2077), .A3(n2078), .A4(n2079), .ZN(n2075)
         );
  OAI221_X1 U1649 ( .B1(n12482), .B2(n12063), .C1(n4160), .C2(n12059), .A(
        n2054), .ZN(n2559) );
  OAI21_X1 U1650 ( .B1(n2055), .B2(n2056), .A(n12057), .ZN(n2054) );
  NAND4_X1 U1651 ( .A1(n2065), .A2(n2066), .A3(n2067), .A4(n2068), .ZN(n2055)
         );
  NAND4_X1 U1652 ( .A1(n2057), .A2(n2058), .A3(n2059), .A4(n2060), .ZN(n2056)
         );
  OAI221_X1 U1653 ( .B1(n12479), .B2(n12063), .C1(n4161), .C2(n12059), .A(
        n2035), .ZN(n2560) );
  OAI21_X1 U1654 ( .B1(n2036), .B2(n2037), .A(n12057), .ZN(n2035) );
  NAND4_X1 U1655 ( .A1(n2046), .A2(n2047), .A3(n2048), .A4(n2049), .ZN(n2036)
         );
  NAND4_X1 U1656 ( .A1(n2038), .A2(n2039), .A3(n2040), .A4(n2041), .ZN(n2037)
         );
  OAI221_X1 U1657 ( .B1(n12503), .B2(n12168), .C1(n4185), .C2(n12165), .A(
        n1524), .ZN(n2584) );
  OAI21_X1 U1658 ( .B1(n1525), .B2(n1526), .A(n12162), .ZN(n1524) );
  NAND4_X1 U1659 ( .A1(n1535), .A2(n1536), .A3(n1537), .A4(n1538), .ZN(n1525)
         );
  NAND4_X1 U1660 ( .A1(n1527), .A2(n1528), .A3(n1529), .A4(n1530), .ZN(n1526)
         );
  OAI221_X1 U1661 ( .B1(n12500), .B2(n12168), .C1(n4186), .C2(n12165), .A(
        n1505), .ZN(n2585) );
  OAI21_X1 U1662 ( .B1(n1506), .B2(n1507), .A(n12162), .ZN(n1505) );
  NAND4_X1 U1663 ( .A1(n1516), .A2(n1517), .A3(n1518), .A4(n1519), .ZN(n1506)
         );
  NAND4_X1 U1664 ( .A1(n1508), .A2(n1509), .A3(n1510), .A4(n1511), .ZN(n1507)
         );
  OAI221_X1 U1665 ( .B1(n12497), .B2(n12168), .C1(n4187), .C2(n12165), .A(
        n1486), .ZN(n2586) );
  OAI21_X1 U1666 ( .B1(n1487), .B2(n1488), .A(n12162), .ZN(n1486) );
  NAND4_X1 U1667 ( .A1(n1497), .A2(n1498), .A3(n1499), .A4(n1500), .ZN(n1487)
         );
  NAND4_X1 U1668 ( .A1(n1489), .A2(n1490), .A3(n1491), .A4(n1492), .ZN(n1488)
         );
  AOI221_X1 U1669 ( .B1(n11995), .B2(n8469), .C1(n11992), .C2(n8013), .A(n1994), .ZN(n1991) );
  OAI22_X1 U1670 ( .A1(n11053), .A2(n11989), .B1(n11309), .B2(n11986), .ZN(
        n1994) );
  AOI221_X1 U1671 ( .B1(n11995), .B2(n9581), .C1(n11992), .C2(n9893), .A(n1975), .ZN(n1972) );
  OAI22_X1 U1672 ( .A1(n11054), .A2(n11989), .B1(n11310), .B2(n11986), .ZN(
        n1975) );
  AOI221_X1 U1673 ( .B1(n11995), .B2(n9584), .C1(n11992), .C2(n9896), .A(n1956), .ZN(n1953) );
  OAI22_X1 U1674 ( .A1(n11055), .A2(n11989), .B1(n11311), .B2(n11986), .ZN(
        n1956) );
  AOI221_X1 U1675 ( .B1(n11995), .B2(n9587), .C1(n11992), .C2(n9899), .A(n1937), .ZN(n1934) );
  OAI22_X1 U1676 ( .A1(n11056), .A2(n11989), .B1(n11312), .B2(n11986), .ZN(
        n1937) );
  AOI221_X1 U1677 ( .B1(n11995), .B2(n9590), .C1(n11992), .C2(n9902), .A(n1918), .ZN(n1915) );
  OAI22_X1 U1678 ( .A1(n11057), .A2(n11989), .B1(n11313), .B2(n11986), .ZN(
        n1918) );
  AOI221_X1 U1679 ( .B1(n11995), .B2(n9593), .C1(n11992), .C2(n9905), .A(n1899), .ZN(n1896) );
  OAI22_X1 U1680 ( .A1(n11058), .A2(n11989), .B1(n11314), .B2(n11986), .ZN(
        n1899) );
  AOI221_X1 U1681 ( .B1(n11995), .B2(n9596), .C1(n11992), .C2(n9908), .A(n1880), .ZN(n1877) );
  OAI22_X1 U1682 ( .A1(n11059), .A2(n11989), .B1(n11315), .B2(n11986), .ZN(
        n1880) );
  AOI221_X1 U1683 ( .B1(n11995), .B2(n9599), .C1(n11992), .C2(n9911), .A(n1851), .ZN(n1842) );
  OAI22_X1 U1684 ( .A1(n11060), .A2(n11989), .B1(n11316), .B2(n11986), .ZN(
        n1851) );
  AOI221_X1 U1685 ( .B1(n12043), .B2(n11468), .C1(n12040), .C2(n8012), .A(
        n1986), .ZN(n1983) );
  OAI22_X1 U1686 ( .A1(n10995), .A2(n12037), .B1(n11251), .B2(n12034), .ZN(
        n1986) );
  AOI221_X1 U1687 ( .B1(n12019), .B2(n8519), .C1(n12016), .C2(n8063), .A(n1988), .ZN(n1981) );
  OAI22_X1 U1688 ( .A1(n11038), .A2(n12013), .B1(n11294), .B2(n12010), .ZN(
        n1988) );
  AOI221_X1 U1689 ( .B1(n11971), .B2(n8521), .C1(n11968), .C2(n8065), .A(n1996), .ZN(n1989) );
  OAI22_X1 U1690 ( .A1(n11037), .A2(n11965), .B1(n11293), .B2(n11962), .ZN(
        n1996) );
  AOI221_X1 U1691 ( .B1(n12043), .B2(n9573), .C1(n12040), .C2(n9885), .A(n1967), .ZN(n1964) );
  OAI22_X1 U1692 ( .A1(n10976), .A2(n12037), .B1(n11232), .B2(n12034), .ZN(
        n1967) );
  AOI221_X1 U1693 ( .B1(n12019), .B2(n9580), .C1(n12016), .C2(n9892), .A(n1969), .ZN(n1962) );
  OAI22_X1 U1694 ( .A1(n11040), .A2(n12013), .B1(n11296), .B2(n12010), .ZN(
        n1969) );
  AOI221_X1 U1695 ( .B1(n11971), .B2(n9582), .C1(n11968), .C2(n9894), .A(n1977), .ZN(n1970) );
  OAI22_X1 U1696 ( .A1(n11039), .A2(n11965), .B1(n11295), .B2(n11962), .ZN(
        n1977) );
  AOI221_X1 U1697 ( .B1(n12043), .B2(n9574), .C1(n12040), .C2(n9886), .A(n1948), .ZN(n1945) );
  OAI22_X1 U1698 ( .A1(n10977), .A2(n12037), .B1(n11233), .B2(n12034), .ZN(
        n1948) );
  AOI221_X1 U1699 ( .B1(n12019), .B2(n9583), .C1(n12016), .C2(n9895), .A(n1950), .ZN(n1943) );
  OAI22_X1 U1700 ( .A1(n11042), .A2(n12013), .B1(n11298), .B2(n12010), .ZN(
        n1950) );
  AOI221_X1 U1701 ( .B1(n11971), .B2(n9585), .C1(n11968), .C2(n9897), .A(n1958), .ZN(n1951) );
  OAI22_X1 U1702 ( .A1(n11041), .A2(n11965), .B1(n11297), .B2(n11962), .ZN(
        n1958) );
  AOI221_X1 U1703 ( .B1(n12043), .B2(n9575), .C1(n12040), .C2(n9887), .A(n1929), .ZN(n1926) );
  OAI22_X1 U1704 ( .A1(n10978), .A2(n12037), .B1(n11234), .B2(n12034), .ZN(
        n1929) );
  AOI221_X1 U1705 ( .B1(n12019), .B2(n9586), .C1(n12016), .C2(n9898), .A(n1931), .ZN(n1924) );
  OAI22_X1 U1706 ( .A1(n11044), .A2(n12013), .B1(n11300), .B2(n12010), .ZN(
        n1931) );
  AOI221_X1 U1707 ( .B1(n11971), .B2(n9588), .C1(n11968), .C2(n9900), .A(n1939), .ZN(n1932) );
  OAI22_X1 U1708 ( .A1(n11043), .A2(n11965), .B1(n11299), .B2(n11962), .ZN(
        n1939) );
  AOI221_X1 U1709 ( .B1(n12043), .B2(n9576), .C1(n12040), .C2(n9888), .A(n1910), .ZN(n1907) );
  OAI22_X1 U1710 ( .A1(n10979), .A2(n12037), .B1(n11235), .B2(n12034), .ZN(
        n1910) );
  AOI221_X1 U1711 ( .B1(n12019), .B2(n9589), .C1(n12016), .C2(n9901), .A(n1912), .ZN(n1905) );
  OAI22_X1 U1712 ( .A1(n11046), .A2(n12013), .B1(n11302), .B2(n12010), .ZN(
        n1912) );
  AOI221_X1 U1713 ( .B1(n11971), .B2(n9591), .C1(n11968), .C2(n9903), .A(n1920), .ZN(n1913) );
  OAI22_X1 U1714 ( .A1(n11045), .A2(n11965), .B1(n11301), .B2(n11962), .ZN(
        n1920) );
  AOI221_X1 U1715 ( .B1(n12043), .B2(n9577), .C1(n12040), .C2(n9889), .A(n1891), .ZN(n1888) );
  OAI22_X1 U1716 ( .A1(n10980), .A2(n12037), .B1(n11236), .B2(n12034), .ZN(
        n1891) );
  AOI221_X1 U1717 ( .B1(n12019), .B2(n9592), .C1(n12016), .C2(n9904), .A(n1893), .ZN(n1886) );
  OAI22_X1 U1718 ( .A1(n11048), .A2(n12013), .B1(n11304), .B2(n12010), .ZN(
        n1893) );
  AOI221_X1 U1719 ( .B1(n11971), .B2(n9594), .C1(n11968), .C2(n9906), .A(n1901), .ZN(n1894) );
  OAI22_X1 U1720 ( .A1(n11047), .A2(n11965), .B1(n11303), .B2(n11962), .ZN(
        n1901) );
  AOI221_X1 U1721 ( .B1(n12043), .B2(n9578), .C1(n12040), .C2(n9890), .A(n1872), .ZN(n1869) );
  OAI22_X1 U1722 ( .A1(n10981), .A2(n12037), .B1(n11237), .B2(n12034), .ZN(
        n1872) );
  AOI221_X1 U1723 ( .B1(n12019), .B2(n9595), .C1(n12016), .C2(n9907), .A(n1874), .ZN(n1867) );
  OAI22_X1 U1724 ( .A1(n11050), .A2(n12013), .B1(n11306), .B2(n12010), .ZN(
        n1874) );
  AOI221_X1 U1725 ( .B1(n11971), .B2(n9597), .C1(n11968), .C2(n9909), .A(n1882), .ZN(n1875) );
  OAI22_X1 U1726 ( .A1(n11049), .A2(n11965), .B1(n11305), .B2(n11962), .ZN(
        n1882) );
  AOI221_X1 U1727 ( .B1(n12019), .B2(n9598), .C1(n12016), .C2(n9910), .A(n1837), .ZN(n1816) );
  OAI22_X1 U1728 ( .A1(n11052), .A2(n12013), .B1(n11308), .B2(n12010), .ZN(
        n1837) );
  AOI221_X1 U1729 ( .B1(n11971), .B2(n9600), .C1(n11968), .C2(n9912), .A(n1861), .ZN(n1840) );
  OAI22_X1 U1730 ( .A1(n11051), .A2(n11965), .B1(n11307), .B2(n11962), .ZN(
        n1861) );
  AOI221_X1 U1731 ( .B1(n12055), .B2(n11486), .C1(n12052), .C2(n7962), .A(
        n1985), .ZN(n1984) );
  OAI22_X1 U1732 ( .A1(n11070), .A2(n12049), .B1(n11326), .B2(n12046), .ZN(
        n1985) );
  AOI221_X1 U1733 ( .B1(n12007), .B2(n8419), .C1(n12004), .C2(n7963), .A(n1993), .ZN(n1992) );
  OAI22_X1 U1734 ( .A1(n11069), .A2(n12001), .B1(n11325), .B2(n11998), .ZN(
        n1993) );
  AOI221_X1 U1735 ( .B1(n12055), .B2(n9601), .C1(n12052), .C2(n9913), .A(n1966), .ZN(n1965) );
  OAI22_X1 U1736 ( .A1(n11072), .A2(n12049), .B1(n11328), .B2(n12046), .ZN(
        n1966) );
  AOI221_X1 U1737 ( .B1(n12007), .B2(n9552), .C1(n12004), .C2(n9864), .A(n1974), .ZN(n1973) );
  OAI22_X1 U1738 ( .A1(n11071), .A2(n12001), .B1(n11327), .B2(n11998), .ZN(
        n1974) );
  AOI221_X1 U1739 ( .B1(n12055), .B2(n9602), .C1(n12052), .C2(n9914), .A(n1947), .ZN(n1946) );
  OAI22_X1 U1740 ( .A1(n11074), .A2(n12049), .B1(n11330), .B2(n12046), .ZN(
        n1947) );
  AOI221_X1 U1741 ( .B1(n12007), .B2(n9553), .C1(n12004), .C2(n9865), .A(n1955), .ZN(n1954) );
  OAI22_X1 U1742 ( .A1(n11073), .A2(n12001), .B1(n11329), .B2(n11998), .ZN(
        n1955) );
  AOI221_X1 U1743 ( .B1(n12055), .B2(n9603), .C1(n12052), .C2(n9915), .A(n1928), .ZN(n1927) );
  OAI22_X1 U1744 ( .A1(n11076), .A2(n12049), .B1(n11332), .B2(n12046), .ZN(
        n1928) );
  AOI221_X1 U1745 ( .B1(n12007), .B2(n9554), .C1(n12004), .C2(n9866), .A(n1936), .ZN(n1935) );
  OAI22_X1 U1746 ( .A1(n11075), .A2(n12001), .B1(n11331), .B2(n11998), .ZN(
        n1936) );
  AOI221_X1 U1747 ( .B1(n12055), .B2(n9604), .C1(n12052), .C2(n9916), .A(n1909), .ZN(n1908) );
  OAI22_X1 U1748 ( .A1(n11078), .A2(n12049), .B1(n11334), .B2(n12046), .ZN(
        n1909) );
  AOI221_X1 U1749 ( .B1(n12007), .B2(n9555), .C1(n12004), .C2(n9867), .A(n1917), .ZN(n1916) );
  OAI22_X1 U1750 ( .A1(n11077), .A2(n12001), .B1(n11333), .B2(n11998), .ZN(
        n1917) );
  AOI221_X1 U1751 ( .B1(n12055), .B2(n9605), .C1(n12052), .C2(n9917), .A(n1890), .ZN(n1889) );
  OAI22_X1 U1752 ( .A1(n11080), .A2(n12049), .B1(n11336), .B2(n12046), .ZN(
        n1890) );
  AOI221_X1 U1753 ( .B1(n12007), .B2(n9556), .C1(n12004), .C2(n9868), .A(n1898), .ZN(n1897) );
  OAI22_X1 U1754 ( .A1(n11079), .A2(n12001), .B1(n11335), .B2(n11998), .ZN(
        n1898) );
  AOI221_X1 U1755 ( .B1(n12055), .B2(n9606), .C1(n12052), .C2(n9918), .A(n1871), .ZN(n1870) );
  OAI22_X1 U1756 ( .A1(n11082), .A2(n12049), .B1(n11338), .B2(n12046), .ZN(
        n1871) );
  AOI221_X1 U1757 ( .B1(n12007), .B2(n9557), .C1(n12004), .C2(n9869), .A(n1879), .ZN(n1878) );
  OAI22_X1 U1758 ( .A1(n11081), .A2(n12001), .B1(n11337), .B2(n11998), .ZN(
        n1879) );
  AOI221_X1 U1759 ( .B1(n12043), .B2(n9579), .C1(n12040), .C2(n9891), .A(n1827), .ZN(n1818) );
  OAI22_X1 U1760 ( .A1(n10982), .A2(n12037), .B1(n11238), .B2(n12034), .ZN(
        n1827) );
  AOI221_X1 U1761 ( .B1(n12055), .B2(n9607), .C1(n12052), .C2(n9919), .A(n1822), .ZN(n1819) );
  OAI22_X1 U1762 ( .A1(n11084), .A2(n12049), .B1(n11340), .B2(n12046), .ZN(
        n1822) );
  AOI221_X1 U1763 ( .B1(n12007), .B2(n9558), .C1(n12004), .C2(n9870), .A(n1846), .ZN(n1843) );
  OAI22_X1 U1764 ( .A1(n11083), .A2(n12001), .B1(n11339), .B2(n11998), .ZN(
        n1846) );
  AOI221_X1 U1765 ( .B1(n12053), .B2(n11487), .C1(n12050), .C2(n7914), .A(
        n2442), .ZN(n2441) );
  OAI22_X1 U1766 ( .A1(n11085), .A2(n12047), .B1(n11341), .B2(n12044), .ZN(
        n2442) );
  AOI221_X1 U1767 ( .B1(n12005), .B2(n11448), .C1(n12002), .C2(n7915), .A(
        n2458), .ZN(n2457) );
  OAI22_X1 U1768 ( .A1(n10951), .A2(n11999), .B1(n11207), .B2(n11996), .ZN(
        n2458) );
  AOI221_X1 U1769 ( .B1(n11993), .B2(n11456), .C1(n11990), .C2(n7965), .A(
        n2461), .ZN(n2456) );
  OAI22_X1 U1770 ( .A1(n10983), .A2(n11987), .B1(n11239), .B2(n11984), .ZN(
        n2461) );
  AOI221_X1 U1771 ( .B1(n12053), .B2(n11491), .C1(n12050), .C2(n7916), .A(
        n2422), .ZN(n2421) );
  OAI22_X1 U1772 ( .A1(n11089), .A2(n12047), .B1(n11345), .B2(n12044), .ZN(
        n2422) );
  AOI221_X1 U1773 ( .B1(n12005), .B2(n11449), .C1(n12002), .C2(n7917), .A(
        n2430), .ZN(n2429) );
  OAI22_X1 U1774 ( .A1(n10952), .A2(n11999), .B1(n11208), .B2(n11996), .ZN(
        n2430) );
  AOI221_X1 U1775 ( .B1(n11993), .B2(n11457), .C1(n11990), .C2(n7967), .A(
        n2431), .ZN(n2428) );
  OAI22_X1 U1776 ( .A1(n10984), .A2(n11987), .B1(n11240), .B2(n11984), .ZN(
        n2431) );
  AOI221_X1 U1777 ( .B1(n12053), .B2(n11495), .C1(n12050), .C2(n7918), .A(
        n2403), .ZN(n2402) );
  OAI22_X1 U1778 ( .A1(n11093), .A2(n12047), .B1(n11349), .B2(n12044), .ZN(
        n2403) );
  AOI221_X1 U1779 ( .B1(n12005), .B2(n11450), .C1(n12002), .C2(n7919), .A(
        n2411), .ZN(n2410) );
  OAI22_X1 U1780 ( .A1(n10953), .A2(n11999), .B1(n11209), .B2(n11996), .ZN(
        n2411) );
  AOI221_X1 U1781 ( .B1(n11993), .B2(n11458), .C1(n11990), .C2(n7969), .A(
        n2412), .ZN(n2409) );
  OAI22_X1 U1782 ( .A1(n10985), .A2(n11987), .B1(n11241), .B2(n11984), .ZN(
        n2412) );
  AOI221_X1 U1783 ( .B1(n12053), .B2(n11499), .C1(n12050), .C2(n7920), .A(
        n2384), .ZN(n2383) );
  OAI22_X1 U1784 ( .A1(n11097), .A2(n12047), .B1(n11353), .B2(n12044), .ZN(
        n2384) );
  AOI221_X1 U1785 ( .B1(n12005), .B2(n11451), .C1(n12002), .C2(n7921), .A(
        n2392), .ZN(n2391) );
  OAI22_X1 U1786 ( .A1(n10954), .A2(n11999), .B1(n11210), .B2(n11996), .ZN(
        n2392) );
  AOI221_X1 U1787 ( .B1(n11993), .B2(n11459), .C1(n11990), .C2(n7971), .A(
        n2393), .ZN(n2390) );
  OAI22_X1 U1788 ( .A1(n10986), .A2(n11987), .B1(n11242), .B2(n11984), .ZN(
        n2393) );
  AOI221_X1 U1789 ( .B1(n12053), .B2(n11503), .C1(n12050), .C2(n7922), .A(
        n2365), .ZN(n2364) );
  OAI22_X1 U1790 ( .A1(n11101), .A2(n12047), .B1(n11357), .B2(n12044), .ZN(
        n2365) );
  AOI221_X1 U1791 ( .B1(n12005), .B2(n11452), .C1(n12002), .C2(n7923), .A(
        n2373), .ZN(n2372) );
  OAI22_X1 U1792 ( .A1(n10955), .A2(n11999), .B1(n11211), .B2(n11996), .ZN(
        n2373) );
  AOI221_X1 U1793 ( .B1(n11993), .B2(n11460), .C1(n11990), .C2(n7973), .A(
        n2374), .ZN(n2371) );
  OAI22_X1 U1794 ( .A1(n10987), .A2(n11987), .B1(n11243), .B2(n11984), .ZN(
        n2374) );
  AOI221_X1 U1795 ( .B1(n12053), .B2(n11507), .C1(n12050), .C2(n7924), .A(
        n2346), .ZN(n2345) );
  OAI22_X1 U1796 ( .A1(n11105), .A2(n12047), .B1(n11361), .B2(n12044), .ZN(
        n2346) );
  AOI221_X1 U1797 ( .B1(n12005), .B2(n11453), .C1(n12002), .C2(n7925), .A(
        n2354), .ZN(n2353) );
  OAI22_X1 U1798 ( .A1(n10956), .A2(n11999), .B1(n11212), .B2(n11996), .ZN(
        n2354) );
  AOI221_X1 U1799 ( .B1(n11993), .B2(n11461), .C1(n11990), .C2(n7975), .A(
        n2355), .ZN(n2352) );
  OAI22_X1 U1800 ( .A1(n10988), .A2(n11987), .B1(n11244), .B2(n11984), .ZN(
        n2355) );
  AOI221_X1 U1801 ( .B1(n12053), .B2(n11511), .C1(n12050), .C2(n7926), .A(
        n2327), .ZN(n2326) );
  OAI22_X1 U1802 ( .A1(n11109), .A2(n12047), .B1(n11365), .B2(n12044), .ZN(
        n2327) );
  AOI221_X1 U1803 ( .B1(n12005), .B2(n11454), .C1(n12002), .C2(n7927), .A(
        n2335), .ZN(n2334) );
  OAI22_X1 U1804 ( .A1(n10957), .A2(n11999), .B1(n11213), .B2(n11996), .ZN(
        n2335) );
  AOI221_X1 U1805 ( .B1(n11993), .B2(n11462), .C1(n11990), .C2(n7977), .A(
        n2336), .ZN(n2333) );
  OAI22_X1 U1806 ( .A1(n10989), .A2(n11987), .B1(n11245), .B2(n11984), .ZN(
        n2336) );
  AOI221_X1 U1807 ( .B1(n12053), .B2(n11515), .C1(n12050), .C2(n7928), .A(
        n2308), .ZN(n2307) );
  OAI22_X1 U1808 ( .A1(n11113), .A2(n12047), .B1(n11369), .B2(n12044), .ZN(
        n2308) );
  AOI221_X1 U1809 ( .B1(n12005), .B2(n11455), .C1(n12002), .C2(n7929), .A(
        n2316), .ZN(n2315) );
  OAI22_X1 U1810 ( .A1(n10958), .A2(n11999), .B1(n11214), .B2(n11996), .ZN(
        n2316) );
  AOI221_X1 U1811 ( .B1(n11993), .B2(n11463), .C1(n11990), .C2(n7979), .A(
        n2317), .ZN(n2314) );
  OAI22_X1 U1812 ( .A1(n10990), .A2(n11987), .B1(n11246), .B2(n11984), .ZN(
        n2317) );
  AOI221_X1 U1813 ( .B1(n12053), .B2(n8386), .C1(n12050), .C2(n7930), .A(n2289), .ZN(n2288) );
  OAI22_X1 U1814 ( .A1(n11117), .A2(n12047), .B1(n11373), .B2(n12044), .ZN(
        n2289) );
  AOI221_X1 U1815 ( .B1(n12005), .B2(n8387), .C1(n12002), .C2(n7931), .A(n2297), .ZN(n2296) );
  OAI22_X1 U1816 ( .A1(n11119), .A2(n11999), .B1(n11375), .B2(n11996), .ZN(
        n2297) );
  AOI221_X1 U1817 ( .B1(n11993), .B2(n8437), .C1(n11990), .C2(n7981), .A(n2298), .ZN(n2295) );
  OAI22_X1 U1818 ( .A1(n10960), .A2(n11987), .B1(n11216), .B2(n11984), .ZN(
        n2298) );
  AOI221_X1 U1819 ( .B1(n12053), .B2(n8388), .C1(n12050), .C2(n7932), .A(n2270), .ZN(n2269) );
  OAI22_X1 U1820 ( .A1(n11122), .A2(n12047), .B1(n11378), .B2(n12044), .ZN(
        n2270) );
  AOI221_X1 U1821 ( .B1(n12005), .B2(n8389), .C1(n12002), .C2(n7933), .A(n2278), .ZN(n2277) );
  OAI22_X1 U1822 ( .A1(n10936), .A2(n11999), .B1(n11192), .B2(n11996), .ZN(
        n2278) );
  AOI221_X1 U1823 ( .B1(n11993), .B2(n8439), .C1(n11990), .C2(n7983), .A(n2279), .ZN(n2276) );
  OAI22_X1 U1824 ( .A1(n10961), .A2(n11987), .B1(n11217), .B2(n11984), .ZN(
        n2279) );
  AOI221_X1 U1825 ( .B1(n12053), .B2(n8390), .C1(n12050), .C2(n7934), .A(n2251), .ZN(n2250) );
  OAI22_X1 U1826 ( .A1(n11127), .A2(n12047), .B1(n11383), .B2(n12044), .ZN(
        n2251) );
  AOI221_X1 U1827 ( .B1(n12005), .B2(n8391), .C1(n12002), .C2(n7935), .A(n2259), .ZN(n2258) );
  OAI22_X1 U1828 ( .A1(n10937), .A2(n11999), .B1(n11193), .B2(n11996), .ZN(
        n2259) );
  AOI221_X1 U1829 ( .B1(n11993), .B2(n8441), .C1(n11990), .C2(n7985), .A(n2260), .ZN(n2257) );
  OAI22_X1 U1830 ( .A1(n10962), .A2(n11987), .B1(n11218), .B2(n11984), .ZN(
        n2260) );
  AOI221_X1 U1831 ( .B1(n12054), .B2(n8392), .C1(n12051), .C2(n7936), .A(n2232), .ZN(n2231) );
  OAI22_X1 U1832 ( .A1(n11132), .A2(n12047), .B1(n11388), .B2(n12044), .ZN(
        n2232) );
  AOI221_X1 U1833 ( .B1(n12006), .B2(n8393), .C1(n12003), .C2(n7937), .A(n2240), .ZN(n2239) );
  OAI22_X1 U1834 ( .A1(n10938), .A2(n11999), .B1(n11194), .B2(n11996), .ZN(
        n2240) );
  AOI221_X1 U1835 ( .B1(n11994), .B2(n8443), .C1(n11991), .C2(n7987), .A(n2241), .ZN(n2238) );
  OAI22_X1 U1836 ( .A1(n10963), .A2(n11987), .B1(n11219), .B2(n11984), .ZN(
        n2241) );
  AOI221_X1 U1837 ( .B1(n11970), .B2(n8506), .C1(n11967), .C2(n8050), .A(n2243), .ZN(n2236) );
  OAI22_X1 U1838 ( .A1(n11135), .A2(n11963), .B1(n11391), .B2(n11960), .ZN(
        n2243) );
  AOI221_X1 U1839 ( .B1(n12054), .B2(n8394), .C1(n12051), .C2(n7938), .A(n2213), .ZN(n2212) );
  OAI22_X1 U1840 ( .A1(n11137), .A2(n12048), .B1(n11393), .B2(n12045), .ZN(
        n2213) );
  AOI221_X1 U1841 ( .B1(n12006), .B2(n8395), .C1(n12003), .C2(n7939), .A(n2221), .ZN(n2220) );
  OAI22_X1 U1842 ( .A1(n10939), .A2(n12000), .B1(n11195), .B2(n11997), .ZN(
        n2221) );
  AOI221_X1 U1843 ( .B1(n11994), .B2(n8445), .C1(n11991), .C2(n7989), .A(n2222), .ZN(n2219) );
  OAI22_X1 U1844 ( .A1(n10964), .A2(n11988), .B1(n11220), .B2(n11985), .ZN(
        n2222) );
  AOI221_X1 U1845 ( .B1(n11970), .B2(n8507), .C1(n11967), .C2(n8051), .A(n2224), .ZN(n2217) );
  OAI22_X1 U1846 ( .A1(n11140), .A2(n11964), .B1(n11396), .B2(n11961), .ZN(
        n2224) );
  AOI221_X1 U1847 ( .B1(n12054), .B2(n8396), .C1(n12051), .C2(n7940), .A(n2194), .ZN(n2193) );
  OAI22_X1 U1848 ( .A1(n11142), .A2(n12048), .B1(n11398), .B2(n12045), .ZN(
        n2194) );
  AOI221_X1 U1849 ( .B1(n12006), .B2(n8397), .C1(n12003), .C2(n7941), .A(n2202), .ZN(n2201) );
  OAI22_X1 U1850 ( .A1(n10940), .A2(n12000), .B1(n11196), .B2(n11997), .ZN(
        n2202) );
  AOI221_X1 U1851 ( .B1(n11994), .B2(n8447), .C1(n11991), .C2(n7991), .A(n2203), .ZN(n2200) );
  OAI22_X1 U1852 ( .A1(n10965), .A2(n11988), .B1(n11221), .B2(n11985), .ZN(
        n2203) );
  AOI221_X1 U1853 ( .B1(n11970), .B2(n8508), .C1(n11967), .C2(n8052), .A(n2205), .ZN(n2198) );
  OAI22_X1 U1854 ( .A1(n11145), .A2(n11964), .B1(n11401), .B2(n11961), .ZN(
        n2205) );
  AOI221_X1 U1855 ( .B1(n12054), .B2(n8398), .C1(n12051), .C2(n7942), .A(n2175), .ZN(n2174) );
  OAI22_X1 U1856 ( .A1(n11147), .A2(n12048), .B1(n11403), .B2(n12045), .ZN(
        n2175) );
  AOI221_X1 U1857 ( .B1(n12006), .B2(n8399), .C1(n12003), .C2(n7943), .A(n2183), .ZN(n2182) );
  OAI22_X1 U1858 ( .A1(n10941), .A2(n12000), .B1(n11197), .B2(n11997), .ZN(
        n2183) );
  AOI221_X1 U1859 ( .B1(n11994), .B2(n8449), .C1(n11991), .C2(n7993), .A(n2184), .ZN(n2181) );
  OAI22_X1 U1860 ( .A1(n10966), .A2(n11988), .B1(n11222), .B2(n11985), .ZN(
        n2184) );
  AOI221_X1 U1861 ( .B1(n11970), .B2(n8509), .C1(n11967), .C2(n8053), .A(n2186), .ZN(n2179) );
  OAI22_X1 U1862 ( .A1(n11150), .A2(n11964), .B1(n11406), .B2(n11961), .ZN(
        n2186) );
  AOI221_X1 U1863 ( .B1(n12054), .B2(n8400), .C1(n12051), .C2(n7944), .A(n2156), .ZN(n2155) );
  OAI22_X1 U1864 ( .A1(n11152), .A2(n12048), .B1(n11408), .B2(n12045), .ZN(
        n2156) );
  AOI221_X1 U1865 ( .B1(n12006), .B2(n8401), .C1(n12003), .C2(n7945), .A(n2164), .ZN(n2163) );
  OAI22_X1 U1866 ( .A1(n10942), .A2(n12000), .B1(n11198), .B2(n11997), .ZN(
        n2164) );
  AOI221_X1 U1867 ( .B1(n11994), .B2(n8451), .C1(n11991), .C2(n7995), .A(n2165), .ZN(n2162) );
  OAI22_X1 U1868 ( .A1(n10967), .A2(n11988), .B1(n11223), .B2(n11985), .ZN(
        n2165) );
  AOI221_X1 U1869 ( .B1(n11970), .B2(n8510), .C1(n11967), .C2(n8054), .A(n2167), .ZN(n2160) );
  OAI22_X1 U1870 ( .A1(n11155), .A2(n11964), .B1(n11411), .B2(n11961), .ZN(
        n2167) );
  AOI221_X1 U1871 ( .B1(n12054), .B2(n8402), .C1(n12051), .C2(n7946), .A(n2137), .ZN(n2136) );
  OAI22_X1 U1872 ( .A1(n11157), .A2(n12048), .B1(n11413), .B2(n12045), .ZN(
        n2137) );
  AOI221_X1 U1873 ( .B1(n12006), .B2(n8403), .C1(n12003), .C2(n7947), .A(n2145), .ZN(n2144) );
  OAI22_X1 U1874 ( .A1(n10943), .A2(n12000), .B1(n11199), .B2(n11997), .ZN(
        n2145) );
  AOI221_X1 U1875 ( .B1(n11994), .B2(n8453), .C1(n11991), .C2(n7997), .A(n2146), .ZN(n2143) );
  OAI22_X1 U1876 ( .A1(n10968), .A2(n11988), .B1(n11224), .B2(n11985), .ZN(
        n2146) );
  AOI221_X1 U1877 ( .B1(n11970), .B2(n8511), .C1(n11967), .C2(n8055), .A(n2148), .ZN(n2141) );
  OAI22_X1 U1878 ( .A1(n11160), .A2(n11964), .B1(n11416), .B2(n11961), .ZN(
        n2148) );
  AOI221_X1 U1879 ( .B1(n12054), .B2(n8404), .C1(n12051), .C2(n7948), .A(n2118), .ZN(n2117) );
  OAI22_X1 U1880 ( .A1(n11162), .A2(n12048), .B1(n11418), .B2(n12045), .ZN(
        n2118) );
  AOI221_X1 U1881 ( .B1(n12006), .B2(n8405), .C1(n12003), .C2(n7949), .A(n2126), .ZN(n2125) );
  OAI22_X1 U1882 ( .A1(n10944), .A2(n12000), .B1(n11200), .B2(n11997), .ZN(
        n2126) );
  AOI221_X1 U1883 ( .B1(n11994), .B2(n8455), .C1(n11991), .C2(n7999), .A(n2127), .ZN(n2124) );
  OAI22_X1 U1884 ( .A1(n10969), .A2(n11988), .B1(n11225), .B2(n11985), .ZN(
        n2127) );
  AOI221_X1 U1885 ( .B1(n11970), .B2(n8512), .C1(n11967), .C2(n8056), .A(n2129), .ZN(n2122) );
  OAI22_X1 U1886 ( .A1(n11165), .A2(n11964), .B1(n11421), .B2(n11961), .ZN(
        n2129) );
  AOI221_X1 U1887 ( .B1(n12054), .B2(n8406), .C1(n12051), .C2(n7950), .A(n2099), .ZN(n2098) );
  OAI22_X1 U1888 ( .A1(n11167), .A2(n12048), .B1(n11423), .B2(n12045), .ZN(
        n2099) );
  AOI221_X1 U1889 ( .B1(n12006), .B2(n8407), .C1(n12003), .C2(n7951), .A(n2107), .ZN(n2106) );
  OAI22_X1 U1890 ( .A1(n10945), .A2(n12000), .B1(n11201), .B2(n11997), .ZN(
        n2107) );
  AOI221_X1 U1891 ( .B1(n11994), .B2(n8457), .C1(n11991), .C2(n8001), .A(n2108), .ZN(n2105) );
  OAI22_X1 U1892 ( .A1(n10970), .A2(n11988), .B1(n11226), .B2(n11985), .ZN(
        n2108) );
  AOI221_X1 U1893 ( .B1(n11970), .B2(n8513), .C1(n11967), .C2(n8057), .A(n2110), .ZN(n2103) );
  OAI22_X1 U1894 ( .A1(n11170), .A2(n11964), .B1(n11426), .B2(n11961), .ZN(
        n2110) );
  AOI221_X1 U1895 ( .B1(n12054), .B2(n8408), .C1(n12051), .C2(n7952), .A(n2080), .ZN(n2079) );
  OAI22_X1 U1896 ( .A1(n11172), .A2(n12048), .B1(n11428), .B2(n12045), .ZN(
        n2080) );
  AOI221_X1 U1897 ( .B1(n12006), .B2(n8409), .C1(n12003), .C2(n7953), .A(n2088), .ZN(n2087) );
  OAI22_X1 U1898 ( .A1(n10946), .A2(n12000), .B1(n11202), .B2(n11997), .ZN(
        n2088) );
  AOI221_X1 U1899 ( .B1(n11994), .B2(n8459), .C1(n11991), .C2(n8003), .A(n2089), .ZN(n2086) );
  OAI22_X1 U1900 ( .A1(n10971), .A2(n11988), .B1(n11227), .B2(n11985), .ZN(
        n2089) );
  AOI221_X1 U1901 ( .B1(n11970), .B2(n8514), .C1(n11967), .C2(n8058), .A(n2091), .ZN(n2084) );
  OAI22_X1 U1902 ( .A1(n11175), .A2(n11964), .B1(n11431), .B2(n11961), .ZN(
        n2091) );
  AOI221_X1 U1903 ( .B1(n12054), .B2(n11520), .C1(n12051), .C2(n7954), .A(
        n2061), .ZN(n2060) );
  OAI22_X1 U1904 ( .A1(n11177), .A2(n12048), .B1(n11433), .B2(n12045), .ZN(
        n2061) );
  AOI221_X1 U1905 ( .B1(n12006), .B2(n8411), .C1(n12003), .C2(n7955), .A(n2069), .ZN(n2068) );
  OAI22_X1 U1906 ( .A1(n10947), .A2(n12000), .B1(n11203), .B2(n11997), .ZN(
        n2069) );
  AOI221_X1 U1907 ( .B1(n11994), .B2(n8461), .C1(n11991), .C2(n8005), .A(n2070), .ZN(n2067) );
  OAI22_X1 U1908 ( .A1(n10972), .A2(n11988), .B1(n11228), .B2(n11985), .ZN(
        n2070) );
  AOI221_X1 U1909 ( .B1(n11970), .B2(n8515), .C1(n11967), .C2(n8059), .A(n2072), .ZN(n2065) );
  OAI22_X1 U1910 ( .A1(n11179), .A2(n11964), .B1(n11435), .B2(n11961), .ZN(
        n2072) );
  AOI221_X1 U1911 ( .B1(n12054), .B2(n11523), .C1(n12051), .C2(n7956), .A(
        n2042), .ZN(n2041) );
  OAI22_X1 U1912 ( .A1(n11181), .A2(n12048), .B1(n11437), .B2(n12045), .ZN(
        n2042) );
  AOI221_X1 U1913 ( .B1(n12006), .B2(n8413), .C1(n12003), .C2(n7957), .A(n2050), .ZN(n2049) );
  OAI22_X1 U1914 ( .A1(n10948), .A2(n12000), .B1(n11204), .B2(n11997), .ZN(
        n2050) );
  AOI221_X1 U1915 ( .B1(n11994), .B2(n8463), .C1(n11991), .C2(n8007), .A(n2051), .ZN(n2048) );
  OAI22_X1 U1916 ( .A1(n10973), .A2(n11988), .B1(n11229), .B2(n11985), .ZN(
        n2051) );
  AOI221_X1 U1917 ( .B1(n11970), .B2(n8516), .C1(n11967), .C2(n8060), .A(n2053), .ZN(n2046) );
  OAI22_X1 U1918 ( .A1(n11183), .A2(n11964), .B1(n11439), .B2(n11961), .ZN(
        n2053) );
  AOI221_X1 U1919 ( .B1(n12055), .B2(n11525), .C1(n12052), .C2(n7958), .A(
        n2023), .ZN(n2022) );
  OAI22_X1 U1920 ( .A1(n11185), .A2(n12048), .B1(n11441), .B2(n12045), .ZN(
        n2023) );
  AOI221_X1 U1921 ( .B1(n12007), .B2(n8415), .C1(n12004), .C2(n7959), .A(n2031), .ZN(n2030) );
  OAI22_X1 U1922 ( .A1(n10949), .A2(n12000), .B1(n11205), .B2(n11997), .ZN(
        n2031) );
  AOI221_X1 U1923 ( .B1(n11995), .B2(n8465), .C1(n11992), .C2(n8009), .A(n2032), .ZN(n2029) );
  OAI22_X1 U1924 ( .A1(n10974), .A2(n11988), .B1(n11230), .B2(n11985), .ZN(
        n2032) );
  AOI221_X1 U1925 ( .B1(n11971), .B2(n8517), .C1(n11968), .C2(n8061), .A(n2034), .ZN(n2027) );
  OAI22_X1 U1926 ( .A1(n11187), .A2(n11964), .B1(n11443), .B2(n11961), .ZN(
        n2034) );
  AOI221_X1 U1927 ( .B1(n12055), .B2(n11527), .C1(n12052), .C2(n7960), .A(
        n2004), .ZN(n2003) );
  OAI22_X1 U1928 ( .A1(n11189), .A2(n12048), .B1(n11445), .B2(n12045), .ZN(
        n2004) );
  AOI221_X1 U1929 ( .B1(n12007), .B2(n8417), .C1(n12004), .C2(n7961), .A(n2012), .ZN(n2011) );
  OAI22_X1 U1930 ( .A1(n10950), .A2(n12000), .B1(n11206), .B2(n11997), .ZN(
        n2012) );
  AOI221_X1 U1931 ( .B1(n11995), .B2(n8467), .C1(n11992), .C2(n8011), .A(n2013), .ZN(n2010) );
  OAI22_X1 U1932 ( .A1(n10975), .A2(n11988), .B1(n11231), .B2(n11985), .ZN(
        n2013) );
  AOI221_X1 U1933 ( .B1(n11971), .B2(n8518), .C1(n11968), .C2(n8062), .A(n2015), .ZN(n2008) );
  OAI22_X1 U1934 ( .A1(n11191), .A2(n11964), .B1(n11447), .B2(n11961), .ZN(
        n2015) );
  OAI22_X1 U1935 ( .A1(n12175), .A2(n12515), .B1(n12170), .B2(n11784), .ZN(
        n2612) );
  OAI22_X1 U1936 ( .A1(n12175), .A2(n12512), .B1(n12170), .B2(n11785), .ZN(
        n2613) );
  OAI22_X1 U1937 ( .A1(n12175), .A2(n12509), .B1(n12170), .B2(n11786), .ZN(
        n2614) );
  OAI22_X1 U1938 ( .A1(n12174), .A2(n12506), .B1(n12170), .B2(n11787), .ZN(
        n2615) );
  OAI22_X1 U1939 ( .A1(n12174), .A2(n12503), .B1(n12170), .B2(n11788), .ZN(
        n2616) );
  OAI22_X1 U1940 ( .A1(n12174), .A2(n12500), .B1(n12170), .B2(n11789), .ZN(
        n2617) );
  OAI22_X1 U1941 ( .A1(n12174), .A2(n12497), .B1(n12170), .B2(n11790), .ZN(
        n2618) );
  OAI22_X1 U1942 ( .A1(n12174), .A2(n12494), .B1(n12170), .B2(n11791), .ZN(
        n2619) );
  OAI22_X1 U1943 ( .A1(n12193), .A2(n12515), .B1(n12188), .B2(n11792), .ZN(
        n2740) );
  OAI22_X1 U1944 ( .A1(n12193), .A2(n12512), .B1(n12188), .B2(n11793), .ZN(
        n2741) );
  OAI22_X1 U1945 ( .A1(n12193), .A2(n12509), .B1(n12188), .B2(n11794), .ZN(
        n2742) );
  OAI22_X1 U1946 ( .A1(n12192), .A2(n12506), .B1(n12188), .B2(n11795), .ZN(
        n2743) );
  OAI22_X1 U1947 ( .A1(n12192), .A2(n12503), .B1(n12188), .B2(n11796), .ZN(
        n2744) );
  OAI22_X1 U1948 ( .A1(n12192), .A2(n12500), .B1(n12188), .B2(n11797), .ZN(
        n2745) );
  OAI22_X1 U1949 ( .A1(n12192), .A2(n12497), .B1(n12188), .B2(n11798), .ZN(
        n2746) );
  OAI22_X1 U1950 ( .A1(n12192), .A2(n12494), .B1(n12188), .B2(n11799), .ZN(
        n2747) );
  OAI22_X1 U1951 ( .A1(n12211), .A2(n12515), .B1(n1142), .B2(n11800), .ZN(
        n2868) );
  OAI22_X1 U1952 ( .A1(n12211), .A2(n12512), .B1(n1142), .B2(n11801), .ZN(
        n2869) );
  OAI22_X1 U1953 ( .A1(n12211), .A2(n12509), .B1(n1142), .B2(n11802), .ZN(
        n2870) );
  OAI22_X1 U1954 ( .A1(n12210), .A2(n12506), .B1(n12206), .B2(n11803), .ZN(
        n2871) );
  OAI22_X1 U1955 ( .A1(n12210), .A2(n12503), .B1(n12206), .B2(n11804), .ZN(
        n2872) );
  OAI22_X1 U1956 ( .A1(n12210), .A2(n12500), .B1(n12206), .B2(n11805), .ZN(
        n2873) );
  OAI22_X1 U1957 ( .A1(n12210), .A2(n12497), .B1(n12206), .B2(n11806), .ZN(
        n2874) );
  OAI22_X1 U1958 ( .A1(n12210), .A2(n12494), .B1(n12206), .B2(n11807), .ZN(
        n2875) );
  OAI22_X1 U1959 ( .A1(n12247), .A2(n12515), .B1(n12242), .B2(n11808), .ZN(
        n2996) );
  OAI22_X1 U1960 ( .A1(n12247), .A2(n12512), .B1(n12242), .B2(n11809), .ZN(
        n2997) );
  OAI22_X1 U1961 ( .A1(n12247), .A2(n12509), .B1(n12242), .B2(n11810), .ZN(
        n2998) );
  OAI22_X1 U1962 ( .A1(n12246), .A2(n12506), .B1(n12242), .B2(n11811), .ZN(
        n2999) );
  OAI22_X1 U1963 ( .A1(n12246), .A2(n12503), .B1(n12242), .B2(n11812), .ZN(
        n3000) );
  OAI22_X1 U1964 ( .A1(n12246), .A2(n12500), .B1(n1138), .B2(n11813), .ZN(
        n3001) );
  OAI22_X1 U1965 ( .A1(n12246), .A2(n12497), .B1(n1138), .B2(n11814), .ZN(
        n3002) );
  OAI22_X1 U1966 ( .A1(n12246), .A2(n12494), .B1(n1138), .B2(n11815), .ZN(
        n3003) );
  OAI22_X1 U1967 ( .A1(n12280), .A2(n12471), .B1(n12278), .B2(n11816), .ZN(
        n3139) );
  OAI22_X1 U1968 ( .A1(n12280), .A2(n12468), .B1(n1133), .B2(n11817), .ZN(
        n3140) );
  OAI22_X1 U1969 ( .A1(n12280), .A2(n12465), .B1(n12278), .B2(n11818), .ZN(
        n3141) );
  OAI22_X1 U1970 ( .A1(n12279), .A2(n12462), .B1(n12278), .B2(n11819), .ZN(
        n3142) );
  OAI22_X1 U1971 ( .A1(n12279), .A2(n12459), .B1(n12278), .B2(n11820), .ZN(
        n3143) );
  OAI22_X1 U1972 ( .A1(n12279), .A2(n12456), .B1(n1133), .B2(n11821), .ZN(
        n3144) );
  OAI22_X1 U1973 ( .A1(n12279), .A2(n12453), .B1(n1133), .B2(n11822), .ZN(
        n3145) );
  OAI22_X1 U1974 ( .A1(n12279), .A2(n12450), .B1(n1133), .B2(n11823), .ZN(
        n3146) );
  OAI22_X1 U1975 ( .A1(n12316), .A2(n12471), .B1(n12314), .B2(n11824), .ZN(
        n3267) );
  OAI22_X1 U1976 ( .A1(n12316), .A2(n12468), .B1(n1129), .B2(n11825), .ZN(
        n3268) );
  OAI22_X1 U1977 ( .A1(n12316), .A2(n12465), .B1(n12314), .B2(n11826), .ZN(
        n3269) );
  OAI22_X1 U1978 ( .A1(n12315), .A2(n12462), .B1(n12314), .B2(n11827), .ZN(
        n3270) );
  OAI22_X1 U1979 ( .A1(n12315), .A2(n12459), .B1(n12314), .B2(n11828), .ZN(
        n3271) );
  OAI22_X1 U1980 ( .A1(n12315), .A2(n12456), .B1(n1129), .B2(n11829), .ZN(
        n3272) );
  OAI22_X1 U1981 ( .A1(n12315), .A2(n12453), .B1(n1129), .B2(n11830), .ZN(
        n3273) );
  OAI22_X1 U1982 ( .A1(n12315), .A2(n12450), .B1(n1129), .B2(n11831), .ZN(
        n3274) );
  OAI22_X1 U1983 ( .A1(n12361), .A2(n12471), .B1(n12359), .B2(n11832), .ZN(
        n3491) );
  OAI22_X1 U1984 ( .A1(n12361), .A2(n12468), .B1(n1123), .B2(n11833), .ZN(
        n3492) );
  OAI22_X1 U1985 ( .A1(n12361), .A2(n12465), .B1(n12359), .B2(n11834), .ZN(
        n3493) );
  OAI22_X1 U1986 ( .A1(n12360), .A2(n12462), .B1(n12359), .B2(n11835), .ZN(
        n3494) );
  OAI22_X1 U1987 ( .A1(n12360), .A2(n12459), .B1(n12359), .B2(n11836), .ZN(
        n3495) );
  OAI22_X1 U1988 ( .A1(n12360), .A2(n12456), .B1(n1123), .B2(n11837), .ZN(
        n3496) );
  OAI22_X1 U1989 ( .A1(n12360), .A2(n12453), .B1(n1123), .B2(n11838), .ZN(
        n3497) );
  OAI22_X1 U1990 ( .A1(n12360), .A2(n12450), .B1(n1123), .B2(n11839), .ZN(
        n3498) );
  OAI22_X1 U1991 ( .A1(n12379), .A2(n12472), .B1(n12377), .B2(n11840), .ZN(
        n3619) );
  OAI22_X1 U1992 ( .A1(n12379), .A2(n12469), .B1(n1121), .B2(n11841), .ZN(
        n3620) );
  OAI22_X1 U1993 ( .A1(n12379), .A2(n12466), .B1(n12377), .B2(n11842), .ZN(
        n3621) );
  OAI22_X1 U1994 ( .A1(n12378), .A2(n12463), .B1(n12377), .B2(n11843), .ZN(
        n3622) );
  OAI22_X1 U1995 ( .A1(n12378), .A2(n12460), .B1(n12377), .B2(n11844), .ZN(
        n3623) );
  OAI22_X1 U1996 ( .A1(n12378), .A2(n12457), .B1(n1121), .B2(n11845), .ZN(
        n3624) );
  OAI22_X1 U1997 ( .A1(n12378), .A2(n12454), .B1(n1121), .B2(n11846), .ZN(
        n3625) );
  OAI22_X1 U1998 ( .A1(n12378), .A2(n12451), .B1(n1121), .B2(n11847), .ZN(
        n3626) );
  OAI22_X1 U1999 ( .A1(n12247), .A2(n12518), .B1(n12242), .B2(n11848), .ZN(
        n2995) );
  OAI22_X1 U2000 ( .A1(n12243), .A2(n12455), .B1(n12242), .B2(n11849), .ZN(
        n3016) );
  OAI22_X1 U2001 ( .A1(n12243), .A2(n12452), .B1(n12242), .B2(n11850), .ZN(
        n3017) );
  OAI22_X1 U2002 ( .A1(n12283), .A2(n12519), .B1(n12278), .B2(n11851), .ZN(
        n3123) );
  OAI22_X1 U2003 ( .A1(n12283), .A2(n12516), .B1(n12278), .B2(n11852), .ZN(
        n3124) );
  OAI22_X1 U2004 ( .A1(n12283), .A2(n12513), .B1(n12278), .B2(n11853), .ZN(
        n3125) );
  OAI22_X1 U2005 ( .A1(n12283), .A2(n12510), .B1(n12278), .B2(n11854), .ZN(
        n3126) );
  OAI22_X1 U2006 ( .A1(n12319), .A2(n12519), .B1(n12314), .B2(n11855), .ZN(
        n3251) );
  OAI22_X1 U2007 ( .A1(n12319), .A2(n12516), .B1(n12314), .B2(n11856), .ZN(
        n3252) );
  OAI22_X1 U2008 ( .A1(n12319), .A2(n12513), .B1(n12314), .B2(n11857), .ZN(
        n3253) );
  OAI22_X1 U2009 ( .A1(n12319), .A2(n12510), .B1(n12314), .B2(n11858), .ZN(
        n3254) );
  OAI22_X1 U2010 ( .A1(n12364), .A2(n12519), .B1(n12359), .B2(n11859), .ZN(
        n3475) );
  OAI22_X1 U2011 ( .A1(n12364), .A2(n12516), .B1(n12359), .B2(n11860), .ZN(
        n3476) );
  OAI22_X1 U2012 ( .A1(n12364), .A2(n12513), .B1(n12359), .B2(n11861), .ZN(
        n3477) );
  OAI22_X1 U2013 ( .A1(n12364), .A2(n12510), .B1(n12359), .B2(n11862), .ZN(
        n3478) );
  OAI22_X1 U2014 ( .A1(n12382), .A2(n12520), .B1(n12377), .B2(n11863), .ZN(
        n3603) );
  OAI22_X1 U2015 ( .A1(n12382), .A2(n12517), .B1(n12377), .B2(n11864), .ZN(
        n3604) );
  OAI22_X1 U2016 ( .A1(n12382), .A2(n12514), .B1(n12377), .B2(n11865), .ZN(
        n3605) );
  OAI22_X1 U2017 ( .A1(n12382), .A2(n12511), .B1(n12377), .B2(n11866), .ZN(
        n3606) );
  OAI22_X1 U2018 ( .A1(n12175), .A2(n12518), .B1(n1146), .B2(n11867), .ZN(
        n2611) );
  OAI22_X1 U2019 ( .A1(n12173), .A2(n12491), .B1(n1146), .B2(n11868), .ZN(
        n2620) );
  OAI22_X1 U2020 ( .A1(n12173), .A2(n12488), .B1(n1146), .B2(n11869), .ZN(
        n2621) );
  OAI22_X1 U2021 ( .A1(n12173), .A2(n12485), .B1(n1146), .B2(n11870), .ZN(
        n2622) );
  OAI22_X1 U2022 ( .A1(n12172), .A2(n12467), .B1(n1146), .B2(n11871), .ZN(
        n2628) );
  OAI22_X1 U2023 ( .A1(n12172), .A2(n12464), .B1(n1146), .B2(n11872), .ZN(
        n2629) );
  OAI22_X1 U2024 ( .A1(n12171), .A2(n12461), .B1(n12170), .B2(n11873), .ZN(
        n2630) );
  OAI22_X1 U2025 ( .A1(n12171), .A2(n12458), .B1(n12170), .B2(n11874), .ZN(
        n2631) );
  OAI22_X1 U2026 ( .A1(n12171), .A2(n12455), .B1(n12170), .B2(n11875), .ZN(
        n2632) );
  OAI22_X1 U2027 ( .A1(n12171), .A2(n12452), .B1(n12170), .B2(n11876), .ZN(
        n2633) );
  OAI22_X1 U2028 ( .A1(n12171), .A2(n12449), .B1(n12170), .B2(n11877), .ZN(
        n2634) );
  OAI22_X1 U2029 ( .A1(n12193), .A2(n12518), .B1(n1144), .B2(n11878), .ZN(
        n2739) );
  OAI22_X1 U2030 ( .A1(n12191), .A2(n12491), .B1(n1144), .B2(n11879), .ZN(
        n2748) );
  OAI22_X1 U2031 ( .A1(n12191), .A2(n12488), .B1(n1144), .B2(n11880), .ZN(
        n2749) );
  OAI22_X1 U2032 ( .A1(n12191), .A2(n12485), .B1(n1144), .B2(n11881), .ZN(
        n2750) );
  OAI22_X1 U2033 ( .A1(n12190), .A2(n12467), .B1(n1144), .B2(n11882), .ZN(
        n2756) );
  OAI22_X1 U2034 ( .A1(n12190), .A2(n12464), .B1(n1144), .B2(n11883), .ZN(
        n2757) );
  OAI22_X1 U2035 ( .A1(n12189), .A2(n12461), .B1(n12188), .B2(n11884), .ZN(
        n2758) );
  OAI22_X1 U2036 ( .A1(n12189), .A2(n12458), .B1(n12188), .B2(n11885), .ZN(
        n2759) );
  OAI22_X1 U2037 ( .A1(n12189), .A2(n12455), .B1(n12188), .B2(n11886), .ZN(
        n2760) );
  OAI22_X1 U2038 ( .A1(n12189), .A2(n12452), .B1(n12188), .B2(n11887), .ZN(
        n2761) );
  OAI22_X1 U2039 ( .A1(n12189), .A2(n12449), .B1(n12188), .B2(n11888), .ZN(
        n2762) );
  OAI22_X1 U2040 ( .A1(n12211), .A2(n12518), .B1(n12206), .B2(n11889), .ZN(
        n2867) );
  OAI22_X1 U2041 ( .A1(n12209), .A2(n12491), .B1(n12206), .B2(n11890), .ZN(
        n2876) );
  OAI22_X1 U2042 ( .A1(n12209), .A2(n12488), .B1(n12206), .B2(n11891), .ZN(
        n2877) );
  OAI22_X1 U2043 ( .A1(n12209), .A2(n12485), .B1(n12206), .B2(n11892), .ZN(
        n2878) );
  OAI22_X1 U2044 ( .A1(n12208), .A2(n12467), .B1(n12206), .B2(n11893), .ZN(
        n2884) );
  OAI22_X1 U2045 ( .A1(n12208), .A2(n12464), .B1(n12206), .B2(n11894), .ZN(
        n2885) );
  OAI22_X1 U2046 ( .A1(n12207), .A2(n12461), .B1(n12206), .B2(n11895), .ZN(
        n2886) );
  OAI22_X1 U2047 ( .A1(n12207), .A2(n12458), .B1(n12206), .B2(n11896), .ZN(
        n2887) );
  OAI22_X1 U2048 ( .A1(n12207), .A2(n12455), .B1(n12206), .B2(n11897), .ZN(
        n2888) );
  OAI22_X1 U2049 ( .A1(n12207), .A2(n12452), .B1(n12206), .B2(n11898), .ZN(
        n2889) );
  OAI22_X1 U2050 ( .A1(n12207), .A2(n12449), .B1(n12206), .B2(n11899), .ZN(
        n2890) );
  OAI22_X1 U2051 ( .A1(n12245), .A2(n12491), .B1(n12242), .B2(n11900), .ZN(
        n3004) );
  OAI22_X1 U2052 ( .A1(n12245), .A2(n12488), .B1(n12242), .B2(n11901), .ZN(
        n3005) );
  OAI22_X1 U2053 ( .A1(n12245), .A2(n12485), .B1(n12242), .B2(n11902), .ZN(
        n3006) );
  OAI22_X1 U2054 ( .A1(n12245), .A2(n12479), .B1(n12242), .B2(n11903), .ZN(
        n3008) );
  OAI22_X1 U2055 ( .A1(n12244), .A2(n12476), .B1(n12242), .B2(n11904), .ZN(
        n3009) );
  OAI22_X1 U2056 ( .A1(n12244), .A2(n12473), .B1(n12242), .B2(n11905), .ZN(
        n3010) );
  OAI22_X1 U2057 ( .A1(n12244), .A2(n12470), .B1(n12242), .B2(n11906), .ZN(
        n3011) );
  OAI22_X1 U2058 ( .A1(n12244), .A2(n12467), .B1(n12242), .B2(n11907), .ZN(
        n3012) );
  OAI22_X1 U2059 ( .A1(n12244), .A2(n12464), .B1(n12242), .B2(n11908), .ZN(
        n3013) );
  OAI22_X1 U2060 ( .A1(n12243), .A2(n12461), .B1(n12242), .B2(n11909), .ZN(
        n3014) );
  OAI22_X1 U2061 ( .A1(n12243), .A2(n12458), .B1(n12242), .B2(n11910), .ZN(
        n3015) );
  OAI22_X1 U2062 ( .A1(n12243), .A2(n12449), .B1(n12242), .B2(n11911), .ZN(
        n3018) );
  OAI22_X1 U2063 ( .A1(n12282), .A2(n12507), .B1(n12278), .B2(n11912), .ZN(
        n3127) );
  OAI22_X1 U2064 ( .A1(n12282), .A2(n12504), .B1(n12278), .B2(n11913), .ZN(
        n3128) );
  OAI22_X1 U2065 ( .A1(n12282), .A2(n12501), .B1(n12278), .B2(n11914), .ZN(
        n3129) );
  OAI22_X1 U2066 ( .A1(n12282), .A2(n12498), .B1(n12278), .B2(n11915), .ZN(
        n3130) );
  OAI22_X1 U2067 ( .A1(n12282), .A2(n12495), .B1(n12278), .B2(n11916), .ZN(
        n3131) );
  OAI22_X1 U2068 ( .A1(n12281), .A2(n12492), .B1(n12278), .B2(n11917), .ZN(
        n3132) );
  OAI22_X1 U2069 ( .A1(n12281), .A2(n12489), .B1(n12278), .B2(n11918), .ZN(
        n3133) );
  OAI22_X1 U2070 ( .A1(n12281), .A2(n12486), .B1(n12278), .B2(n11919), .ZN(
        n3134) );
  OAI22_X1 U2071 ( .A1(n12281), .A2(n12483), .B1(n12278), .B2(n11920), .ZN(
        n3135) );
  OAI22_X1 U2072 ( .A1(n12281), .A2(n12480), .B1(n12278), .B2(n11921), .ZN(
        n3136) );
  OAI22_X1 U2073 ( .A1(n12280), .A2(n12477), .B1(n12278), .B2(n11922), .ZN(
        n3137) );
  OAI22_X1 U2074 ( .A1(n12280), .A2(n12474), .B1(n12278), .B2(n11923), .ZN(
        n3138) );
  OAI22_X1 U2075 ( .A1(n12318), .A2(n12507), .B1(n12314), .B2(n11924), .ZN(
        n3255) );
  OAI22_X1 U2076 ( .A1(n12318), .A2(n12504), .B1(n12314), .B2(n11925), .ZN(
        n3256) );
  OAI22_X1 U2077 ( .A1(n12318), .A2(n12501), .B1(n12314), .B2(n11926), .ZN(
        n3257) );
  OAI22_X1 U2078 ( .A1(n12318), .A2(n12498), .B1(n12314), .B2(n11927), .ZN(
        n3258) );
  OAI22_X1 U2079 ( .A1(n12318), .A2(n12495), .B1(n12314), .B2(n11928), .ZN(
        n3259) );
  OAI22_X1 U2080 ( .A1(n12317), .A2(n12492), .B1(n12314), .B2(n11929), .ZN(
        n3260) );
  OAI22_X1 U2081 ( .A1(n12317), .A2(n12489), .B1(n12314), .B2(n11930), .ZN(
        n3261) );
  OAI22_X1 U2082 ( .A1(n12317), .A2(n12486), .B1(n12314), .B2(n11931), .ZN(
        n3262) );
  OAI22_X1 U2083 ( .A1(n12317), .A2(n12483), .B1(n12314), .B2(n11932), .ZN(
        n3263) );
  OAI22_X1 U2084 ( .A1(n12317), .A2(n12480), .B1(n12314), .B2(n11933), .ZN(
        n3264) );
  OAI22_X1 U2085 ( .A1(n12316), .A2(n12477), .B1(n12314), .B2(n11934), .ZN(
        n3265) );
  OAI22_X1 U2086 ( .A1(n12316), .A2(n12474), .B1(n12314), .B2(n11935), .ZN(
        n3266) );
  OAI22_X1 U2087 ( .A1(n12363), .A2(n12507), .B1(n12359), .B2(n11936), .ZN(
        n3479) );
  OAI22_X1 U2088 ( .A1(n12363), .A2(n12504), .B1(n12359), .B2(n11937), .ZN(
        n3480) );
  OAI22_X1 U2089 ( .A1(n12363), .A2(n12501), .B1(n12359), .B2(n11938), .ZN(
        n3481) );
  OAI22_X1 U2090 ( .A1(n12363), .A2(n12498), .B1(n12359), .B2(n11939), .ZN(
        n3482) );
  OAI22_X1 U2091 ( .A1(n12363), .A2(n12495), .B1(n12359), .B2(n11940), .ZN(
        n3483) );
  OAI22_X1 U2092 ( .A1(n12362), .A2(n12492), .B1(n12359), .B2(n11941), .ZN(
        n3484) );
  OAI22_X1 U2093 ( .A1(n12362), .A2(n12489), .B1(n12359), .B2(n11942), .ZN(
        n3485) );
  OAI22_X1 U2094 ( .A1(n12362), .A2(n12486), .B1(n12359), .B2(n11943), .ZN(
        n3486) );
  OAI22_X1 U2095 ( .A1(n12362), .A2(n12483), .B1(n12359), .B2(n11944), .ZN(
        n3487) );
  OAI22_X1 U2096 ( .A1(n12362), .A2(n12480), .B1(n12359), .B2(n11945), .ZN(
        n3488) );
  OAI22_X1 U2097 ( .A1(n12361), .A2(n12477), .B1(n12359), .B2(n11946), .ZN(
        n3489) );
  OAI22_X1 U2098 ( .A1(n12361), .A2(n12474), .B1(n12359), .B2(n11947), .ZN(
        n3490) );
  OAI22_X1 U2099 ( .A1(n12381), .A2(n12508), .B1(n12377), .B2(n11948), .ZN(
        n3607) );
  OAI22_X1 U2100 ( .A1(n12381), .A2(n12505), .B1(n12377), .B2(n11949), .ZN(
        n3608) );
  OAI22_X1 U2101 ( .A1(n12381), .A2(n12502), .B1(n12377), .B2(n11950), .ZN(
        n3609) );
  OAI22_X1 U2102 ( .A1(n12381), .A2(n12499), .B1(n12377), .B2(n11951), .ZN(
        n3610) );
  OAI22_X1 U2103 ( .A1(n12381), .A2(n12496), .B1(n12377), .B2(n11952), .ZN(
        n3611) );
  OAI22_X1 U2104 ( .A1(n12380), .A2(n12493), .B1(n12377), .B2(n11953), .ZN(
        n3612) );
  OAI22_X1 U2105 ( .A1(n12380), .A2(n12490), .B1(n12377), .B2(n11954), .ZN(
        n3613) );
  OAI22_X1 U2106 ( .A1(n12380), .A2(n12487), .B1(n12377), .B2(n11955), .ZN(
        n3614) );
  OAI22_X1 U2107 ( .A1(n12380), .A2(n12484), .B1(n12377), .B2(n11956), .ZN(
        n3615) );
  OAI22_X1 U2108 ( .A1(n12380), .A2(n12481), .B1(n12377), .B2(n11957), .ZN(
        n3616) );
  OAI22_X1 U2109 ( .A1(n12379), .A2(n12478), .B1(n12377), .B2(n11958), .ZN(
        n3617) );
  OAI22_X1 U2110 ( .A1(n12379), .A2(n12475), .B1(n12377), .B2(n11959), .ZN(
        n3618) );
  OAI22_X1 U2111 ( .A1(n12186), .A2(n12551), .B1(n12179), .B2(n11528), .ZN(
        n2635) );
  OAI22_X1 U2112 ( .A1(n12186), .A2(n12539), .B1(n12179), .B2(n11529), .ZN(
        n2636) );
  OAI22_X1 U2113 ( .A1(n12185), .A2(n12536), .B1(n12179), .B2(n11530), .ZN(
        n2637) );
  OAI22_X1 U2114 ( .A1(n12185), .A2(n12533), .B1(n12179), .B2(n11531), .ZN(
        n2638) );
  OAI22_X1 U2115 ( .A1(n12185), .A2(n12530), .B1(n12179), .B2(n11532), .ZN(
        n2639) );
  OAI22_X1 U2116 ( .A1(n12185), .A2(n12527), .B1(n12179), .B2(n11533), .ZN(
        n2640) );
  OAI22_X1 U2117 ( .A1(n12185), .A2(n12524), .B1(n12179), .B2(n11534), .ZN(
        n2641) );
  OAI22_X1 U2118 ( .A1(n12184), .A2(n12521), .B1(n12179), .B2(n11535), .ZN(
        n2642) );
  OAI22_X1 U2119 ( .A1(n12184), .A2(n12518), .B1(n12179), .B2(n11536), .ZN(
        n2643) );
  OAI22_X1 U2120 ( .A1(n12184), .A2(n12515), .B1(n12179), .B2(n11537), .ZN(
        n2644) );
  OAI22_X1 U2121 ( .A1(n12184), .A2(n12512), .B1(n12179), .B2(n11538), .ZN(
        n2645) );
  OAI22_X1 U2122 ( .A1(n12184), .A2(n12509), .B1(n12179), .B2(n11539), .ZN(
        n2646) );
  OAI22_X1 U2123 ( .A1(n12183), .A2(n12506), .B1(n1145), .B2(n11540), .ZN(
        n2647) );
  OAI22_X1 U2124 ( .A1(n12183), .A2(n12503), .B1(n1145), .B2(n11541), .ZN(
        n2648) );
  OAI22_X1 U2125 ( .A1(n12183), .A2(n12500), .B1(n1145), .B2(n11542), .ZN(
        n2649) );
  OAI22_X1 U2126 ( .A1(n12183), .A2(n12497), .B1(n1145), .B2(n11543), .ZN(
        n2650) );
  OAI22_X1 U2127 ( .A1(n12183), .A2(n12494), .B1(n12179), .B2(n11544), .ZN(
        n2651) );
  OAI22_X1 U2128 ( .A1(n12182), .A2(n12491), .B1(n12179), .B2(n11545), .ZN(
        n2652) );
  OAI22_X1 U2129 ( .A1(n12182), .A2(n12488), .B1(n12179), .B2(n11546), .ZN(
        n2653) );
  OAI22_X1 U2130 ( .A1(n12182), .A2(n12485), .B1(n12179), .B2(n11547), .ZN(
        n2654) );
  OAI22_X1 U2131 ( .A1(n12182), .A2(n12482), .B1(n12179), .B2(n11548), .ZN(
        n2655) );
  OAI22_X1 U2132 ( .A1(n12182), .A2(n12479), .B1(n12179), .B2(n11549), .ZN(
        n2656) );
  OAI22_X1 U2133 ( .A1(n12204), .A2(n12551), .B1(n12197), .B2(n11550), .ZN(
        n2763) );
  OAI22_X1 U2134 ( .A1(n12204), .A2(n12539), .B1(n12197), .B2(n11551), .ZN(
        n2764) );
  OAI22_X1 U2135 ( .A1(n12203), .A2(n12536), .B1(n12197), .B2(n11552), .ZN(
        n2765) );
  OAI22_X1 U2136 ( .A1(n12203), .A2(n12533), .B1(n12197), .B2(n11553), .ZN(
        n2766) );
  OAI22_X1 U2137 ( .A1(n12203), .A2(n12530), .B1(n12197), .B2(n11554), .ZN(
        n2767) );
  OAI22_X1 U2138 ( .A1(n12203), .A2(n12527), .B1(n12197), .B2(n11555), .ZN(
        n2768) );
  OAI22_X1 U2139 ( .A1(n12203), .A2(n12524), .B1(n12197), .B2(n11556), .ZN(
        n2769) );
  OAI22_X1 U2140 ( .A1(n12202), .A2(n12521), .B1(n12197), .B2(n11557), .ZN(
        n2770) );
  OAI22_X1 U2141 ( .A1(n12202), .A2(n12518), .B1(n12197), .B2(n11558), .ZN(
        n2771) );
  OAI22_X1 U2142 ( .A1(n12202), .A2(n12515), .B1(n12197), .B2(n11559), .ZN(
        n2772) );
  OAI22_X1 U2143 ( .A1(n12202), .A2(n12512), .B1(n12197), .B2(n11560), .ZN(
        n2773) );
  OAI22_X1 U2144 ( .A1(n12202), .A2(n12509), .B1(n12197), .B2(n11561), .ZN(
        n2774) );
  OAI22_X1 U2145 ( .A1(n12201), .A2(n12506), .B1(n1143), .B2(n11562), .ZN(
        n2775) );
  OAI22_X1 U2146 ( .A1(n12201), .A2(n12503), .B1(n1143), .B2(n11563), .ZN(
        n2776) );
  OAI22_X1 U2147 ( .A1(n12201), .A2(n12500), .B1(n1143), .B2(n11564), .ZN(
        n2777) );
  OAI22_X1 U2148 ( .A1(n12201), .A2(n12497), .B1(n1143), .B2(n11565), .ZN(
        n2778) );
  OAI22_X1 U2149 ( .A1(n12201), .A2(n12494), .B1(n12197), .B2(n11566), .ZN(
        n2779) );
  OAI22_X1 U2150 ( .A1(n12200), .A2(n12491), .B1(n12197), .B2(n11567), .ZN(
        n2780) );
  OAI22_X1 U2151 ( .A1(n12200), .A2(n12488), .B1(n12197), .B2(n11568), .ZN(
        n2781) );
  OAI22_X1 U2152 ( .A1(n12200), .A2(n12485), .B1(n12197), .B2(n11569), .ZN(
        n2782) );
  OAI22_X1 U2153 ( .A1(n12200), .A2(n12482), .B1(n12197), .B2(n11570), .ZN(
        n2783) );
  OAI22_X1 U2154 ( .A1(n12200), .A2(n12479), .B1(n12197), .B2(n11571), .ZN(
        n2784) );
  OAI22_X1 U2155 ( .A1(n12222), .A2(n12551), .B1(n12215), .B2(n11572), .ZN(
        n2891) );
  OAI22_X1 U2156 ( .A1(n12222), .A2(n12539), .B1(n12215), .B2(n11573), .ZN(
        n2892) );
  OAI22_X1 U2157 ( .A1(n12221), .A2(n12536), .B1(n12215), .B2(n11574), .ZN(
        n2893) );
  OAI22_X1 U2158 ( .A1(n12221), .A2(n12533), .B1(n12215), .B2(n11575), .ZN(
        n2894) );
  OAI22_X1 U2159 ( .A1(n12221), .A2(n12530), .B1(n12215), .B2(n11576), .ZN(
        n2895) );
  OAI22_X1 U2160 ( .A1(n12221), .A2(n12527), .B1(n12215), .B2(n11577), .ZN(
        n2896) );
  OAI22_X1 U2161 ( .A1(n12221), .A2(n12524), .B1(n12215), .B2(n11578), .ZN(
        n2897) );
  OAI22_X1 U2162 ( .A1(n12220), .A2(n12521), .B1(n12215), .B2(n11579), .ZN(
        n2898) );
  OAI22_X1 U2163 ( .A1(n12220), .A2(n12518), .B1(n12215), .B2(n11580), .ZN(
        n2899) );
  OAI22_X1 U2164 ( .A1(n12220), .A2(n12515), .B1(n12215), .B2(n11581), .ZN(
        n2900) );
  OAI22_X1 U2165 ( .A1(n12220), .A2(n12512), .B1(n12215), .B2(n11582), .ZN(
        n2901) );
  OAI22_X1 U2166 ( .A1(n12220), .A2(n12509), .B1(n12215), .B2(n11583), .ZN(
        n2902) );
  OAI22_X1 U2167 ( .A1(n12219), .A2(n12506), .B1(n1141), .B2(n11584), .ZN(
        n2903) );
  OAI22_X1 U2168 ( .A1(n12219), .A2(n12503), .B1(n1141), .B2(n11585), .ZN(
        n2904) );
  OAI22_X1 U2169 ( .A1(n12219), .A2(n12500), .B1(n1141), .B2(n11586), .ZN(
        n2905) );
  OAI22_X1 U2170 ( .A1(n12219), .A2(n12497), .B1(n1141), .B2(n11587), .ZN(
        n2906) );
  OAI22_X1 U2171 ( .A1(n12219), .A2(n12494), .B1(n12215), .B2(n11588), .ZN(
        n2907) );
  OAI22_X1 U2172 ( .A1(n12218), .A2(n12491), .B1(n12215), .B2(n11589), .ZN(
        n2908) );
  OAI22_X1 U2173 ( .A1(n12218), .A2(n12488), .B1(n12215), .B2(n11590), .ZN(
        n2909) );
  OAI22_X1 U2174 ( .A1(n12218), .A2(n12485), .B1(n12215), .B2(n11591), .ZN(
        n2910) );
  OAI22_X1 U2175 ( .A1(n12218), .A2(n12482), .B1(n12215), .B2(n11592), .ZN(
        n2911) );
  OAI22_X1 U2176 ( .A1(n12218), .A2(n12479), .B1(n12215), .B2(n11593), .ZN(
        n2912) );
  OAI22_X1 U2177 ( .A1(n12258), .A2(n12551), .B1(n12251), .B2(n11594), .ZN(
        n3019) );
  OAI22_X1 U2178 ( .A1(n12258), .A2(n12539), .B1(n12251), .B2(n11595), .ZN(
        n3020) );
  OAI22_X1 U2179 ( .A1(n12257), .A2(n12536), .B1(n12251), .B2(n11596), .ZN(
        n3021) );
  OAI22_X1 U2180 ( .A1(n12257), .A2(n12533), .B1(n12251), .B2(n11597), .ZN(
        n3022) );
  OAI22_X1 U2181 ( .A1(n12257), .A2(n12530), .B1(n12251), .B2(n11598), .ZN(
        n3023) );
  OAI22_X1 U2182 ( .A1(n12257), .A2(n12527), .B1(n12251), .B2(n11599), .ZN(
        n3024) );
  OAI22_X1 U2183 ( .A1(n12257), .A2(n12524), .B1(n12251), .B2(n11600), .ZN(
        n3025) );
  OAI22_X1 U2184 ( .A1(n12256), .A2(n12521), .B1(n12251), .B2(n11601), .ZN(
        n3026) );
  OAI22_X1 U2185 ( .A1(n12256), .A2(n12518), .B1(n12251), .B2(n11602), .ZN(
        n3027) );
  OAI22_X1 U2186 ( .A1(n12256), .A2(n12515), .B1(n12251), .B2(n11603), .ZN(
        n3028) );
  OAI22_X1 U2187 ( .A1(n12256), .A2(n12512), .B1(n12251), .B2(n11604), .ZN(
        n3029) );
  OAI22_X1 U2188 ( .A1(n12256), .A2(n12509), .B1(n12251), .B2(n11605), .ZN(
        n3030) );
  OAI22_X1 U2189 ( .A1(n12255), .A2(n12506), .B1(n1137), .B2(n11606), .ZN(
        n3031) );
  OAI22_X1 U2190 ( .A1(n12255), .A2(n12503), .B1(n1137), .B2(n11607), .ZN(
        n3032) );
  OAI22_X1 U2191 ( .A1(n12255), .A2(n12500), .B1(n1137), .B2(n11608), .ZN(
        n3033) );
  OAI22_X1 U2192 ( .A1(n12255), .A2(n12497), .B1(n1137), .B2(n11609), .ZN(
        n3034) );
  OAI22_X1 U2193 ( .A1(n12255), .A2(n12494), .B1(n12251), .B2(n11610), .ZN(
        n3035) );
  OAI22_X1 U2194 ( .A1(n12254), .A2(n12491), .B1(n12251), .B2(n11611), .ZN(
        n3036) );
  OAI22_X1 U2195 ( .A1(n12254), .A2(n12488), .B1(n12251), .B2(n11612), .ZN(
        n3037) );
  OAI22_X1 U2196 ( .A1(n12254), .A2(n12485), .B1(n12251), .B2(n11613), .ZN(
        n3038) );
  OAI22_X1 U2197 ( .A1(n12254), .A2(n12482), .B1(n12251), .B2(n11614), .ZN(
        n3039) );
  OAI22_X1 U2198 ( .A1(n12254), .A2(n12479), .B1(n12251), .B2(n11615), .ZN(
        n3040) );
  OAI22_X1 U2199 ( .A1(n12294), .A2(n12552), .B1(n12287), .B2(n11616), .ZN(
        n3147) );
  OAI22_X1 U2200 ( .A1(n12294), .A2(n12540), .B1(n12287), .B2(n11617), .ZN(
        n3148) );
  OAI22_X1 U2201 ( .A1(n12293), .A2(n12537), .B1(n12287), .B2(n11618), .ZN(
        n3149) );
  OAI22_X1 U2202 ( .A1(n12293), .A2(n12534), .B1(n12287), .B2(n11619), .ZN(
        n3150) );
  OAI22_X1 U2203 ( .A1(n12293), .A2(n12531), .B1(n12287), .B2(n11620), .ZN(
        n3151) );
  OAI22_X1 U2204 ( .A1(n12293), .A2(n12528), .B1(n12287), .B2(n11621), .ZN(
        n3152) );
  OAI22_X1 U2205 ( .A1(n12293), .A2(n12525), .B1(n12287), .B2(n11622), .ZN(
        n3153) );
  OAI22_X1 U2206 ( .A1(n12292), .A2(n12522), .B1(n12287), .B2(n11623), .ZN(
        n3154) );
  OAI22_X1 U2207 ( .A1(n12292), .A2(n12519), .B1(n12287), .B2(n11624), .ZN(
        n3155) );
  OAI22_X1 U2208 ( .A1(n12292), .A2(n12516), .B1(n12287), .B2(n11625), .ZN(
        n3156) );
  OAI22_X1 U2209 ( .A1(n12292), .A2(n12513), .B1(n12287), .B2(n11626), .ZN(
        n3157) );
  OAI22_X1 U2210 ( .A1(n12292), .A2(n12510), .B1(n12287), .B2(n11627), .ZN(
        n3158) );
  OAI22_X1 U2211 ( .A1(n12291), .A2(n12507), .B1(n1132), .B2(n11628), .ZN(
        n3159) );
  OAI22_X1 U2212 ( .A1(n12291), .A2(n12504), .B1(n1132), .B2(n11629), .ZN(
        n3160) );
  OAI22_X1 U2213 ( .A1(n12291), .A2(n12501), .B1(n1132), .B2(n11630), .ZN(
        n3161) );
  OAI22_X1 U2214 ( .A1(n12291), .A2(n12498), .B1(n1132), .B2(n11631), .ZN(
        n3162) );
  OAI22_X1 U2215 ( .A1(n12291), .A2(n12495), .B1(n12287), .B2(n11632), .ZN(
        n3163) );
  OAI22_X1 U2216 ( .A1(n12290), .A2(n12492), .B1(n12287), .B2(n11633), .ZN(
        n3164) );
  OAI22_X1 U2217 ( .A1(n12290), .A2(n12489), .B1(n12287), .B2(n11634), .ZN(
        n3165) );
  OAI22_X1 U2218 ( .A1(n12290), .A2(n12486), .B1(n12287), .B2(n11635), .ZN(
        n3166) );
  OAI22_X1 U2219 ( .A1(n12290), .A2(n12483), .B1(n12287), .B2(n11636), .ZN(
        n3167) );
  OAI22_X1 U2220 ( .A1(n12290), .A2(n12480), .B1(n12287), .B2(n11637), .ZN(
        n3168) );
  OAI22_X1 U2221 ( .A1(n12330), .A2(n12552), .B1(n12323), .B2(n11638), .ZN(
        n3275) );
  OAI22_X1 U2222 ( .A1(n12330), .A2(n12540), .B1(n12323), .B2(n11639), .ZN(
        n3276) );
  OAI22_X1 U2223 ( .A1(n12329), .A2(n12537), .B1(n12323), .B2(n11640), .ZN(
        n3277) );
  OAI22_X1 U2224 ( .A1(n12329), .A2(n12534), .B1(n12323), .B2(n11641), .ZN(
        n3278) );
  OAI22_X1 U2225 ( .A1(n12329), .A2(n12531), .B1(n12323), .B2(n11642), .ZN(
        n3279) );
  OAI22_X1 U2226 ( .A1(n12329), .A2(n12528), .B1(n12323), .B2(n11643), .ZN(
        n3280) );
  OAI22_X1 U2227 ( .A1(n12329), .A2(n12525), .B1(n12323), .B2(n11644), .ZN(
        n3281) );
  OAI22_X1 U2228 ( .A1(n12328), .A2(n12522), .B1(n12323), .B2(n11645), .ZN(
        n3282) );
  OAI22_X1 U2229 ( .A1(n12328), .A2(n12519), .B1(n12323), .B2(n11646), .ZN(
        n3283) );
  OAI22_X1 U2230 ( .A1(n12328), .A2(n12516), .B1(n12323), .B2(n11647), .ZN(
        n3284) );
  OAI22_X1 U2231 ( .A1(n12328), .A2(n12513), .B1(n12323), .B2(n11648), .ZN(
        n3285) );
  OAI22_X1 U2232 ( .A1(n12328), .A2(n12510), .B1(n12323), .B2(n11649), .ZN(
        n3286) );
  OAI22_X1 U2233 ( .A1(n12327), .A2(n12507), .B1(n1128), .B2(n11650), .ZN(
        n3287) );
  OAI22_X1 U2234 ( .A1(n12327), .A2(n12504), .B1(n1128), .B2(n11651), .ZN(
        n3288) );
  OAI22_X1 U2235 ( .A1(n12327), .A2(n12501), .B1(n1128), .B2(n11652), .ZN(
        n3289) );
  OAI22_X1 U2236 ( .A1(n12327), .A2(n12498), .B1(n1128), .B2(n11653), .ZN(
        n3290) );
  OAI22_X1 U2237 ( .A1(n12327), .A2(n12495), .B1(n12323), .B2(n11654), .ZN(
        n3291) );
  OAI22_X1 U2238 ( .A1(n12326), .A2(n12492), .B1(n12323), .B2(n11655), .ZN(
        n3292) );
  OAI22_X1 U2239 ( .A1(n12326), .A2(n12489), .B1(n12323), .B2(n11656), .ZN(
        n3293) );
  OAI22_X1 U2240 ( .A1(n12326), .A2(n12486), .B1(n12323), .B2(n11657), .ZN(
        n3294) );
  OAI22_X1 U2241 ( .A1(n12326), .A2(n12483), .B1(n12323), .B2(n11658), .ZN(
        n3295) );
  OAI22_X1 U2242 ( .A1(n12326), .A2(n12480), .B1(n12323), .B2(n11659), .ZN(
        n3296) );
  OAI22_X1 U2243 ( .A1(n12357), .A2(n12552), .B1(n12350), .B2(n11660), .ZN(
        n3435) );
  OAI22_X1 U2244 ( .A1(n12357), .A2(n12540), .B1(n12350), .B2(n11661), .ZN(
        n3436) );
  OAI22_X1 U2245 ( .A1(n12356), .A2(n12537), .B1(n12350), .B2(n11662), .ZN(
        n3437) );
  OAI22_X1 U2246 ( .A1(n12356), .A2(n12534), .B1(n12350), .B2(n11663), .ZN(
        n3438) );
  OAI22_X1 U2247 ( .A1(n12356), .A2(n12531), .B1(n12350), .B2(n11664), .ZN(
        n3439) );
  OAI22_X1 U2248 ( .A1(n12356), .A2(n12528), .B1(n12350), .B2(n11665), .ZN(
        n3440) );
  OAI22_X1 U2249 ( .A1(n12356), .A2(n12525), .B1(n12350), .B2(n11666), .ZN(
        n3441) );
  OAI22_X1 U2250 ( .A1(n12355), .A2(n12522), .B1(n12350), .B2(n11667), .ZN(
        n3442) );
  OAI22_X1 U2251 ( .A1(n12355), .A2(n12519), .B1(n12350), .B2(n11668), .ZN(
        n3443) );
  OAI22_X1 U2252 ( .A1(n12355), .A2(n12516), .B1(n12350), .B2(n11669), .ZN(
        n3444) );
  OAI22_X1 U2253 ( .A1(n12355), .A2(n12513), .B1(n12350), .B2(n11670), .ZN(
        n3445) );
  OAI22_X1 U2254 ( .A1(n12355), .A2(n12510), .B1(n12350), .B2(n11671), .ZN(
        n3446) );
  OAI22_X1 U2255 ( .A1(n12354), .A2(n12507), .B1(n1124), .B2(n11672), .ZN(
        n3447) );
  OAI22_X1 U2256 ( .A1(n12354), .A2(n12504), .B1(n1124), .B2(n11673), .ZN(
        n3448) );
  OAI22_X1 U2257 ( .A1(n12354), .A2(n12501), .B1(n1124), .B2(n11674), .ZN(
        n3449) );
  OAI22_X1 U2258 ( .A1(n12354), .A2(n12498), .B1(n1124), .B2(n11675), .ZN(
        n3450) );
  OAI22_X1 U2259 ( .A1(n12354), .A2(n12495), .B1(n12350), .B2(n11676), .ZN(
        n3451) );
  OAI22_X1 U2260 ( .A1(n12353), .A2(n12492), .B1(n12350), .B2(n11677), .ZN(
        n3452) );
  OAI22_X1 U2261 ( .A1(n12353), .A2(n12489), .B1(n12350), .B2(n11678), .ZN(
        n3453) );
  OAI22_X1 U2262 ( .A1(n12353), .A2(n12486), .B1(n12350), .B2(n11679), .ZN(
        n3454) );
  OAI22_X1 U2263 ( .A1(n12353), .A2(n12483), .B1(n12350), .B2(n11680), .ZN(
        n3455) );
  OAI22_X1 U2264 ( .A1(n12353), .A2(n12480), .B1(n12350), .B2(n11681), .ZN(
        n3456) );
  OAI22_X1 U2265 ( .A1(n12375), .A2(n12553), .B1(n12368), .B2(n11682), .ZN(
        n3563) );
  OAI22_X1 U2266 ( .A1(n12375), .A2(n12541), .B1(n12368), .B2(n11683), .ZN(
        n3564) );
  OAI22_X1 U2267 ( .A1(n12374), .A2(n12538), .B1(n12368), .B2(n11684), .ZN(
        n3565) );
  OAI22_X1 U2268 ( .A1(n12374), .A2(n12535), .B1(n12368), .B2(n11685), .ZN(
        n3566) );
  OAI22_X1 U2269 ( .A1(n12374), .A2(n12532), .B1(n12368), .B2(n11686), .ZN(
        n3567) );
  OAI22_X1 U2270 ( .A1(n12374), .A2(n12529), .B1(n12368), .B2(n11687), .ZN(
        n3568) );
  OAI22_X1 U2271 ( .A1(n12374), .A2(n12526), .B1(n12368), .B2(n11688), .ZN(
        n3569) );
  OAI22_X1 U2272 ( .A1(n12373), .A2(n12523), .B1(n12368), .B2(n11689), .ZN(
        n3570) );
  OAI22_X1 U2273 ( .A1(n12373), .A2(n12520), .B1(n12368), .B2(n11690), .ZN(
        n3571) );
  OAI22_X1 U2274 ( .A1(n12373), .A2(n12517), .B1(n12368), .B2(n11691), .ZN(
        n3572) );
  OAI22_X1 U2275 ( .A1(n12373), .A2(n12514), .B1(n12368), .B2(n11692), .ZN(
        n3573) );
  OAI22_X1 U2276 ( .A1(n12373), .A2(n12511), .B1(n12368), .B2(n11693), .ZN(
        n3574) );
  OAI22_X1 U2277 ( .A1(n12372), .A2(n12508), .B1(n1122), .B2(n11694), .ZN(
        n3575) );
  OAI22_X1 U2278 ( .A1(n12372), .A2(n12505), .B1(n1122), .B2(n11695), .ZN(
        n3576) );
  OAI22_X1 U2279 ( .A1(n12372), .A2(n12502), .B1(n1122), .B2(n11696), .ZN(
        n3577) );
  OAI22_X1 U2280 ( .A1(n12372), .A2(n12499), .B1(n1122), .B2(n11697), .ZN(
        n3578) );
  OAI22_X1 U2281 ( .A1(n12372), .A2(n12496), .B1(n12368), .B2(n11698), .ZN(
        n3579) );
  OAI22_X1 U2282 ( .A1(n12371), .A2(n12493), .B1(n12368), .B2(n11699), .ZN(
        n3580) );
  OAI22_X1 U2283 ( .A1(n12371), .A2(n12490), .B1(n12368), .B2(n11700), .ZN(
        n3581) );
  OAI22_X1 U2284 ( .A1(n12371), .A2(n12487), .B1(n12368), .B2(n11701), .ZN(
        n3582) );
  OAI22_X1 U2285 ( .A1(n12371), .A2(n12484), .B1(n12368), .B2(n11702), .ZN(
        n3583) );
  OAI22_X1 U2286 ( .A1(n12371), .A2(n12481), .B1(n12368), .B2(n11703), .ZN(
        n3584) );
  OAI22_X1 U2287 ( .A1(n12177), .A2(n12551), .B1(n9920), .B2(n12170), .ZN(
        n2603) );
  OAI22_X1 U2288 ( .A1(n12177), .A2(n12539), .B1(n9921), .B2(n12170), .ZN(
        n2604) );
  OAI22_X1 U2289 ( .A1(n12176), .A2(n12536), .B1(n9922), .B2(n12170), .ZN(
        n2605) );
  OAI22_X1 U2290 ( .A1(n12176), .A2(n12533), .B1(n9923), .B2(n12170), .ZN(
        n2606) );
  OAI22_X1 U2291 ( .A1(n12176), .A2(n12530), .B1(n9924), .B2(n12170), .ZN(
        n2607) );
  OAI22_X1 U2292 ( .A1(n12176), .A2(n12527), .B1(n9925), .B2(n12170), .ZN(
        n2608) );
  OAI22_X1 U2293 ( .A1(n12176), .A2(n12524), .B1(n9926), .B2(n12170), .ZN(
        n2609) );
  OAI22_X1 U2294 ( .A1(n12175), .A2(n12521), .B1(n9927), .B2(n12170), .ZN(
        n2610) );
  OAI22_X1 U2295 ( .A1(n12173), .A2(n12482), .B1(n9984), .B2(n12170), .ZN(
        n2623) );
  OAI22_X1 U2296 ( .A1(n12172), .A2(n12476), .B1(n9986), .B2(n1146), .ZN(n2625) );
  OAI22_X1 U2297 ( .A1(n12172), .A2(n12473), .B1(n9987), .B2(n1146), .ZN(n2626) );
  OAI22_X1 U2298 ( .A1(n12172), .A2(n12470), .B1(n9988), .B2(n1146), .ZN(n2627) );
  OAI22_X1 U2299 ( .A1(n12195), .A2(n12551), .B1(n9928), .B2(n12188), .ZN(
        n2731) );
  OAI22_X1 U2300 ( .A1(n12195), .A2(n12539), .B1(n9929), .B2(n12188), .ZN(
        n2732) );
  OAI22_X1 U2301 ( .A1(n12194), .A2(n12536), .B1(n9930), .B2(n12188), .ZN(
        n2733) );
  OAI22_X1 U2302 ( .A1(n12194), .A2(n12533), .B1(n9931), .B2(n12188), .ZN(
        n2734) );
  OAI22_X1 U2303 ( .A1(n12194), .A2(n12530), .B1(n9932), .B2(n12188), .ZN(
        n2735) );
  OAI22_X1 U2304 ( .A1(n12194), .A2(n12527), .B1(n9933), .B2(n12188), .ZN(
        n2736) );
  OAI22_X1 U2305 ( .A1(n12194), .A2(n12524), .B1(n9934), .B2(n12188), .ZN(
        n2737) );
  OAI22_X1 U2306 ( .A1(n12193), .A2(n12521), .B1(n9935), .B2(n12188), .ZN(
        n2738) );
  OAI22_X1 U2307 ( .A1(n12191), .A2(n12482), .B1(n9989), .B2(n12188), .ZN(
        n2751) );
  OAI22_X1 U2308 ( .A1(n12190), .A2(n12476), .B1(n9991), .B2(n1144), .ZN(n2753) );
  OAI22_X1 U2309 ( .A1(n12190), .A2(n12473), .B1(n9992), .B2(n1144), .ZN(n2754) );
  OAI22_X1 U2310 ( .A1(n12190), .A2(n12470), .B1(n9993), .B2(n1144), .ZN(n2755) );
  OAI22_X1 U2311 ( .A1(n12213), .A2(n12551), .B1(n9936), .B2(n12206), .ZN(
        n2859) );
  OAI22_X1 U2312 ( .A1(n12213), .A2(n12539), .B1(n9937), .B2(n12206), .ZN(
        n2860) );
  OAI22_X1 U2313 ( .A1(n12212), .A2(n12536), .B1(n9938), .B2(n12206), .ZN(
        n2861) );
  OAI22_X1 U2314 ( .A1(n12212), .A2(n12533), .B1(n9939), .B2(n1142), .ZN(n2862) );
  OAI22_X1 U2315 ( .A1(n12212), .A2(n12530), .B1(n9940), .B2(n1142), .ZN(n2863) );
  OAI22_X1 U2316 ( .A1(n12212), .A2(n12527), .B1(n9941), .B2(n12206), .ZN(
        n2864) );
  OAI22_X1 U2317 ( .A1(n12212), .A2(n12524), .B1(n9942), .B2(n1142), .ZN(n2865) );
  OAI22_X1 U2318 ( .A1(n12211), .A2(n12521), .B1(n9943), .B2(n12206), .ZN(
        n2866) );
  OAI22_X1 U2319 ( .A1(n12209), .A2(n12482), .B1(n9994), .B2(n1142), .ZN(n2879) );
  OAI22_X1 U2320 ( .A1(n12208), .A2(n12476), .B1(n9996), .B2(n1142), .ZN(n2881) );
  OAI22_X1 U2321 ( .A1(n12208), .A2(n12473), .B1(n9997), .B2(n1142), .ZN(n2882) );
  OAI22_X1 U2322 ( .A1(n12208), .A2(n12470), .B1(n9998), .B2(n1142), .ZN(n2883) );
  OAI22_X1 U2323 ( .A1(n12249), .A2(n12551), .B1(n9944), .B2(n12242), .ZN(
        n2987) );
  OAI22_X1 U2324 ( .A1(n12249), .A2(n12539), .B1(n9945), .B2(n12242), .ZN(
        n2988) );
  OAI22_X1 U2325 ( .A1(n12248), .A2(n12536), .B1(n9946), .B2(n1138), .ZN(n2989) );
  OAI22_X1 U2326 ( .A1(n12248), .A2(n12533), .B1(n9947), .B2(n1138), .ZN(n2990) );
  OAI22_X1 U2327 ( .A1(n12248), .A2(n12530), .B1(n9948), .B2(n1138), .ZN(n2991) );
  OAI22_X1 U2328 ( .A1(n12248), .A2(n12527), .B1(n9949), .B2(n1138), .ZN(n2992) );
  OAI22_X1 U2329 ( .A1(n12248), .A2(n12524), .B1(n9950), .B2(n1138), .ZN(n2993) );
  OAI22_X1 U2330 ( .A1(n12247), .A2(n12521), .B1(n9951), .B2(n1138), .ZN(n2994) );
  OAI22_X1 U2331 ( .A1(n12245), .A2(n12482), .B1(n9999), .B2(n1138), .ZN(n3007) );
  OAI22_X1 U2332 ( .A1(n12285), .A2(n12552), .B1(n9952), .B2(n12278), .ZN(
        n3115) );
  OAI22_X1 U2333 ( .A1(n12285), .A2(n12540), .B1(n9953), .B2(n12278), .ZN(
        n3116) );
  OAI22_X1 U2334 ( .A1(n12284), .A2(n12537), .B1(n9954), .B2(n1133), .ZN(n3117) );
  OAI22_X1 U2335 ( .A1(n12284), .A2(n12534), .B1(n9955), .B2(n1133), .ZN(n3118) );
  OAI22_X1 U2336 ( .A1(n12284), .A2(n12531), .B1(n9956), .B2(n1133), .ZN(n3119) );
  OAI22_X1 U2337 ( .A1(n12284), .A2(n12528), .B1(n9957), .B2(n1133), .ZN(n3120) );
  OAI22_X1 U2338 ( .A1(n12284), .A2(n12525), .B1(n9958), .B2(n1133), .ZN(n3121) );
  OAI22_X1 U2339 ( .A1(n12283), .A2(n12522), .B1(n9959), .B2(n1133), .ZN(n3122) );
  OAI22_X1 U2340 ( .A1(n12321), .A2(n12552), .B1(n9960), .B2(n12314), .ZN(
        n3243) );
  OAI22_X1 U2341 ( .A1(n12321), .A2(n12540), .B1(n9961), .B2(n12314), .ZN(
        n3244) );
  OAI22_X1 U2342 ( .A1(n12320), .A2(n12537), .B1(n9962), .B2(n1129), .ZN(n3245) );
  OAI22_X1 U2343 ( .A1(n12320), .A2(n12534), .B1(n9963), .B2(n1129), .ZN(n3246) );
  OAI22_X1 U2344 ( .A1(n12320), .A2(n12531), .B1(n9964), .B2(n1129), .ZN(n3247) );
  OAI22_X1 U2345 ( .A1(n12320), .A2(n12528), .B1(n9965), .B2(n1129), .ZN(n3248) );
  OAI22_X1 U2346 ( .A1(n12320), .A2(n12525), .B1(n9966), .B2(n1129), .ZN(n3249) );
  OAI22_X1 U2347 ( .A1(n12319), .A2(n12522), .B1(n9967), .B2(n1129), .ZN(n3250) );
  OAI22_X1 U2348 ( .A1(n12366), .A2(n12552), .B1(n9968), .B2(n12359), .ZN(
        n3467) );
  OAI22_X1 U2349 ( .A1(n12366), .A2(n12540), .B1(n9969), .B2(n12359), .ZN(
        n3468) );
  OAI22_X1 U2350 ( .A1(n12365), .A2(n12537), .B1(n9970), .B2(n1123), .ZN(n3469) );
  OAI22_X1 U2351 ( .A1(n12365), .A2(n12534), .B1(n9971), .B2(n1123), .ZN(n3470) );
  OAI22_X1 U2352 ( .A1(n12365), .A2(n12531), .B1(n9972), .B2(n1123), .ZN(n3471) );
  OAI22_X1 U2353 ( .A1(n12365), .A2(n12528), .B1(n9973), .B2(n1123), .ZN(n3472) );
  OAI22_X1 U2354 ( .A1(n12365), .A2(n12525), .B1(n9974), .B2(n1123), .ZN(n3473) );
  OAI22_X1 U2355 ( .A1(n12364), .A2(n12522), .B1(n9975), .B2(n1123), .ZN(n3474) );
  OAI22_X1 U2356 ( .A1(n12384), .A2(n12553), .B1(n9976), .B2(n12377), .ZN(
        n3595) );
  OAI22_X1 U2357 ( .A1(n12384), .A2(n12541), .B1(n9977), .B2(n12377), .ZN(
        n3596) );
  OAI22_X1 U2358 ( .A1(n12383), .A2(n12538), .B1(n9978), .B2(n1121), .ZN(n3597) );
  OAI22_X1 U2359 ( .A1(n12383), .A2(n12535), .B1(n9979), .B2(n1121), .ZN(n3598) );
  OAI22_X1 U2360 ( .A1(n12383), .A2(n12532), .B1(n9980), .B2(n1121), .ZN(n3599) );
  OAI22_X1 U2361 ( .A1(n12383), .A2(n12529), .B1(n9981), .B2(n1121), .ZN(n3600) );
  OAI22_X1 U2362 ( .A1(n12383), .A2(n12526), .B1(n9982), .B2(n1121), .ZN(n3601) );
  OAI22_X1 U2363 ( .A1(n12382), .A2(n12523), .B1(n9983), .B2(n1121), .ZN(n3602) );
  OAI22_X1 U2364 ( .A1(n12173), .A2(n12479), .B1(n9985), .B2(n1146), .ZN(n2624) );
  OAI22_X1 U2365 ( .A1(n12191), .A2(n12479), .B1(n9990), .B2(n1144), .ZN(n2752) );
  OAI22_X1 U2366 ( .A1(n12209), .A2(n12479), .B1(n9995), .B2(n12206), .ZN(
        n2880) );
  OAI22_X1 U2367 ( .A1(n12181), .A2(n12476), .B1(n12179), .B2(n11704), .ZN(
        n2657) );
  OAI22_X1 U2368 ( .A1(n12181), .A2(n12473), .B1(n12179), .B2(n11705), .ZN(
        n2658) );
  OAI22_X1 U2369 ( .A1(n12181), .A2(n12470), .B1(n12179), .B2(n11706), .ZN(
        n2659) );
  OAI22_X1 U2370 ( .A1(n12181), .A2(n12467), .B1(n12179), .B2(n11707), .ZN(
        n2660) );
  OAI22_X1 U2371 ( .A1(n12181), .A2(n12464), .B1(n1145), .B2(n11708), .ZN(
        n2661) );
  OAI22_X1 U2372 ( .A1(n12180), .A2(n12461), .B1(n1145), .B2(n11709), .ZN(
        n2662) );
  OAI22_X1 U2373 ( .A1(n12180), .A2(n12458), .B1(n1145), .B2(n11710), .ZN(
        n2663) );
  OAI22_X1 U2374 ( .A1(n12180), .A2(n12455), .B1(n1145), .B2(n11711), .ZN(
        n2664) );
  OAI22_X1 U2375 ( .A1(n12180), .A2(n12452), .B1(n1145), .B2(n11712), .ZN(
        n2665) );
  OAI22_X1 U2376 ( .A1(n12180), .A2(n12449), .B1(n1145), .B2(n11713), .ZN(
        n2666) );
  OAI22_X1 U2377 ( .A1(n12199), .A2(n12476), .B1(n12197), .B2(n11714), .ZN(
        n2785) );
  OAI22_X1 U2378 ( .A1(n12199), .A2(n12473), .B1(n12197), .B2(n11715), .ZN(
        n2786) );
  OAI22_X1 U2379 ( .A1(n12199), .A2(n12470), .B1(n12197), .B2(n11716), .ZN(
        n2787) );
  OAI22_X1 U2380 ( .A1(n12199), .A2(n12467), .B1(n12197), .B2(n11717), .ZN(
        n2788) );
  OAI22_X1 U2381 ( .A1(n12199), .A2(n12464), .B1(n1143), .B2(n11718), .ZN(
        n2789) );
  OAI22_X1 U2382 ( .A1(n12198), .A2(n12461), .B1(n1143), .B2(n11719), .ZN(
        n2790) );
  OAI22_X1 U2383 ( .A1(n12198), .A2(n12458), .B1(n1143), .B2(n11720), .ZN(
        n2791) );
  OAI22_X1 U2384 ( .A1(n12198), .A2(n12455), .B1(n1143), .B2(n11721), .ZN(
        n2792) );
  OAI22_X1 U2385 ( .A1(n12198), .A2(n12452), .B1(n1143), .B2(n11722), .ZN(
        n2793) );
  OAI22_X1 U2386 ( .A1(n12198), .A2(n12449), .B1(n1143), .B2(n11723), .ZN(
        n2794) );
  OAI22_X1 U2387 ( .A1(n12217), .A2(n12476), .B1(n12215), .B2(n11724), .ZN(
        n2913) );
  OAI22_X1 U2388 ( .A1(n12217), .A2(n12473), .B1(n12215), .B2(n11725), .ZN(
        n2914) );
  OAI22_X1 U2389 ( .A1(n12217), .A2(n12470), .B1(n12215), .B2(n11726), .ZN(
        n2915) );
  OAI22_X1 U2390 ( .A1(n12217), .A2(n12467), .B1(n12215), .B2(n11727), .ZN(
        n2916) );
  OAI22_X1 U2391 ( .A1(n12217), .A2(n12464), .B1(n1141), .B2(n11728), .ZN(
        n2917) );
  OAI22_X1 U2392 ( .A1(n12216), .A2(n12461), .B1(n1141), .B2(n11729), .ZN(
        n2918) );
  OAI22_X1 U2393 ( .A1(n12216), .A2(n12458), .B1(n1141), .B2(n11730), .ZN(
        n2919) );
  OAI22_X1 U2394 ( .A1(n12216), .A2(n12455), .B1(n1141), .B2(n11731), .ZN(
        n2920) );
  OAI22_X1 U2395 ( .A1(n12216), .A2(n12452), .B1(n1141), .B2(n11732), .ZN(
        n2921) );
  OAI22_X1 U2396 ( .A1(n12216), .A2(n12449), .B1(n1141), .B2(n11733), .ZN(
        n2922) );
  OAI22_X1 U2397 ( .A1(n12253), .A2(n12476), .B1(n12251), .B2(n11734), .ZN(
        n3041) );
  OAI22_X1 U2398 ( .A1(n12253), .A2(n12473), .B1(n12251), .B2(n11735), .ZN(
        n3042) );
  OAI22_X1 U2399 ( .A1(n12253), .A2(n12470), .B1(n12251), .B2(n11736), .ZN(
        n3043) );
  OAI22_X1 U2400 ( .A1(n12253), .A2(n12467), .B1(n12251), .B2(n11737), .ZN(
        n3044) );
  OAI22_X1 U2401 ( .A1(n12253), .A2(n12464), .B1(n1137), .B2(n11738), .ZN(
        n3045) );
  OAI22_X1 U2402 ( .A1(n12252), .A2(n12461), .B1(n1137), .B2(n11739), .ZN(
        n3046) );
  OAI22_X1 U2403 ( .A1(n12252), .A2(n12458), .B1(n1137), .B2(n11740), .ZN(
        n3047) );
  OAI22_X1 U2404 ( .A1(n12252), .A2(n12455), .B1(n1137), .B2(n11741), .ZN(
        n3048) );
  OAI22_X1 U2405 ( .A1(n12252), .A2(n12452), .B1(n1137), .B2(n11742), .ZN(
        n3049) );
  OAI22_X1 U2406 ( .A1(n12252), .A2(n12449), .B1(n1137), .B2(n11743), .ZN(
        n3050) );
  OAI22_X1 U2407 ( .A1(n12289), .A2(n12477), .B1(n12287), .B2(n11744), .ZN(
        n3169) );
  OAI22_X1 U2408 ( .A1(n12289), .A2(n12474), .B1(n12287), .B2(n11745), .ZN(
        n3170) );
  OAI22_X1 U2409 ( .A1(n12289), .A2(n12471), .B1(n12287), .B2(n11746), .ZN(
        n3171) );
  OAI22_X1 U2410 ( .A1(n12289), .A2(n12468), .B1(n12287), .B2(n11747), .ZN(
        n3172) );
  OAI22_X1 U2411 ( .A1(n12289), .A2(n12465), .B1(n1132), .B2(n11748), .ZN(
        n3173) );
  OAI22_X1 U2412 ( .A1(n12288), .A2(n12462), .B1(n1132), .B2(n11749), .ZN(
        n3174) );
  OAI22_X1 U2413 ( .A1(n12288), .A2(n12459), .B1(n1132), .B2(n11750), .ZN(
        n3175) );
  OAI22_X1 U2414 ( .A1(n12288), .A2(n12456), .B1(n1132), .B2(n11751), .ZN(
        n3176) );
  OAI22_X1 U2415 ( .A1(n12288), .A2(n12453), .B1(n1132), .B2(n11752), .ZN(
        n3177) );
  OAI22_X1 U2416 ( .A1(n12288), .A2(n12450), .B1(n1132), .B2(n11753), .ZN(
        n3178) );
  OAI22_X1 U2417 ( .A1(n12325), .A2(n12477), .B1(n12323), .B2(n11754), .ZN(
        n3297) );
  OAI22_X1 U2418 ( .A1(n12325), .A2(n12474), .B1(n12323), .B2(n11755), .ZN(
        n3298) );
  OAI22_X1 U2419 ( .A1(n12325), .A2(n12471), .B1(n12323), .B2(n11756), .ZN(
        n3299) );
  OAI22_X1 U2420 ( .A1(n12325), .A2(n12468), .B1(n12323), .B2(n11757), .ZN(
        n3300) );
  OAI22_X1 U2421 ( .A1(n12325), .A2(n12465), .B1(n1128), .B2(n11758), .ZN(
        n3301) );
  OAI22_X1 U2422 ( .A1(n12324), .A2(n12462), .B1(n1128), .B2(n11759), .ZN(
        n3302) );
  OAI22_X1 U2423 ( .A1(n12324), .A2(n12459), .B1(n1128), .B2(n11760), .ZN(
        n3303) );
  OAI22_X1 U2424 ( .A1(n12324), .A2(n12456), .B1(n1128), .B2(n11761), .ZN(
        n3304) );
  OAI22_X1 U2425 ( .A1(n12324), .A2(n12453), .B1(n1128), .B2(n11762), .ZN(
        n3305) );
  OAI22_X1 U2426 ( .A1(n12324), .A2(n12450), .B1(n1128), .B2(n11763), .ZN(
        n3306) );
  OAI22_X1 U2427 ( .A1(n12352), .A2(n12477), .B1(n12350), .B2(n11764), .ZN(
        n3457) );
  OAI22_X1 U2428 ( .A1(n12352), .A2(n12474), .B1(n12350), .B2(n11765), .ZN(
        n3458) );
  OAI22_X1 U2429 ( .A1(n12352), .A2(n12471), .B1(n12350), .B2(n11766), .ZN(
        n3459) );
  OAI22_X1 U2430 ( .A1(n12352), .A2(n12468), .B1(n12350), .B2(n11767), .ZN(
        n3460) );
  OAI22_X1 U2431 ( .A1(n12352), .A2(n12465), .B1(n1124), .B2(n11768), .ZN(
        n3461) );
  OAI22_X1 U2432 ( .A1(n12351), .A2(n12462), .B1(n1124), .B2(n11769), .ZN(
        n3462) );
  OAI22_X1 U2433 ( .A1(n12351), .A2(n12459), .B1(n1124), .B2(n11770), .ZN(
        n3463) );
  OAI22_X1 U2434 ( .A1(n12351), .A2(n12456), .B1(n1124), .B2(n11771), .ZN(
        n3464) );
  OAI22_X1 U2435 ( .A1(n12351), .A2(n12453), .B1(n1124), .B2(n11772), .ZN(
        n3465) );
  OAI22_X1 U2436 ( .A1(n12351), .A2(n12450), .B1(n1124), .B2(n11773), .ZN(
        n3466) );
  OAI22_X1 U2437 ( .A1(n12370), .A2(n12478), .B1(n12368), .B2(n11774), .ZN(
        n3585) );
  OAI22_X1 U2438 ( .A1(n12370), .A2(n12475), .B1(n12368), .B2(n11775), .ZN(
        n3586) );
  OAI22_X1 U2439 ( .A1(n12370), .A2(n12472), .B1(n12368), .B2(n11776), .ZN(
        n3587) );
  OAI22_X1 U2440 ( .A1(n12370), .A2(n12469), .B1(n12368), .B2(n11777), .ZN(
        n3588) );
  OAI22_X1 U2441 ( .A1(n12370), .A2(n12466), .B1(n1122), .B2(n11778), .ZN(
        n3589) );
  OAI22_X1 U2442 ( .A1(n12369), .A2(n12463), .B1(n1122), .B2(n11779), .ZN(
        n3590) );
  OAI22_X1 U2443 ( .A1(n12369), .A2(n12460), .B1(n1122), .B2(n11780), .ZN(
        n3591) );
  OAI22_X1 U2444 ( .A1(n12369), .A2(n12457), .B1(n1122), .B2(n11781), .ZN(
        n3592) );
  OAI22_X1 U2445 ( .A1(n12369), .A2(n12454), .B1(n1122), .B2(n11782), .ZN(
        n3593) );
  OAI22_X1 U2446 ( .A1(n12369), .A2(n12451), .B1(n1122), .B2(n11783), .ZN(
        n3594) );
  INV_X1 U2447 ( .A(ADD_WR[4]), .ZN(n12566) );
  INV_X1 U2448 ( .A(ADD_WR[3]), .ZN(n12560) );
  NAND4_X1 U2449 ( .A1(n2467), .A2(n2468), .A3(n2469), .A4(n2470), .ZN(n2437)
         );
  XNOR2_X1 U2450 ( .A(ADD_RD2[1]), .B(ADD_WR[1]), .ZN(n2467) );
  XNOR2_X1 U2451 ( .A(ADD_RD2[2]), .B(ADD_WR[2]), .ZN(n2469) );
  XNOR2_X1 U2452 ( .A(ADD_WR[3]), .B(ADD_RD2[3]), .ZN(n2468) );
  NAND2_X1 U2453 ( .A1(DATAIN[25]), .A2(n12554), .ZN(n1097) );
  NAND2_X1 U2454 ( .A1(DATAIN[26]), .A2(n12554), .ZN(n1098) );
  NAND2_X1 U2455 ( .A1(DATAIN[29]), .A2(n12554), .ZN(n1101) );
  NAND2_X1 U2456 ( .A1(DATAIN[30]), .A2(n12554), .ZN(n1102) );
  NAND2_X1 U2457 ( .A1(DATAIN[23]), .A2(n12554), .ZN(n1095) );
  NOR2_X1 U2458 ( .A1(n12573), .A2(ADD_RD1[2]), .ZN(n1786) );
  NOR3_X1 U2459 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n12572), .ZN(n1796) );
  NOR3_X1 U2460 ( .A1(n12571), .A2(ADD_RD1[4]), .A3(n12572), .ZN(n1797) );
  NOR3_X1 U2461 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(n1801) );
  NOR3_X1 U2462 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n12571), .ZN(n1800) );
  AOI221_X1 U2463 ( .B1(n12110), .B2(n8389), .C1(n12107), .C2(n7933), .A(n1615), .ZN(n1614) );
  OAI22_X1 U2464 ( .A1(n10936), .A2(n12104), .B1(n11192), .B2(n12101), .ZN(
        n1615) );
  AOI221_X1 U2465 ( .B1(n12110), .B2(n8391), .C1(n12107), .C2(n7935), .A(n1596), .ZN(n1595) );
  OAI22_X1 U2466 ( .A1(n10937), .A2(n12104), .B1(n11193), .B2(n12101), .ZN(
        n1596) );
  AOI221_X1 U2467 ( .B1(n12111), .B2(n8393), .C1(n12108), .C2(n7937), .A(n1577), .ZN(n1576) );
  OAI22_X1 U2468 ( .A1(n10938), .A2(n12104), .B1(n11194), .B2(n12101), .ZN(
        n1577) );
  AOI221_X1 U2469 ( .B1(n12111), .B2(n8395), .C1(n12108), .C2(n7939), .A(n1558), .ZN(n1557) );
  OAI22_X1 U2470 ( .A1(n10939), .A2(n12105), .B1(n11195), .B2(n12102), .ZN(
        n1558) );
  AOI221_X1 U2471 ( .B1(n12111), .B2(n8397), .C1(n12108), .C2(n7941), .A(n1539), .ZN(n1538) );
  OAI22_X1 U2472 ( .A1(n10940), .A2(n12105), .B1(n11196), .B2(n12102), .ZN(
        n1539) );
  AOI221_X1 U2473 ( .B1(n12111), .B2(n8399), .C1(n12108), .C2(n7943), .A(n1520), .ZN(n1519) );
  OAI22_X1 U2474 ( .A1(n10941), .A2(n12105), .B1(n11197), .B2(n12102), .ZN(
        n1520) );
  AOI221_X1 U2475 ( .B1(n12111), .B2(n8401), .C1(n12108), .C2(n7945), .A(n1501), .ZN(n1500) );
  OAI22_X1 U2476 ( .A1(n10942), .A2(n12105), .B1(n11198), .B2(n12102), .ZN(
        n1501) );
  AOI221_X1 U2477 ( .B1(n12111), .B2(n8403), .C1(n12108), .C2(n7947), .A(n1482), .ZN(n1481) );
  OAI22_X1 U2478 ( .A1(n10943), .A2(n12105), .B1(n11199), .B2(n12102), .ZN(
        n1482) );
  AOI221_X1 U2479 ( .B1(n12111), .B2(n8405), .C1(n12108), .C2(n7949), .A(n1463), .ZN(n1462) );
  OAI22_X1 U2480 ( .A1(n10944), .A2(n12105), .B1(n11200), .B2(n12102), .ZN(
        n1463) );
  AOI221_X1 U2481 ( .B1(n12111), .B2(n8407), .C1(n12108), .C2(n7951), .A(n1444), .ZN(n1443) );
  OAI22_X1 U2482 ( .A1(n10945), .A2(n12105), .B1(n11201), .B2(n12102), .ZN(
        n1444) );
  AOI221_X1 U2483 ( .B1(n12111), .B2(n8409), .C1(n12108), .C2(n7953), .A(n1425), .ZN(n1424) );
  OAI22_X1 U2484 ( .A1(n10946), .A2(n12105), .B1(n11202), .B2(n12102), .ZN(
        n1425) );
  AOI221_X1 U2485 ( .B1(n12111), .B2(n8411), .C1(n12108), .C2(n7955), .A(n1406), .ZN(n1405) );
  OAI22_X1 U2486 ( .A1(n10947), .A2(n12105), .B1(n11203), .B2(n12102), .ZN(
        n1406) );
  AOI221_X1 U2487 ( .B1(n12111), .B2(n8413), .C1(n12108), .C2(n7957), .A(n1387), .ZN(n1386) );
  OAI22_X1 U2488 ( .A1(n10948), .A2(n12105), .B1(n11204), .B2(n12102), .ZN(
        n1387) );
  AOI221_X1 U2489 ( .B1(n12112), .B2(n8415), .C1(n12109), .C2(n7959), .A(n1368), .ZN(n1367) );
  OAI22_X1 U2490 ( .A1(n10949), .A2(n12105), .B1(n11205), .B2(n12102), .ZN(
        n1368) );
  AOI221_X1 U2491 ( .B1(n12112), .B2(n8417), .C1(n12109), .C2(n7961), .A(n1349), .ZN(n1348) );
  OAI22_X1 U2492 ( .A1(n10950), .A2(n12105), .B1(n11206), .B2(n12102), .ZN(
        n1349) );
  AOI221_X1 U2493 ( .B1(n12110), .B2(n11448), .C1(n12107), .C2(n7915), .A(
        n1795), .ZN(n1794) );
  OAI22_X1 U2494 ( .A1(n10951), .A2(n12104), .B1(n11207), .B2(n12101), .ZN(
        n1795) );
  AOI221_X1 U2495 ( .B1(n12110), .B2(n11449), .C1(n12107), .C2(n7917), .A(
        n1767), .ZN(n1766) );
  OAI22_X1 U2496 ( .A1(n10952), .A2(n12104), .B1(n11208), .B2(n12101), .ZN(
        n1767) );
  AOI221_X1 U2497 ( .B1(n12110), .B2(n11450), .C1(n12107), .C2(n7919), .A(
        n1748), .ZN(n1747) );
  OAI22_X1 U2498 ( .A1(n10953), .A2(n12104), .B1(n11209), .B2(n12101), .ZN(
        n1748) );
  AOI221_X1 U2499 ( .B1(n12110), .B2(n11451), .C1(n12107), .C2(n7921), .A(
        n1729), .ZN(n1728) );
  OAI22_X1 U2500 ( .A1(n10954), .A2(n12104), .B1(n11210), .B2(n12101), .ZN(
        n1729) );
  AOI221_X1 U2501 ( .B1(n12110), .B2(n11452), .C1(n12107), .C2(n7923), .A(
        n1710), .ZN(n1709) );
  OAI22_X1 U2502 ( .A1(n10955), .A2(n12104), .B1(n11211), .B2(n12101), .ZN(
        n1710) );
  AOI221_X1 U2503 ( .B1(n12110), .B2(n11453), .C1(n12107), .C2(n7925), .A(
        n1691), .ZN(n1690) );
  OAI22_X1 U2504 ( .A1(n10956), .A2(n12104), .B1(n11212), .B2(n12101), .ZN(
        n1691) );
  AOI221_X1 U2505 ( .B1(n12110), .B2(n11454), .C1(n12107), .C2(n7927), .A(
        n1672), .ZN(n1671) );
  OAI22_X1 U2506 ( .A1(n10957), .A2(n12104), .B1(n11213), .B2(n12101), .ZN(
        n1672) );
  AOI221_X1 U2507 ( .B1(n12110), .B2(n11455), .C1(n12107), .C2(n7929), .A(
        n1653), .ZN(n1652) );
  OAI22_X1 U2508 ( .A1(n10958), .A2(n12104), .B1(n11214), .B2(n12101), .ZN(
        n1653) );
  AOI221_X1 U2509 ( .B1(n12146), .B2(n8436), .C1(n12143), .C2(n7980), .A(n1627), .ZN(n1624) );
  OAI22_X1 U2510 ( .A1(n10959), .A2(n12140), .B1(n11215), .B2(n12137), .ZN(
        n1627) );
  AOI221_X1 U2511 ( .B1(n12098), .B2(n8437), .C1(n12095), .C2(n7981), .A(n1635), .ZN(n1632) );
  OAI22_X1 U2512 ( .A1(n10960), .A2(n12092), .B1(n11216), .B2(n12089), .ZN(
        n1635) );
  AOI221_X1 U2513 ( .B1(n12098), .B2(n8439), .C1(n12095), .C2(n7983), .A(n1616), .ZN(n1613) );
  OAI22_X1 U2514 ( .A1(n10961), .A2(n12092), .B1(n11217), .B2(n12089), .ZN(
        n1616) );
  AOI221_X1 U2515 ( .B1(n12098), .B2(n8441), .C1(n12095), .C2(n7985), .A(n1597), .ZN(n1594) );
  OAI22_X1 U2516 ( .A1(n10962), .A2(n12092), .B1(n11218), .B2(n12089), .ZN(
        n1597) );
  AOI221_X1 U2517 ( .B1(n12099), .B2(n8443), .C1(n12096), .C2(n7987), .A(n1578), .ZN(n1575) );
  OAI22_X1 U2518 ( .A1(n10963), .A2(n12092), .B1(n11219), .B2(n12089), .ZN(
        n1578) );
  AOI221_X1 U2519 ( .B1(n12099), .B2(n8445), .C1(n12096), .C2(n7989), .A(n1559), .ZN(n1556) );
  OAI22_X1 U2520 ( .A1(n10964), .A2(n12093), .B1(n11220), .B2(n12090), .ZN(
        n1559) );
  AOI221_X1 U2521 ( .B1(n12099), .B2(n8447), .C1(n12096), .C2(n7991), .A(n1540), .ZN(n1537) );
  OAI22_X1 U2522 ( .A1(n10965), .A2(n12093), .B1(n11221), .B2(n12090), .ZN(
        n1540) );
  AOI221_X1 U2523 ( .B1(n12099), .B2(n8449), .C1(n12096), .C2(n7993), .A(n1521), .ZN(n1518) );
  OAI22_X1 U2524 ( .A1(n10966), .A2(n12093), .B1(n11222), .B2(n12090), .ZN(
        n1521) );
  AOI221_X1 U2525 ( .B1(n12099), .B2(n8451), .C1(n12096), .C2(n7995), .A(n1502), .ZN(n1499) );
  OAI22_X1 U2526 ( .A1(n10967), .A2(n12093), .B1(n11223), .B2(n12090), .ZN(
        n1502) );
  AOI221_X1 U2527 ( .B1(n12099), .B2(n8453), .C1(n12096), .C2(n7997), .A(n1483), .ZN(n1480) );
  OAI22_X1 U2528 ( .A1(n10968), .A2(n12093), .B1(n11224), .B2(n12090), .ZN(
        n1483) );
  AOI221_X1 U2529 ( .B1(n12099), .B2(n8455), .C1(n12096), .C2(n7999), .A(n1464), .ZN(n1461) );
  OAI22_X1 U2530 ( .A1(n10969), .A2(n12093), .B1(n11225), .B2(n12090), .ZN(
        n1464) );
  AOI221_X1 U2531 ( .B1(n12099), .B2(n8457), .C1(n12096), .C2(n8001), .A(n1445), .ZN(n1442) );
  OAI22_X1 U2532 ( .A1(n10970), .A2(n12093), .B1(n11226), .B2(n12090), .ZN(
        n1445) );
  AOI221_X1 U2533 ( .B1(n12099), .B2(n8459), .C1(n12096), .C2(n8003), .A(n1426), .ZN(n1423) );
  OAI22_X1 U2534 ( .A1(n10971), .A2(n12093), .B1(n11227), .B2(n12090), .ZN(
        n1426) );
  AOI221_X1 U2535 ( .B1(n12099), .B2(n8461), .C1(n12096), .C2(n8005), .A(n1407), .ZN(n1404) );
  OAI22_X1 U2536 ( .A1(n10972), .A2(n12093), .B1(n11228), .B2(n12090), .ZN(
        n1407) );
  AOI221_X1 U2537 ( .B1(n12099), .B2(n8463), .C1(n12096), .C2(n8007), .A(n1388), .ZN(n1385) );
  OAI22_X1 U2538 ( .A1(n10973), .A2(n12093), .B1(n11229), .B2(n12090), .ZN(
        n1388) );
  AOI221_X1 U2539 ( .B1(n12100), .B2(n8465), .C1(n12097), .C2(n8009), .A(n1369), .ZN(n1366) );
  OAI22_X1 U2540 ( .A1(n10974), .A2(n12093), .B1(n11230), .B2(n12090), .ZN(
        n1369) );
  AOI221_X1 U2541 ( .B1(n12100), .B2(n8467), .C1(n12097), .C2(n8011), .A(n1350), .ZN(n1347) );
  OAI22_X1 U2542 ( .A1(n10975), .A2(n12093), .B1(n11231), .B2(n12090), .ZN(
        n1350) );
  AOI221_X1 U2543 ( .B1(n12148), .B2(n9573), .C1(n12145), .C2(n9885), .A(n1304), .ZN(n1301) );
  OAI22_X1 U2544 ( .A1(n10976), .A2(n12142), .B1(n11232), .B2(n12139), .ZN(
        n1304) );
  AOI221_X1 U2545 ( .B1(n12148), .B2(n9574), .C1(n12145), .C2(n9886), .A(n1285), .ZN(n1282) );
  OAI22_X1 U2546 ( .A1(n10977), .A2(n12142), .B1(n11233), .B2(n12139), .ZN(
        n1285) );
  AOI221_X1 U2547 ( .B1(n12148), .B2(n9575), .C1(n12145), .C2(n9887), .A(n1266), .ZN(n1263) );
  OAI22_X1 U2548 ( .A1(n10978), .A2(n12142), .B1(n11234), .B2(n12139), .ZN(
        n1266) );
  AOI221_X1 U2549 ( .B1(n12148), .B2(n9576), .C1(n12145), .C2(n9888), .A(n1247), .ZN(n1244) );
  OAI22_X1 U2550 ( .A1(n10979), .A2(n12142), .B1(n11235), .B2(n12139), .ZN(
        n1247) );
  AOI221_X1 U2551 ( .B1(n12148), .B2(n9577), .C1(n12145), .C2(n9889), .A(n1228), .ZN(n1225) );
  OAI22_X1 U2552 ( .A1(n10980), .A2(n12142), .B1(n11236), .B2(n12139), .ZN(
        n1228) );
  AOI221_X1 U2553 ( .B1(n12148), .B2(n9578), .C1(n12145), .C2(n9890), .A(n1209), .ZN(n1206) );
  OAI22_X1 U2554 ( .A1(n10981), .A2(n12142), .B1(n11237), .B2(n12139), .ZN(
        n1209) );
  AOI221_X1 U2555 ( .B1(n12148), .B2(n9579), .C1(n12145), .C2(n9891), .A(n1164), .ZN(n1155) );
  OAI22_X1 U2556 ( .A1(n10982), .A2(n12142), .B1(n11238), .B2(n12139), .ZN(
        n1164) );
  AOI221_X1 U2557 ( .B1(n12098), .B2(n11456), .C1(n12095), .C2(n7965), .A(
        n1798), .ZN(n1793) );
  OAI22_X1 U2558 ( .A1(n10983), .A2(n12092), .B1(n11239), .B2(n12089), .ZN(
        n1798) );
  AOI221_X1 U2559 ( .B1(n12098), .B2(n11457), .C1(n12095), .C2(n7967), .A(
        n1768), .ZN(n1765) );
  OAI22_X1 U2560 ( .A1(n10984), .A2(n12092), .B1(n11240), .B2(n12089), .ZN(
        n1768) );
  AOI221_X1 U2561 ( .B1(n12098), .B2(n11458), .C1(n12095), .C2(n7969), .A(
        n1749), .ZN(n1746) );
  OAI22_X1 U2562 ( .A1(n10985), .A2(n12092), .B1(n11241), .B2(n12089), .ZN(
        n1749) );
  AOI221_X1 U2563 ( .B1(n12098), .B2(n11459), .C1(n12095), .C2(n7971), .A(
        n1730), .ZN(n1727) );
  OAI22_X1 U2564 ( .A1(n10986), .A2(n12092), .B1(n11242), .B2(n12089), .ZN(
        n1730) );
  AOI221_X1 U2565 ( .B1(n12098), .B2(n11460), .C1(n12095), .C2(n7973), .A(
        n1711), .ZN(n1708) );
  OAI22_X1 U2566 ( .A1(n10987), .A2(n12092), .B1(n11243), .B2(n12089), .ZN(
        n1711) );
  AOI221_X1 U2567 ( .B1(n12098), .B2(n11461), .C1(n12095), .C2(n7975), .A(
        n1692), .ZN(n1689) );
  OAI22_X1 U2568 ( .A1(n10988), .A2(n12092), .B1(n11244), .B2(n12089), .ZN(
        n1692) );
  AOI221_X1 U2569 ( .B1(n12098), .B2(n11462), .C1(n12095), .C2(n7977), .A(
        n1673), .ZN(n1670) );
  OAI22_X1 U2570 ( .A1(n10989), .A2(n12092), .B1(n11245), .B2(n12089), .ZN(
        n1673) );
  AOI221_X1 U2571 ( .B1(n12098), .B2(n11463), .C1(n12095), .C2(n7979), .A(
        n1654), .ZN(n1651) );
  OAI22_X1 U2572 ( .A1(n10990), .A2(n12092), .B1(n11246), .B2(n12089), .ZN(
        n1654) );
  AOI221_X1 U2573 ( .B1(n12147), .B2(n11464), .C1(n12144), .C2(n8004), .A(
        n1399), .ZN(n1396) );
  OAI22_X1 U2574 ( .A1(n10991), .A2(n12141), .B1(n11247), .B2(n12138), .ZN(
        n1399) );
  AOI221_X1 U2575 ( .B1(n12147), .B2(n11465), .C1(n12144), .C2(n8006), .A(
        n1380), .ZN(n1377) );
  OAI22_X1 U2576 ( .A1(n10992), .A2(n12141), .B1(n11248), .B2(n12138), .ZN(
        n1380) );
  AOI221_X1 U2577 ( .B1(n12148), .B2(n11466), .C1(n12145), .C2(n8008), .A(
        n1361), .ZN(n1358) );
  OAI22_X1 U2578 ( .A1(n10993), .A2(n12141), .B1(n11249), .B2(n12138), .ZN(
        n1361) );
  AOI221_X1 U2579 ( .B1(n12148), .B2(n11467), .C1(n12145), .C2(n8010), .A(
        n1342), .ZN(n1339) );
  OAI22_X1 U2580 ( .A1(n10994), .A2(n12141), .B1(n11250), .B2(n12138), .ZN(
        n1342) );
  AOI221_X1 U2581 ( .B1(n12148), .B2(n11468), .C1(n12145), .C2(n8012), .A(
        n1323), .ZN(n1320) );
  OAI22_X1 U2582 ( .A1(n10995), .A2(n12142), .B1(n11251), .B2(n12139), .ZN(
        n1323) );
  AOI221_X1 U2583 ( .B1(n12134), .B2(n8538), .C1(n12131), .C2(n8082), .A(n1628), .ZN(n1623) );
  OAI22_X1 U2584 ( .A1(n10996), .A2(n12128), .B1(n11252), .B2(n12125), .ZN(
        n1628) );
  AOI221_X1 U2585 ( .B1(n12086), .B2(n8478), .C1(n12083), .C2(n8022), .A(n1636), .ZN(n1631) );
  OAI22_X1 U2586 ( .A1(n10997), .A2(n12080), .B1(n11253), .B2(n12077), .ZN(
        n1636) );
  AOI221_X1 U2587 ( .B1(n12086), .B2(n8479), .C1(n12083), .C2(n8023), .A(n1617), .ZN(n1612) );
  OAI22_X1 U2588 ( .A1(n10998), .A2(n12080), .B1(n11254), .B2(n12077), .ZN(
        n1617) );
  AOI221_X1 U2589 ( .B1(n12086), .B2(n8480), .C1(n12083), .C2(n8024), .A(n1598), .ZN(n1593) );
  OAI22_X1 U2590 ( .A1(n10999), .A2(n12080), .B1(n11255), .B2(n12077), .ZN(
        n1598) );
  AOI221_X1 U2591 ( .B1(n12087), .B2(n8481), .C1(n12084), .C2(n8025), .A(n1579), .ZN(n1574) );
  OAI22_X1 U2592 ( .A1(n11000), .A2(n12080), .B1(n11256), .B2(n12077), .ZN(
        n1579) );
  AOI221_X1 U2593 ( .B1(n12087), .B2(n8482), .C1(n12084), .C2(n8026), .A(n1560), .ZN(n1555) );
  OAI22_X1 U2594 ( .A1(n11001), .A2(n12081), .B1(n11257), .B2(n12078), .ZN(
        n1560) );
  AOI221_X1 U2595 ( .B1(n12087), .B2(n8483), .C1(n12084), .C2(n8027), .A(n1541), .ZN(n1536) );
  OAI22_X1 U2596 ( .A1(n11002), .A2(n12081), .B1(n11258), .B2(n12078), .ZN(
        n1541) );
  AOI221_X1 U2597 ( .B1(n12087), .B2(n8484), .C1(n12084), .C2(n8028), .A(n1522), .ZN(n1517) );
  OAI22_X1 U2598 ( .A1(n11003), .A2(n12081), .B1(n11259), .B2(n12078), .ZN(
        n1522) );
  AOI221_X1 U2599 ( .B1(n12087), .B2(n8485), .C1(n12084), .C2(n8029), .A(n1503), .ZN(n1498) );
  OAI22_X1 U2600 ( .A1(n11004), .A2(n12081), .B1(n11260), .B2(n12078), .ZN(
        n1503) );
  AOI221_X1 U2601 ( .B1(n12087), .B2(n8486), .C1(n12084), .C2(n8030), .A(n1484), .ZN(n1479) );
  OAI22_X1 U2602 ( .A1(n11005), .A2(n12081), .B1(n11261), .B2(n12078), .ZN(
        n1484) );
  AOI221_X1 U2603 ( .B1(n12087), .B2(n8487), .C1(n12084), .C2(n8031), .A(n1465), .ZN(n1460) );
  OAI22_X1 U2604 ( .A1(n11006), .A2(n12081), .B1(n11262), .B2(n12078), .ZN(
        n1465) );
  AOI221_X1 U2605 ( .B1(n12087), .B2(n8488), .C1(n12084), .C2(n8032), .A(n1446), .ZN(n1441) );
  OAI22_X1 U2606 ( .A1(n11007), .A2(n12081), .B1(n11263), .B2(n12078), .ZN(
        n1446) );
  AOI221_X1 U2607 ( .B1(n12087), .B2(n8489), .C1(n12084), .C2(n8033), .A(n1427), .ZN(n1422) );
  OAI22_X1 U2608 ( .A1(n11008), .A2(n12081), .B1(n11264), .B2(n12078), .ZN(
        n1427) );
  AOI221_X1 U2609 ( .B1(n12087), .B2(n8490), .C1(n12084), .C2(n8034), .A(n1408), .ZN(n1403) );
  OAI22_X1 U2610 ( .A1(n11009), .A2(n12081), .B1(n11265), .B2(n12078), .ZN(
        n1408) );
  AOI221_X1 U2611 ( .B1(n12087), .B2(n8491), .C1(n12084), .C2(n8035), .A(n1389), .ZN(n1384) );
  OAI22_X1 U2612 ( .A1(n11010), .A2(n12081), .B1(n11266), .B2(n12078), .ZN(
        n1389) );
  AOI221_X1 U2613 ( .B1(n12088), .B2(n8492), .C1(n12085), .C2(n8036), .A(n1370), .ZN(n1365) );
  OAI22_X1 U2614 ( .A1(n11011), .A2(n12081), .B1(n11267), .B2(n12078), .ZN(
        n1370) );
  AOI221_X1 U2615 ( .B1(n12088), .B2(n8493), .C1(n12085), .C2(n8037), .A(n1351), .ZN(n1346) );
  OAI22_X1 U2616 ( .A1(n11012), .A2(n12081), .B1(n11268), .B2(n12078), .ZN(
        n1351) );
  AOI221_X1 U2617 ( .B1(n12136), .B2(n9559), .C1(n12133), .C2(n9871), .A(n1305), .ZN(n1300) );
  OAI22_X1 U2618 ( .A1(n11013), .A2(n12130), .B1(n11269), .B2(n12127), .ZN(
        n1305) );
  AOI221_X1 U2619 ( .B1(n12136), .B2(n9561), .C1(n12133), .C2(n9873), .A(n1286), .ZN(n1281) );
  OAI22_X1 U2620 ( .A1(n11014), .A2(n12130), .B1(n11270), .B2(n12127), .ZN(
        n1286) );
  AOI221_X1 U2621 ( .B1(n12136), .B2(n9563), .C1(n12133), .C2(n9875), .A(n1267), .ZN(n1262) );
  OAI22_X1 U2622 ( .A1(n11015), .A2(n12130), .B1(n11271), .B2(n12127), .ZN(
        n1267) );
  AOI221_X1 U2623 ( .B1(n12136), .B2(n9565), .C1(n12133), .C2(n9877), .A(n1248), .ZN(n1243) );
  OAI22_X1 U2624 ( .A1(n11016), .A2(n12130), .B1(n11272), .B2(n12127), .ZN(
        n1248) );
  AOI221_X1 U2625 ( .B1(n12136), .B2(n9567), .C1(n12133), .C2(n9879), .A(n1229), .ZN(n1224) );
  OAI22_X1 U2626 ( .A1(n11017), .A2(n12130), .B1(n11273), .B2(n12127), .ZN(
        n1229) );
  AOI221_X1 U2627 ( .B1(n12136), .B2(n9569), .C1(n12133), .C2(n9881), .A(n1210), .ZN(n1205) );
  OAI22_X1 U2628 ( .A1(n11018), .A2(n12130), .B1(n11274), .B2(n12127), .ZN(
        n1210) );
  AOI221_X1 U2629 ( .B1(n12136), .B2(n9571), .C1(n12133), .C2(n9883), .A(n1169), .ZN(n1154) );
  OAI22_X1 U2630 ( .A1(n11019), .A2(n12130), .B1(n11275), .B2(n12127), .ZN(
        n1169) );
  AOI221_X1 U2631 ( .B1(n12134), .B2(n11469), .C1(n12131), .C2(n8066), .A(
        n1787), .ZN(n1776) );
  OAI22_X1 U2632 ( .A1(n11020), .A2(n12128), .B1(n11276), .B2(n12125), .ZN(
        n1787) );
  AOI221_X1 U2633 ( .B1(n12086), .B2(n11470), .C1(n12083), .C2(n8014), .A(
        n1799), .ZN(n1792) );
  OAI22_X1 U2634 ( .A1(n11021), .A2(n12080), .B1(n11277), .B2(n12077), .ZN(
        n1799) );
  AOI221_X1 U2635 ( .B1(n12134), .B2(n11471), .C1(n12131), .C2(n8068), .A(
        n1761), .ZN(n1756) );
  OAI22_X1 U2636 ( .A1(n11022), .A2(n12128), .B1(n11278), .B2(n12125), .ZN(
        n1761) );
  AOI221_X1 U2637 ( .B1(n12086), .B2(n11472), .C1(n12083), .C2(n8015), .A(
        n1769), .ZN(n1764) );
  OAI22_X1 U2638 ( .A1(n11023), .A2(n12080), .B1(n11279), .B2(n12077), .ZN(
        n1769) );
  AOI221_X1 U2639 ( .B1(n12134), .B2(n11473), .C1(n12131), .C2(n8070), .A(
        n1742), .ZN(n1737) );
  OAI22_X1 U2640 ( .A1(n11024), .A2(n12128), .B1(n11280), .B2(n12125), .ZN(
        n1742) );
  AOI221_X1 U2641 ( .B1(n12086), .B2(n11474), .C1(n12083), .C2(n8016), .A(
        n1750), .ZN(n1745) );
  OAI22_X1 U2642 ( .A1(n11025), .A2(n12080), .B1(n11281), .B2(n12077), .ZN(
        n1750) );
  AOI221_X1 U2643 ( .B1(n12134), .B2(n11475), .C1(n12131), .C2(n8072), .A(
        n1723), .ZN(n1718) );
  OAI22_X1 U2644 ( .A1(n11026), .A2(n12128), .B1(n11282), .B2(n12125), .ZN(
        n1723) );
  AOI221_X1 U2645 ( .B1(n12086), .B2(n11476), .C1(n12083), .C2(n8017), .A(
        n1731), .ZN(n1726) );
  OAI22_X1 U2646 ( .A1(n11027), .A2(n12080), .B1(n11283), .B2(n12077), .ZN(
        n1731) );
  AOI221_X1 U2647 ( .B1(n12134), .B2(n11477), .C1(n12131), .C2(n8074), .A(
        n1704), .ZN(n1699) );
  OAI22_X1 U2648 ( .A1(n11028), .A2(n12128), .B1(n11284), .B2(n12125), .ZN(
        n1704) );
  AOI221_X1 U2649 ( .B1(n12086), .B2(n11478), .C1(n12083), .C2(n8018), .A(
        n1712), .ZN(n1707) );
  OAI22_X1 U2650 ( .A1(n11029), .A2(n12080), .B1(n11285), .B2(n12077), .ZN(
        n1712) );
  AOI221_X1 U2651 ( .B1(n12134), .B2(n11479), .C1(n12131), .C2(n8076), .A(
        n1685), .ZN(n1680) );
  OAI22_X1 U2652 ( .A1(n11030), .A2(n12128), .B1(n11286), .B2(n12125), .ZN(
        n1685) );
  AOI221_X1 U2653 ( .B1(n12086), .B2(n11480), .C1(n12083), .C2(n8019), .A(
        n1693), .ZN(n1688) );
  OAI22_X1 U2654 ( .A1(n11031), .A2(n12080), .B1(n11287), .B2(n12077), .ZN(
        n1693) );
  AOI221_X1 U2655 ( .B1(n12134), .B2(n11481), .C1(n12131), .C2(n8078), .A(
        n1666), .ZN(n1661) );
  OAI22_X1 U2656 ( .A1(n11032), .A2(n12128), .B1(n11288), .B2(n12125), .ZN(
        n1666) );
  AOI221_X1 U2657 ( .B1(n12086), .B2(n11482), .C1(n12083), .C2(n8020), .A(
        n1674), .ZN(n1669) );
  OAI22_X1 U2658 ( .A1(n11033), .A2(n12080), .B1(n11289), .B2(n12077), .ZN(
        n1674) );
  AOI221_X1 U2659 ( .B1(n12134), .B2(n11483), .C1(n12131), .C2(n8080), .A(
        n1647), .ZN(n1642) );
  OAI22_X1 U2660 ( .A1(n11034), .A2(n12128), .B1(n11290), .B2(n12125), .ZN(
        n1647) );
  AOI221_X1 U2661 ( .B1(n12086), .B2(n11484), .C1(n12083), .C2(n8021), .A(
        n1655), .ZN(n1650) );
  OAI22_X1 U2662 ( .A1(n11035), .A2(n12080), .B1(n11291), .B2(n12077), .ZN(
        n1655) );
  AOI221_X1 U2663 ( .B1(n12136), .B2(n11485), .C1(n12133), .C2(n8038), .A(
        n1324), .ZN(n1319) );
  OAI22_X1 U2664 ( .A1(n11036), .A2(n12130), .B1(n11292), .B2(n12127), .ZN(
        n1324) );
  AOI221_X1 U2665 ( .B1(n12076), .B2(n8521), .C1(n12073), .C2(n8065), .A(n1333), .ZN(n1326) );
  OAI22_X1 U2666 ( .A1(n11037), .A2(n12070), .B1(n11293), .B2(n12067), .ZN(
        n1333) );
  AOI221_X1 U2667 ( .B1(n12124), .B2(n8519), .C1(n12121), .C2(n8063), .A(n1325), .ZN(n1318) );
  OAI22_X1 U2668 ( .A1(n11038), .A2(n12118), .B1(n11294), .B2(n12115), .ZN(
        n1325) );
  AOI221_X1 U2669 ( .B1(n12076), .B2(n9582), .C1(n12073), .C2(n9894), .A(n1314), .ZN(n1307) );
  OAI22_X1 U2670 ( .A1(n11039), .A2(n12070), .B1(n11295), .B2(n12067), .ZN(
        n1314) );
  AOI221_X1 U2671 ( .B1(n12124), .B2(n9580), .C1(n12121), .C2(n9892), .A(n1306), .ZN(n1299) );
  OAI22_X1 U2672 ( .A1(n11040), .A2(n12118), .B1(n11296), .B2(n12115), .ZN(
        n1306) );
  AOI221_X1 U2673 ( .B1(n12076), .B2(n9585), .C1(n12073), .C2(n9897), .A(n1295), .ZN(n1288) );
  OAI22_X1 U2674 ( .A1(n11041), .A2(n12070), .B1(n11297), .B2(n12067), .ZN(
        n1295) );
  AOI221_X1 U2675 ( .B1(n12124), .B2(n9583), .C1(n12121), .C2(n9895), .A(n1287), .ZN(n1280) );
  OAI22_X1 U2676 ( .A1(n11042), .A2(n12118), .B1(n11298), .B2(n12115), .ZN(
        n1287) );
  AOI221_X1 U2677 ( .B1(n12076), .B2(n9588), .C1(n12073), .C2(n9900), .A(n1276), .ZN(n1269) );
  OAI22_X1 U2678 ( .A1(n11043), .A2(n12070), .B1(n11299), .B2(n12067), .ZN(
        n1276) );
  AOI221_X1 U2679 ( .B1(n12124), .B2(n9586), .C1(n12121), .C2(n9898), .A(n1268), .ZN(n1261) );
  OAI22_X1 U2680 ( .A1(n11044), .A2(n12118), .B1(n11300), .B2(n12115), .ZN(
        n1268) );
  AOI221_X1 U2681 ( .B1(n12076), .B2(n9591), .C1(n12073), .C2(n9903), .A(n1257), .ZN(n1250) );
  OAI22_X1 U2682 ( .A1(n11045), .A2(n12070), .B1(n11301), .B2(n12067), .ZN(
        n1257) );
  AOI221_X1 U2683 ( .B1(n12124), .B2(n9589), .C1(n12121), .C2(n9901), .A(n1249), .ZN(n1242) );
  OAI22_X1 U2684 ( .A1(n11046), .A2(n12118), .B1(n11302), .B2(n12115), .ZN(
        n1249) );
  AOI221_X1 U2685 ( .B1(n12076), .B2(n9594), .C1(n12073), .C2(n9906), .A(n1238), .ZN(n1231) );
  OAI22_X1 U2686 ( .A1(n11047), .A2(n12070), .B1(n11303), .B2(n12067), .ZN(
        n1238) );
  AOI221_X1 U2687 ( .B1(n12124), .B2(n9592), .C1(n12121), .C2(n9904), .A(n1230), .ZN(n1223) );
  OAI22_X1 U2688 ( .A1(n11048), .A2(n12118), .B1(n11304), .B2(n12115), .ZN(
        n1230) );
  AOI221_X1 U2689 ( .B1(n12076), .B2(n9597), .C1(n12073), .C2(n9909), .A(n1219), .ZN(n1212) );
  OAI22_X1 U2690 ( .A1(n11049), .A2(n12070), .B1(n11305), .B2(n12067), .ZN(
        n1219) );
  AOI221_X1 U2691 ( .B1(n12124), .B2(n9595), .C1(n12121), .C2(n9907), .A(n1211), .ZN(n1204) );
  OAI22_X1 U2692 ( .A1(n11050), .A2(n12118), .B1(n11306), .B2(n12115), .ZN(
        n1211) );
  AOI221_X1 U2693 ( .B1(n12076), .B2(n9600), .C1(n12073), .C2(n9912), .A(n1198), .ZN(n1177) );
  OAI22_X1 U2694 ( .A1(n11051), .A2(n12070), .B1(n11307), .B2(n12067), .ZN(
        n1198) );
  AOI221_X1 U2695 ( .B1(n12124), .B2(n9598), .C1(n12121), .C2(n9910), .A(n1174), .ZN(n1153) );
  OAI22_X1 U2696 ( .A1(n11052), .A2(n12118), .B1(n11308), .B2(n12115), .ZN(
        n1174) );
  AND2_X1 U2697 ( .A1(ADD_RD1[2]), .A2(n12573), .ZN(n1781) );
  OAI221_X1 U2698 ( .B1(n12551), .B2(n12167), .C1(n4172), .C2(n12166), .A(
        n1771), .ZN(n2571) );
  OAI21_X1 U2699 ( .B1(n1772), .B2(n1773), .A(n12161), .ZN(n1771) );
  NAND4_X1 U2700 ( .A1(n1791), .A2(n1792), .A3(n1793), .A4(n1794), .ZN(n1772)
         );
  NAND4_X1 U2701 ( .A1(n1775), .A2(n1776), .A3(n1777), .A4(n1778), .ZN(n1773)
         );
  OAI221_X1 U2702 ( .B1(n12539), .B2(n12167), .C1(n4173), .C2(n12166), .A(
        n1752), .ZN(n2572) );
  OAI21_X1 U2703 ( .B1(n1753), .B2(n1754), .A(n12161), .ZN(n1752) );
  NAND4_X1 U2704 ( .A1(n1763), .A2(n1764), .A3(n1765), .A4(n1766), .ZN(n1753)
         );
  NAND4_X1 U2705 ( .A1(n1755), .A2(n1756), .A3(n1757), .A4(n1758), .ZN(n1754)
         );
  OAI221_X1 U2706 ( .B1(n12536), .B2(n12167), .C1(n4174), .C2(n12166), .A(
        n1733), .ZN(n2573) );
  OAI21_X1 U2707 ( .B1(n1734), .B2(n1735), .A(n12161), .ZN(n1733) );
  NAND4_X1 U2708 ( .A1(n1744), .A2(n1745), .A3(n1746), .A4(n1747), .ZN(n1734)
         );
  NAND4_X1 U2709 ( .A1(n1736), .A2(n1737), .A3(n1738), .A4(n1739), .ZN(n1735)
         );
  OAI221_X1 U2710 ( .B1(n12533), .B2(n12167), .C1(n4175), .C2(n12166), .A(
        n1714), .ZN(n2574) );
  OAI21_X1 U2711 ( .B1(n1715), .B2(n1716), .A(n12161), .ZN(n1714) );
  NAND4_X1 U2712 ( .A1(n1725), .A2(n1726), .A3(n1727), .A4(n1728), .ZN(n1715)
         );
  NAND4_X1 U2713 ( .A1(n1717), .A2(n1718), .A3(n1719), .A4(n1720), .ZN(n1716)
         );
  OAI221_X1 U2714 ( .B1(n12530), .B2(n12167), .C1(n4176), .C2(n12166), .A(
        n1695), .ZN(n2575) );
  OAI21_X1 U2715 ( .B1(n1696), .B2(n1697), .A(n12161), .ZN(n1695) );
  NAND4_X1 U2716 ( .A1(n1706), .A2(n1707), .A3(n1708), .A4(n1709), .ZN(n1696)
         );
  NAND4_X1 U2717 ( .A1(n1698), .A2(n1699), .A3(n1700), .A4(n1701), .ZN(n1697)
         );
  OAI221_X1 U2718 ( .B1(n12527), .B2(n12167), .C1(n4177), .C2(n12166), .A(
        n1676), .ZN(n2576) );
  OAI21_X1 U2719 ( .B1(n1677), .B2(n1678), .A(n12161), .ZN(n1676) );
  NAND4_X1 U2720 ( .A1(n1687), .A2(n1688), .A3(n1689), .A4(n1690), .ZN(n1677)
         );
  NAND4_X1 U2721 ( .A1(n1679), .A2(n1680), .A3(n1681), .A4(n1682), .ZN(n1678)
         );
  OAI221_X1 U2722 ( .B1(n12524), .B2(n12167), .C1(n4178), .C2(n12166), .A(
        n1657), .ZN(n2577) );
  OAI21_X1 U2723 ( .B1(n1658), .B2(n1659), .A(n12161), .ZN(n1657) );
  NAND4_X1 U2724 ( .A1(n1668), .A2(n1669), .A3(n1670), .A4(n1671), .ZN(n1658)
         );
  NAND4_X1 U2725 ( .A1(n1660), .A2(n1661), .A3(n1662), .A4(n1663), .ZN(n1659)
         );
  OAI221_X1 U2726 ( .B1(n12521), .B2(n12167), .C1(n4179), .C2(n12166), .A(
        n1638), .ZN(n2578) );
  OAI21_X1 U2727 ( .B1(n1639), .B2(n1640), .A(n12161), .ZN(n1638) );
  NAND4_X1 U2728 ( .A1(n1649), .A2(n1650), .A3(n1651), .A4(n1652), .ZN(n1639)
         );
  NAND4_X1 U2729 ( .A1(n1641), .A2(n1642), .A3(n1643), .A4(n1644), .ZN(n1640)
         );
  OAI221_X1 U2730 ( .B1(n12518), .B2(n12167), .C1(n4180), .C2(n12166), .A(
        n1619), .ZN(n2579) );
  OAI21_X1 U2731 ( .B1(n1620), .B2(n1621), .A(n12161), .ZN(n1619) );
  NAND4_X1 U2732 ( .A1(n1630), .A2(n1631), .A3(n1632), .A4(n1633), .ZN(n1620)
         );
  NAND4_X1 U2733 ( .A1(n1622), .A2(n1623), .A3(n1624), .A4(n1625), .ZN(n1621)
         );
  OAI221_X1 U2734 ( .B1(n12515), .B2(n12167), .C1(n4181), .C2(n12165), .A(
        n1600), .ZN(n2580) );
  OAI21_X1 U2735 ( .B1(n1601), .B2(n1602), .A(n12161), .ZN(n1600) );
  NAND4_X1 U2736 ( .A1(n1611), .A2(n1612), .A3(n1613), .A4(n1614), .ZN(n1601)
         );
  NAND4_X1 U2737 ( .A1(n1603), .A2(n1604), .A3(n1605), .A4(n1606), .ZN(n1602)
         );
  OAI221_X1 U2738 ( .B1(n12512), .B2(n12167), .C1(n4182), .C2(n12165), .A(
        n1581), .ZN(n2581) );
  OAI21_X1 U2739 ( .B1(n1582), .B2(n1583), .A(n12161), .ZN(n1581) );
  NAND4_X1 U2740 ( .A1(n1592), .A2(n1593), .A3(n1594), .A4(n1595), .ZN(n1582)
         );
  NAND4_X1 U2741 ( .A1(n1584), .A2(n1585), .A3(n1586), .A4(n1587), .ZN(n1583)
         );
  OAI221_X1 U2742 ( .B1(n12476), .B2(n12169), .C1(n4194), .C2(n12164), .A(
        n1353), .ZN(n2593) );
  OAI21_X1 U2743 ( .B1(n1354), .B2(n1355), .A(n12163), .ZN(n1353) );
  NAND4_X1 U2744 ( .A1(n1364), .A2(n1365), .A3(n1366), .A4(n1367), .ZN(n1354)
         );
  NAND4_X1 U2745 ( .A1(n1356), .A2(n1357), .A3(n1358), .A4(n1359), .ZN(n1355)
         );
  OAI221_X1 U2746 ( .B1(n12470), .B2(n12169), .C1(n4196), .C2(n12164), .A(
        n1315), .ZN(n2595) );
  OAI21_X1 U2747 ( .B1(n1316), .B2(n1317), .A(n12163), .ZN(n1315) );
  NAND4_X1 U2748 ( .A1(n1318), .A2(n1319), .A3(n1320), .A4(n1321), .ZN(n1317)
         );
  NAND4_X1 U2749 ( .A1(n1326), .A2(n1327), .A3(n1328), .A4(n1329), .ZN(n1316)
         );
  OAI221_X1 U2750 ( .B1(n12509), .B2(n12168), .C1(n4183), .C2(n12165), .A(
        n1562), .ZN(n2582) );
  OAI21_X1 U2751 ( .B1(n1563), .B2(n1564), .A(n12162), .ZN(n1562) );
  NAND4_X1 U2752 ( .A1(n1573), .A2(n1574), .A3(n1575), .A4(n1576), .ZN(n1563)
         );
  NAND4_X1 U2753 ( .A1(n1565), .A2(n1566), .A3(n1567), .A4(n1568), .ZN(n1564)
         );
  OAI221_X1 U2754 ( .B1(n12506), .B2(n12168), .C1(n4184), .C2(n12165), .A(
        n1543), .ZN(n2583) );
  OAI21_X1 U2755 ( .B1(n1544), .B2(n1545), .A(n12162), .ZN(n1543) );
  NAND4_X1 U2756 ( .A1(n1554), .A2(n1555), .A3(n1556), .A4(n1557), .ZN(n1544)
         );
  NAND4_X1 U2757 ( .A1(n1546), .A2(n1547), .A3(n1548), .A4(n1549), .ZN(n1545)
         );
  OAI221_X1 U2758 ( .B1(n12494), .B2(n12168), .C1(n4188), .C2(n12165), .A(
        n1467), .ZN(n2587) );
  OAI21_X1 U2759 ( .B1(n1468), .B2(n1469), .A(n12162), .ZN(n1467) );
  NAND4_X1 U2760 ( .A1(n1478), .A2(n1479), .A3(n1480), .A4(n1481), .ZN(n1468)
         );
  NAND4_X1 U2761 ( .A1(n1470), .A2(n1471), .A3(n1472), .A4(n1473), .ZN(n1469)
         );
  OAI221_X1 U2762 ( .B1(n12491), .B2(n12168), .C1(n4189), .C2(n12165), .A(
        n1448), .ZN(n2588) );
  OAI21_X1 U2763 ( .B1(n1449), .B2(n1450), .A(n12162), .ZN(n1448) );
  NAND4_X1 U2764 ( .A1(n1459), .A2(n1460), .A3(n1461), .A4(n1462), .ZN(n1449)
         );
  NAND4_X1 U2765 ( .A1(n1451), .A2(n1452), .A3(n1453), .A4(n1454), .ZN(n1450)
         );
  OAI221_X1 U2766 ( .B1(n12488), .B2(n12168), .C1(n4190), .C2(n12165), .A(
        n1429), .ZN(n2589) );
  OAI21_X1 U2767 ( .B1(n1430), .B2(n1431), .A(n12162), .ZN(n1429) );
  NAND4_X1 U2768 ( .A1(n1440), .A2(n1441), .A3(n1442), .A4(n1443), .ZN(n1430)
         );
  NAND4_X1 U2769 ( .A1(n1432), .A2(n1433), .A3(n1434), .A4(n1435), .ZN(n1431)
         );
  OAI221_X1 U2770 ( .B1(n12485), .B2(n12168), .C1(n4191), .C2(n12165), .A(
        n1410), .ZN(n2590) );
  OAI21_X1 U2771 ( .B1(n1411), .B2(n1412), .A(n12162), .ZN(n1410) );
  NAND4_X1 U2772 ( .A1(n1421), .A2(n1422), .A3(n1423), .A4(n1424), .ZN(n1411)
         );
  NAND4_X1 U2773 ( .A1(n1413), .A2(n1414), .A3(n1415), .A4(n1416), .ZN(n1412)
         );
  OAI221_X1 U2774 ( .B1(n12482), .B2(n12168), .C1(n4192), .C2(n12164), .A(
        n1391), .ZN(n2591) );
  OAI21_X1 U2775 ( .B1(n1392), .B2(n1393), .A(n12162), .ZN(n1391) );
  NAND4_X1 U2776 ( .A1(n1402), .A2(n1403), .A3(n1404), .A4(n1405), .ZN(n1392)
         );
  NAND4_X1 U2777 ( .A1(n1394), .A2(n1395), .A3(n1396), .A4(n1397), .ZN(n1393)
         );
  OAI221_X1 U2778 ( .B1(n12479), .B2(n12168), .C1(n4193), .C2(n12164), .A(
        n1372), .ZN(n2592) );
  OAI21_X1 U2779 ( .B1(n1373), .B2(n1374), .A(n12162), .ZN(n1372) );
  NAND4_X1 U2780 ( .A1(n1383), .A2(n1384), .A3(n1385), .A4(n1386), .ZN(n1373)
         );
  NAND4_X1 U2781 ( .A1(n1375), .A2(n1376), .A3(n1377), .A4(n1378), .ZN(n1374)
         );
  AOI221_X1 U2782 ( .B1(n12100), .B2(n8469), .C1(n12097), .C2(n8013), .A(n1331), .ZN(n1328) );
  OAI22_X1 U2783 ( .A1(n11053), .A2(n12094), .B1(n11309), .B2(n12091), .ZN(
        n1331) );
  AOI221_X1 U2784 ( .B1(n12100), .B2(n9581), .C1(n12097), .C2(n9893), .A(n1312), .ZN(n1309) );
  OAI22_X1 U2785 ( .A1(n11054), .A2(n12094), .B1(n11310), .B2(n12091), .ZN(
        n1312) );
  AOI221_X1 U2786 ( .B1(n12100), .B2(n9584), .C1(n12097), .C2(n9896), .A(n1293), .ZN(n1290) );
  OAI22_X1 U2787 ( .A1(n11055), .A2(n12094), .B1(n11311), .B2(n12091), .ZN(
        n1293) );
  AOI221_X1 U2788 ( .B1(n12100), .B2(n9587), .C1(n12097), .C2(n9899), .A(n1274), .ZN(n1271) );
  OAI22_X1 U2789 ( .A1(n11056), .A2(n12094), .B1(n11312), .B2(n12091), .ZN(
        n1274) );
  AOI221_X1 U2790 ( .B1(n12100), .B2(n9590), .C1(n12097), .C2(n9902), .A(n1255), .ZN(n1252) );
  OAI22_X1 U2791 ( .A1(n11057), .A2(n12094), .B1(n11313), .B2(n12091), .ZN(
        n1255) );
  AOI221_X1 U2792 ( .B1(n12100), .B2(n9593), .C1(n12097), .C2(n9905), .A(n1236), .ZN(n1233) );
  OAI22_X1 U2793 ( .A1(n11058), .A2(n12094), .B1(n11314), .B2(n12091), .ZN(
        n1236) );
  AOI221_X1 U2794 ( .B1(n12100), .B2(n9596), .C1(n12097), .C2(n9908), .A(n1217), .ZN(n1214) );
  OAI22_X1 U2795 ( .A1(n11059), .A2(n12094), .B1(n11315), .B2(n12091), .ZN(
        n1217) );
  AOI221_X1 U2796 ( .B1(n12100), .B2(n9599), .C1(n12097), .C2(n9911), .A(n1188), .ZN(n1179) );
  OAI22_X1 U2797 ( .A1(n11060), .A2(n12094), .B1(n11316), .B2(n12091), .ZN(
        n1188) );
  AOI221_X1 U2798 ( .B1(n12088), .B2(n8520), .C1(n12085), .C2(n8064), .A(n1332), .ZN(n1327) );
  OAI22_X1 U2799 ( .A1(n11061), .A2(n12082), .B1(n11317), .B2(n12079), .ZN(
        n1332) );
  AOI221_X1 U2800 ( .B1(n12088), .B2(n9560), .C1(n12085), .C2(n9872), .A(n1313), .ZN(n1308) );
  OAI22_X1 U2801 ( .A1(n11062), .A2(n12082), .B1(n11318), .B2(n12079), .ZN(
        n1313) );
  AOI221_X1 U2802 ( .B1(n12088), .B2(n9562), .C1(n12085), .C2(n9874), .A(n1294), .ZN(n1289) );
  OAI22_X1 U2803 ( .A1(n11063), .A2(n12082), .B1(n11319), .B2(n12079), .ZN(
        n1294) );
  AOI221_X1 U2804 ( .B1(n12088), .B2(n9564), .C1(n12085), .C2(n9876), .A(n1275), .ZN(n1270) );
  OAI22_X1 U2805 ( .A1(n11064), .A2(n12082), .B1(n11320), .B2(n12079), .ZN(
        n1275) );
  AOI221_X1 U2806 ( .B1(n12088), .B2(n9566), .C1(n12085), .C2(n9878), .A(n1256), .ZN(n1251) );
  OAI22_X1 U2807 ( .A1(n11065), .A2(n12082), .B1(n11321), .B2(n12079), .ZN(
        n1256) );
  AOI221_X1 U2808 ( .B1(n12088), .B2(n9568), .C1(n12085), .C2(n9880), .A(n1237), .ZN(n1232) );
  OAI22_X1 U2809 ( .A1(n11066), .A2(n12082), .B1(n11322), .B2(n12079), .ZN(
        n1237) );
  AOI221_X1 U2810 ( .B1(n12088), .B2(n9570), .C1(n12085), .C2(n9882), .A(n1218), .ZN(n1213) );
  OAI22_X1 U2811 ( .A1(n11067), .A2(n12082), .B1(n11323), .B2(n12079), .ZN(
        n1218) );
  AOI221_X1 U2812 ( .B1(n12088), .B2(n9572), .C1(n12085), .C2(n9884), .A(n1193), .ZN(n1178) );
  OAI22_X1 U2813 ( .A1(n11068), .A2(n12082), .B1(n11324), .B2(n12079), .ZN(
        n1193) );
  AOI221_X1 U2814 ( .B1(n12112), .B2(n8419), .C1(n12109), .C2(n7963), .A(n1330), .ZN(n1329) );
  OAI22_X1 U2815 ( .A1(n11069), .A2(n12106), .B1(n11325), .B2(n12103), .ZN(
        n1330) );
  AOI221_X1 U2816 ( .B1(n12160), .B2(n11486), .C1(n12157), .C2(n7962), .A(
        n1322), .ZN(n1321) );
  OAI22_X1 U2817 ( .A1(n11070), .A2(n12154), .B1(n11326), .B2(n12151), .ZN(
        n1322) );
  AOI221_X1 U2818 ( .B1(n12112), .B2(n9552), .C1(n12109), .C2(n9864), .A(n1311), .ZN(n1310) );
  OAI22_X1 U2819 ( .A1(n11071), .A2(n12106), .B1(n11327), .B2(n12103), .ZN(
        n1311) );
  AOI221_X1 U2820 ( .B1(n12160), .B2(n9601), .C1(n12157), .C2(n9913), .A(n1303), .ZN(n1302) );
  OAI22_X1 U2821 ( .A1(n11072), .A2(n12154), .B1(n11328), .B2(n12151), .ZN(
        n1303) );
  AOI221_X1 U2822 ( .B1(n12112), .B2(n9553), .C1(n12109), .C2(n9865), .A(n1292), .ZN(n1291) );
  OAI22_X1 U2823 ( .A1(n11073), .A2(n12106), .B1(n11329), .B2(n12103), .ZN(
        n1292) );
  AOI221_X1 U2824 ( .B1(n12160), .B2(n9602), .C1(n12157), .C2(n9914), .A(n1284), .ZN(n1283) );
  OAI22_X1 U2825 ( .A1(n11074), .A2(n12154), .B1(n11330), .B2(n12151), .ZN(
        n1284) );
  AOI221_X1 U2826 ( .B1(n12112), .B2(n9554), .C1(n12109), .C2(n9866), .A(n1273), .ZN(n1272) );
  OAI22_X1 U2827 ( .A1(n11075), .A2(n12106), .B1(n11331), .B2(n12103), .ZN(
        n1273) );
  AOI221_X1 U2828 ( .B1(n12160), .B2(n9603), .C1(n12157), .C2(n9915), .A(n1265), .ZN(n1264) );
  OAI22_X1 U2829 ( .A1(n11076), .A2(n12154), .B1(n11332), .B2(n12151), .ZN(
        n1265) );
  AOI221_X1 U2830 ( .B1(n12112), .B2(n9555), .C1(n12109), .C2(n9867), .A(n1254), .ZN(n1253) );
  OAI22_X1 U2831 ( .A1(n11077), .A2(n12106), .B1(n11333), .B2(n12103), .ZN(
        n1254) );
  AOI221_X1 U2832 ( .B1(n12160), .B2(n9604), .C1(n12157), .C2(n9916), .A(n1246), .ZN(n1245) );
  OAI22_X1 U2833 ( .A1(n11078), .A2(n12154), .B1(n11334), .B2(n12151), .ZN(
        n1246) );
  AOI221_X1 U2834 ( .B1(n12112), .B2(n9556), .C1(n12109), .C2(n9868), .A(n1235), .ZN(n1234) );
  OAI22_X1 U2835 ( .A1(n11079), .A2(n12106), .B1(n11335), .B2(n12103), .ZN(
        n1235) );
  AOI221_X1 U2836 ( .B1(n12160), .B2(n9605), .C1(n12157), .C2(n9917), .A(n1227), .ZN(n1226) );
  OAI22_X1 U2837 ( .A1(n11080), .A2(n12154), .B1(n11336), .B2(n12151), .ZN(
        n1227) );
  AOI221_X1 U2838 ( .B1(n12112), .B2(n9557), .C1(n12109), .C2(n9869), .A(n1216), .ZN(n1215) );
  OAI22_X1 U2839 ( .A1(n11081), .A2(n12106), .B1(n11337), .B2(n12103), .ZN(
        n1216) );
  AOI221_X1 U2840 ( .B1(n12160), .B2(n9606), .C1(n12157), .C2(n9918), .A(n1208), .ZN(n1207) );
  OAI22_X1 U2841 ( .A1(n11082), .A2(n12154), .B1(n11338), .B2(n12151), .ZN(
        n1208) );
  AOI221_X1 U2842 ( .B1(n12112), .B2(n9558), .C1(n12109), .C2(n9870), .A(n1183), .ZN(n1180) );
  OAI22_X1 U2843 ( .A1(n11083), .A2(n12106), .B1(n11339), .B2(n12103), .ZN(
        n1183) );
  AOI221_X1 U2844 ( .B1(n12160), .B2(n9607), .C1(n12157), .C2(n9919), .A(n1159), .ZN(n1156) );
  OAI22_X1 U2845 ( .A1(n11084), .A2(n12154), .B1(n11340), .B2(n12151), .ZN(
        n1159) );
  AOI221_X1 U2846 ( .B1(n12158), .B2(n11487), .C1(n12155), .C2(n7914), .A(
        n1779), .ZN(n1778) );
  OAI22_X1 U2847 ( .A1(n11085), .A2(n12152), .B1(n11341), .B2(n12149), .ZN(
        n1779) );
  AOI221_X1 U2848 ( .B1(n12146), .B2(n11488), .C1(n12143), .C2(n7964), .A(
        n1784), .ZN(n1777) );
  OAI22_X1 U2849 ( .A1(n11086), .A2(n12140), .B1(n11342), .B2(n12137), .ZN(
        n1784) );
  AOI221_X1 U2850 ( .B1(n12122), .B2(n11489), .C1(n12119), .C2(n8067), .A(
        n1790), .ZN(n1775) );
  OAI22_X1 U2851 ( .A1(n11087), .A2(n12116), .B1(n11343), .B2(n12113), .ZN(
        n1790) );
  AOI221_X1 U2852 ( .B1(n12074), .B2(n11490), .C1(n12071), .C2(n8039), .A(
        n1802), .ZN(n1791) );
  OAI22_X1 U2853 ( .A1(n11088), .A2(n12068), .B1(n11344), .B2(n12065), .ZN(
        n1802) );
  AOI221_X1 U2854 ( .B1(n12158), .B2(n11491), .C1(n12155), .C2(n7916), .A(
        n1759), .ZN(n1758) );
  OAI22_X1 U2855 ( .A1(n11089), .A2(n12152), .B1(n11345), .B2(n12149), .ZN(
        n1759) );
  AOI221_X1 U2856 ( .B1(n12146), .B2(n11492), .C1(n12143), .C2(n7966), .A(
        n1760), .ZN(n1757) );
  OAI22_X1 U2857 ( .A1(n11090), .A2(n12140), .B1(n11346), .B2(n12137), .ZN(
        n1760) );
  AOI221_X1 U2858 ( .B1(n12122), .B2(n11493), .C1(n12119), .C2(n8069), .A(
        n1762), .ZN(n1755) );
  OAI22_X1 U2859 ( .A1(n11091), .A2(n12116), .B1(n11347), .B2(n12113), .ZN(
        n1762) );
  AOI221_X1 U2860 ( .B1(n12074), .B2(n11494), .C1(n12071), .C2(n8040), .A(
        n1770), .ZN(n1763) );
  OAI22_X1 U2861 ( .A1(n11092), .A2(n12068), .B1(n11348), .B2(n12065), .ZN(
        n1770) );
  AOI221_X1 U2862 ( .B1(n12158), .B2(n11495), .C1(n12155), .C2(n7918), .A(
        n1740), .ZN(n1739) );
  OAI22_X1 U2863 ( .A1(n11093), .A2(n12152), .B1(n11349), .B2(n12149), .ZN(
        n1740) );
  AOI221_X1 U2864 ( .B1(n12146), .B2(n11496), .C1(n12143), .C2(n7968), .A(
        n1741), .ZN(n1738) );
  OAI22_X1 U2865 ( .A1(n11094), .A2(n12140), .B1(n11350), .B2(n12137), .ZN(
        n1741) );
  AOI221_X1 U2866 ( .B1(n12122), .B2(n11497), .C1(n12119), .C2(n8071), .A(
        n1743), .ZN(n1736) );
  OAI22_X1 U2867 ( .A1(n11095), .A2(n12116), .B1(n11351), .B2(n12113), .ZN(
        n1743) );
  AOI221_X1 U2868 ( .B1(n12074), .B2(n11498), .C1(n12071), .C2(n8041), .A(
        n1751), .ZN(n1744) );
  OAI22_X1 U2869 ( .A1(n11096), .A2(n12068), .B1(n11352), .B2(n12065), .ZN(
        n1751) );
  AOI221_X1 U2870 ( .B1(n12158), .B2(n11499), .C1(n12155), .C2(n7920), .A(
        n1721), .ZN(n1720) );
  OAI22_X1 U2871 ( .A1(n11097), .A2(n12152), .B1(n11353), .B2(n12149), .ZN(
        n1721) );
  AOI221_X1 U2872 ( .B1(n12146), .B2(n11500), .C1(n12143), .C2(n7970), .A(
        n1722), .ZN(n1719) );
  OAI22_X1 U2873 ( .A1(n11098), .A2(n12140), .B1(n11354), .B2(n12137), .ZN(
        n1722) );
  AOI221_X1 U2874 ( .B1(n12122), .B2(n11501), .C1(n12119), .C2(n8073), .A(
        n1724), .ZN(n1717) );
  OAI22_X1 U2875 ( .A1(n11099), .A2(n12116), .B1(n11355), .B2(n12113), .ZN(
        n1724) );
  AOI221_X1 U2876 ( .B1(n12074), .B2(n11502), .C1(n12071), .C2(n8042), .A(
        n1732), .ZN(n1725) );
  OAI22_X1 U2877 ( .A1(n11100), .A2(n12068), .B1(n11356), .B2(n12065), .ZN(
        n1732) );
  AOI221_X1 U2878 ( .B1(n12158), .B2(n11503), .C1(n12155), .C2(n7922), .A(
        n1702), .ZN(n1701) );
  OAI22_X1 U2879 ( .A1(n11101), .A2(n12152), .B1(n11357), .B2(n12149), .ZN(
        n1702) );
  AOI221_X1 U2880 ( .B1(n12146), .B2(n11504), .C1(n12143), .C2(n7972), .A(
        n1703), .ZN(n1700) );
  OAI22_X1 U2881 ( .A1(n11102), .A2(n12140), .B1(n11358), .B2(n12137), .ZN(
        n1703) );
  AOI221_X1 U2882 ( .B1(n12122), .B2(n11505), .C1(n12119), .C2(n8075), .A(
        n1705), .ZN(n1698) );
  OAI22_X1 U2883 ( .A1(n11103), .A2(n12116), .B1(n11359), .B2(n12113), .ZN(
        n1705) );
  AOI221_X1 U2884 ( .B1(n12074), .B2(n11506), .C1(n12071), .C2(n8043), .A(
        n1713), .ZN(n1706) );
  OAI22_X1 U2885 ( .A1(n11104), .A2(n12068), .B1(n11360), .B2(n12065), .ZN(
        n1713) );
  AOI221_X1 U2886 ( .B1(n12158), .B2(n11507), .C1(n12155), .C2(n7924), .A(
        n1683), .ZN(n1682) );
  OAI22_X1 U2887 ( .A1(n11105), .A2(n12152), .B1(n11361), .B2(n12149), .ZN(
        n1683) );
  AOI221_X1 U2888 ( .B1(n12146), .B2(n11508), .C1(n12143), .C2(n7974), .A(
        n1684), .ZN(n1681) );
  OAI22_X1 U2889 ( .A1(n11106), .A2(n12140), .B1(n11362), .B2(n12137), .ZN(
        n1684) );
  AOI221_X1 U2890 ( .B1(n12122), .B2(n11509), .C1(n12119), .C2(n8077), .A(
        n1686), .ZN(n1679) );
  OAI22_X1 U2891 ( .A1(n11107), .A2(n12116), .B1(n11363), .B2(n12113), .ZN(
        n1686) );
  AOI221_X1 U2892 ( .B1(n12074), .B2(n11510), .C1(n12071), .C2(n8044), .A(
        n1694), .ZN(n1687) );
  OAI22_X1 U2893 ( .A1(n11108), .A2(n12068), .B1(n11364), .B2(n12065), .ZN(
        n1694) );
  AOI221_X1 U2894 ( .B1(n12158), .B2(n11511), .C1(n12155), .C2(n7926), .A(
        n1664), .ZN(n1663) );
  OAI22_X1 U2895 ( .A1(n11109), .A2(n12152), .B1(n11365), .B2(n12149), .ZN(
        n1664) );
  AOI221_X1 U2896 ( .B1(n12146), .B2(n11512), .C1(n12143), .C2(n7976), .A(
        n1665), .ZN(n1662) );
  OAI22_X1 U2897 ( .A1(n11110), .A2(n12140), .B1(n11366), .B2(n12137), .ZN(
        n1665) );
  AOI221_X1 U2898 ( .B1(n12122), .B2(n11513), .C1(n12119), .C2(n8079), .A(
        n1667), .ZN(n1660) );
  OAI22_X1 U2899 ( .A1(n11111), .A2(n12116), .B1(n11367), .B2(n12113), .ZN(
        n1667) );
  AOI221_X1 U2900 ( .B1(n12074), .B2(n11514), .C1(n12071), .C2(n8045), .A(
        n1675), .ZN(n1668) );
  OAI22_X1 U2901 ( .A1(n11112), .A2(n12068), .B1(n11368), .B2(n12065), .ZN(
        n1675) );
  AOI221_X1 U2902 ( .B1(n12158), .B2(n11515), .C1(n12155), .C2(n7928), .A(
        n1645), .ZN(n1644) );
  OAI22_X1 U2903 ( .A1(n11113), .A2(n12152), .B1(n11369), .B2(n12149), .ZN(
        n1645) );
  AOI221_X1 U2904 ( .B1(n12146), .B2(n11516), .C1(n12143), .C2(n7978), .A(
        n1646), .ZN(n1643) );
  OAI22_X1 U2905 ( .A1(n11114), .A2(n12140), .B1(n11370), .B2(n12137), .ZN(
        n1646) );
  AOI221_X1 U2906 ( .B1(n12122), .B2(n11517), .C1(n12119), .C2(n8081), .A(
        n1648), .ZN(n1641) );
  OAI22_X1 U2907 ( .A1(n11115), .A2(n12116), .B1(n11371), .B2(n12113), .ZN(
        n1648) );
  AOI221_X1 U2908 ( .B1(n12074), .B2(n11518), .C1(n12071), .C2(n8046), .A(
        n1656), .ZN(n1649) );
  OAI22_X1 U2909 ( .A1(n11116), .A2(n12068), .B1(n11372), .B2(n12065), .ZN(
        n1656) );
  AOI221_X1 U2910 ( .B1(n12158), .B2(n8386), .C1(n12155), .C2(n7930), .A(n1626), .ZN(n1625) );
  OAI22_X1 U2911 ( .A1(n11117), .A2(n12152), .B1(n11373), .B2(n12149), .ZN(
        n1626) );
  AOI221_X1 U2912 ( .B1(n12122), .B2(n8539), .C1(n12119), .C2(n8083), .A(n1629), .ZN(n1622) );
  OAI22_X1 U2913 ( .A1(n11118), .A2(n12116), .B1(n11374), .B2(n12113), .ZN(
        n1629) );
  AOI221_X1 U2914 ( .B1(n12110), .B2(n8387), .C1(n12107), .C2(n7931), .A(n1634), .ZN(n1633) );
  OAI22_X1 U2915 ( .A1(n11119), .A2(n12104), .B1(n11375), .B2(n12101), .ZN(
        n1634) );
  AOI221_X1 U2916 ( .B1(n12074), .B2(n8503), .C1(n12071), .C2(n8047), .A(n1637), .ZN(n1630) );
  OAI22_X1 U2917 ( .A1(n11120), .A2(n12068), .B1(n11376), .B2(n12065), .ZN(
        n1637) );
  AOI221_X1 U2918 ( .B1(n12134), .B2(n8540), .C1(n12131), .C2(n8084), .A(n1609), .ZN(n1604) );
  OAI22_X1 U2919 ( .A1(n11121), .A2(n12128), .B1(n11377), .B2(n12125), .ZN(
        n1609) );
  AOI221_X1 U2920 ( .B1(n12158), .B2(n8388), .C1(n12155), .C2(n7932), .A(n1607), .ZN(n1606) );
  OAI22_X1 U2921 ( .A1(n11122), .A2(n12152), .B1(n11378), .B2(n12149), .ZN(
        n1607) );
  AOI221_X1 U2922 ( .B1(n12146), .B2(n8438), .C1(n12143), .C2(n7982), .A(n1608), .ZN(n1605) );
  OAI22_X1 U2923 ( .A1(n11123), .A2(n12140), .B1(n11379), .B2(n12137), .ZN(
        n1608) );
  AOI221_X1 U2924 ( .B1(n12122), .B2(n8541), .C1(n12119), .C2(n8085), .A(n1610), .ZN(n1603) );
  OAI22_X1 U2925 ( .A1(n11124), .A2(n12116), .B1(n11380), .B2(n12113), .ZN(
        n1610) );
  AOI221_X1 U2926 ( .B1(n12074), .B2(n8504), .C1(n12071), .C2(n8048), .A(n1618), .ZN(n1611) );
  OAI22_X1 U2927 ( .A1(n11125), .A2(n12068), .B1(n11381), .B2(n12065), .ZN(
        n1618) );
  AOI221_X1 U2928 ( .B1(n12134), .B2(n8542), .C1(n12131), .C2(n8086), .A(n1590), .ZN(n1585) );
  OAI22_X1 U2929 ( .A1(n11126), .A2(n12128), .B1(n11382), .B2(n12125), .ZN(
        n1590) );
  AOI221_X1 U2930 ( .B1(n12158), .B2(n8390), .C1(n12155), .C2(n7934), .A(n1588), .ZN(n1587) );
  OAI22_X1 U2931 ( .A1(n11127), .A2(n12152), .B1(n11383), .B2(n12149), .ZN(
        n1588) );
  AOI221_X1 U2932 ( .B1(n12146), .B2(n8440), .C1(n12143), .C2(n7984), .A(n1589), .ZN(n1586) );
  OAI22_X1 U2933 ( .A1(n11128), .A2(n12140), .B1(n11384), .B2(n12137), .ZN(
        n1589) );
  AOI221_X1 U2934 ( .B1(n12122), .B2(n8543), .C1(n12119), .C2(n8087), .A(n1591), .ZN(n1584) );
  OAI22_X1 U2935 ( .A1(n11129), .A2(n12116), .B1(n11385), .B2(n12113), .ZN(
        n1591) );
  AOI221_X1 U2936 ( .B1(n12074), .B2(n8505), .C1(n12071), .C2(n8049), .A(n1599), .ZN(n1592) );
  OAI22_X1 U2937 ( .A1(n11130), .A2(n12068), .B1(n11386), .B2(n12065), .ZN(
        n1599) );
  AOI221_X1 U2938 ( .B1(n12135), .B2(n8544), .C1(n12132), .C2(n8088), .A(n1571), .ZN(n1566) );
  OAI22_X1 U2939 ( .A1(n11131), .A2(n12128), .B1(n11387), .B2(n12125), .ZN(
        n1571) );
  AOI221_X1 U2940 ( .B1(n12159), .B2(n8392), .C1(n12156), .C2(n7936), .A(n1569), .ZN(n1568) );
  OAI22_X1 U2941 ( .A1(n11132), .A2(n12152), .B1(n11388), .B2(n12149), .ZN(
        n1569) );
  AOI221_X1 U2942 ( .B1(n12147), .B2(n8442), .C1(n12144), .C2(n7986), .A(n1570), .ZN(n1567) );
  OAI22_X1 U2943 ( .A1(n11133), .A2(n12140), .B1(n11389), .B2(n12137), .ZN(
        n1570) );
  AOI221_X1 U2944 ( .B1(n12123), .B2(n8545), .C1(n12120), .C2(n8089), .A(n1572), .ZN(n1565) );
  OAI22_X1 U2945 ( .A1(n11134), .A2(n12116), .B1(n11390), .B2(n12113), .ZN(
        n1572) );
  AOI221_X1 U2946 ( .B1(n12075), .B2(n8506), .C1(n12072), .C2(n8050), .A(n1580), .ZN(n1573) );
  OAI22_X1 U2947 ( .A1(n11135), .A2(n12068), .B1(n11391), .B2(n12065), .ZN(
        n1580) );
  AOI221_X1 U2948 ( .B1(n12135), .B2(n8546), .C1(n12132), .C2(n8090), .A(n1552), .ZN(n1547) );
  OAI22_X1 U2949 ( .A1(n11136), .A2(n12129), .B1(n11392), .B2(n12126), .ZN(
        n1552) );
  AOI221_X1 U2950 ( .B1(n12159), .B2(n8394), .C1(n12156), .C2(n7938), .A(n1550), .ZN(n1549) );
  OAI22_X1 U2951 ( .A1(n11137), .A2(n12153), .B1(n11393), .B2(n12150), .ZN(
        n1550) );
  AOI221_X1 U2952 ( .B1(n12147), .B2(n8444), .C1(n12144), .C2(n7988), .A(n1551), .ZN(n1548) );
  OAI22_X1 U2953 ( .A1(n11138), .A2(n12141), .B1(n11394), .B2(n12138), .ZN(
        n1551) );
  AOI221_X1 U2954 ( .B1(n12123), .B2(n8547), .C1(n12120), .C2(n8091), .A(n1553), .ZN(n1546) );
  OAI22_X1 U2955 ( .A1(n11139), .A2(n12117), .B1(n11395), .B2(n12114), .ZN(
        n1553) );
  AOI221_X1 U2956 ( .B1(n12075), .B2(n8507), .C1(n12072), .C2(n8051), .A(n1561), .ZN(n1554) );
  OAI22_X1 U2957 ( .A1(n11140), .A2(n12069), .B1(n11396), .B2(n12066), .ZN(
        n1561) );
  AOI221_X1 U2958 ( .B1(n12135), .B2(n8548), .C1(n12132), .C2(n8092), .A(n1533), .ZN(n1528) );
  OAI22_X1 U2959 ( .A1(n11141), .A2(n12129), .B1(n11397), .B2(n12126), .ZN(
        n1533) );
  AOI221_X1 U2960 ( .B1(n12159), .B2(n8396), .C1(n12156), .C2(n7940), .A(n1531), .ZN(n1530) );
  OAI22_X1 U2961 ( .A1(n11142), .A2(n12153), .B1(n11398), .B2(n12150), .ZN(
        n1531) );
  AOI221_X1 U2962 ( .B1(n12147), .B2(n8446), .C1(n12144), .C2(n7990), .A(n1532), .ZN(n1529) );
  OAI22_X1 U2963 ( .A1(n11143), .A2(n12141), .B1(n11399), .B2(n12138), .ZN(
        n1532) );
  AOI221_X1 U2964 ( .B1(n12123), .B2(n8549), .C1(n12120), .C2(n8093), .A(n1534), .ZN(n1527) );
  OAI22_X1 U2965 ( .A1(n11144), .A2(n12117), .B1(n11400), .B2(n12114), .ZN(
        n1534) );
  AOI221_X1 U2966 ( .B1(n12075), .B2(n8508), .C1(n12072), .C2(n8052), .A(n1542), .ZN(n1535) );
  OAI22_X1 U2967 ( .A1(n11145), .A2(n12069), .B1(n11401), .B2(n12066), .ZN(
        n1542) );
  AOI221_X1 U2968 ( .B1(n12135), .B2(n8550), .C1(n12132), .C2(n8094), .A(n1514), .ZN(n1509) );
  OAI22_X1 U2969 ( .A1(n11146), .A2(n12129), .B1(n11402), .B2(n12126), .ZN(
        n1514) );
  AOI221_X1 U2970 ( .B1(n12159), .B2(n8398), .C1(n12156), .C2(n7942), .A(n1512), .ZN(n1511) );
  OAI22_X1 U2971 ( .A1(n11147), .A2(n12153), .B1(n11403), .B2(n12150), .ZN(
        n1512) );
  AOI221_X1 U2972 ( .B1(n12147), .B2(n8448), .C1(n12144), .C2(n7992), .A(n1513), .ZN(n1510) );
  OAI22_X1 U2973 ( .A1(n11148), .A2(n12141), .B1(n11404), .B2(n12138), .ZN(
        n1513) );
  AOI221_X1 U2974 ( .B1(n12123), .B2(n8551), .C1(n12120), .C2(n8095), .A(n1515), .ZN(n1508) );
  OAI22_X1 U2975 ( .A1(n11149), .A2(n12117), .B1(n11405), .B2(n12114), .ZN(
        n1515) );
  AOI221_X1 U2976 ( .B1(n12075), .B2(n8509), .C1(n12072), .C2(n8053), .A(n1523), .ZN(n1516) );
  OAI22_X1 U2977 ( .A1(n11150), .A2(n12069), .B1(n11406), .B2(n12066), .ZN(
        n1523) );
  AOI221_X1 U2978 ( .B1(n12135), .B2(n8552), .C1(n12132), .C2(n8096), .A(n1495), .ZN(n1490) );
  OAI22_X1 U2979 ( .A1(n11151), .A2(n12129), .B1(n11407), .B2(n12126), .ZN(
        n1495) );
  AOI221_X1 U2980 ( .B1(n12159), .B2(n8400), .C1(n12156), .C2(n7944), .A(n1493), .ZN(n1492) );
  OAI22_X1 U2981 ( .A1(n11152), .A2(n12153), .B1(n11408), .B2(n12150), .ZN(
        n1493) );
  AOI221_X1 U2982 ( .B1(n12147), .B2(n8450), .C1(n12144), .C2(n7994), .A(n1494), .ZN(n1491) );
  OAI22_X1 U2983 ( .A1(n11153), .A2(n12141), .B1(n11409), .B2(n12138), .ZN(
        n1494) );
  AOI221_X1 U2984 ( .B1(n12123), .B2(n8553), .C1(n12120), .C2(n8097), .A(n1496), .ZN(n1489) );
  OAI22_X1 U2985 ( .A1(n11154), .A2(n12117), .B1(n11410), .B2(n12114), .ZN(
        n1496) );
  AOI221_X1 U2986 ( .B1(n12075), .B2(n8510), .C1(n12072), .C2(n8054), .A(n1504), .ZN(n1497) );
  OAI22_X1 U2987 ( .A1(n11155), .A2(n12069), .B1(n11411), .B2(n12066), .ZN(
        n1504) );
  AOI221_X1 U2988 ( .B1(n12135), .B2(n8554), .C1(n12132), .C2(n8098), .A(n1476), .ZN(n1471) );
  OAI22_X1 U2989 ( .A1(n11156), .A2(n12129), .B1(n11412), .B2(n12126), .ZN(
        n1476) );
  AOI221_X1 U2990 ( .B1(n12159), .B2(n8402), .C1(n12156), .C2(n7946), .A(n1474), .ZN(n1473) );
  OAI22_X1 U2991 ( .A1(n11157), .A2(n12153), .B1(n11413), .B2(n12150), .ZN(
        n1474) );
  AOI221_X1 U2992 ( .B1(n12147), .B2(n8452), .C1(n12144), .C2(n7996), .A(n1475), .ZN(n1472) );
  OAI22_X1 U2993 ( .A1(n11158), .A2(n12141), .B1(n11414), .B2(n12138), .ZN(
        n1475) );
  AOI221_X1 U2994 ( .B1(n12123), .B2(n8555), .C1(n12120), .C2(n8099), .A(n1477), .ZN(n1470) );
  OAI22_X1 U2995 ( .A1(n11159), .A2(n12117), .B1(n11415), .B2(n12114), .ZN(
        n1477) );
  AOI221_X1 U2996 ( .B1(n12075), .B2(n8511), .C1(n12072), .C2(n8055), .A(n1485), .ZN(n1478) );
  OAI22_X1 U2997 ( .A1(n11160), .A2(n12069), .B1(n11416), .B2(n12066), .ZN(
        n1485) );
  AOI221_X1 U2998 ( .B1(n12135), .B2(n8556), .C1(n12132), .C2(n8100), .A(n1457), .ZN(n1452) );
  OAI22_X1 U2999 ( .A1(n11161), .A2(n12129), .B1(n11417), .B2(n12126), .ZN(
        n1457) );
  AOI221_X1 U3000 ( .B1(n12159), .B2(n8404), .C1(n12156), .C2(n7948), .A(n1455), .ZN(n1454) );
  OAI22_X1 U3001 ( .A1(n11162), .A2(n12153), .B1(n11418), .B2(n12150), .ZN(
        n1455) );
  AOI221_X1 U3002 ( .B1(n12147), .B2(n8454), .C1(n12144), .C2(n7998), .A(n1456), .ZN(n1453) );
  OAI22_X1 U3003 ( .A1(n11163), .A2(n12141), .B1(n11419), .B2(n12138), .ZN(
        n1456) );
  AOI221_X1 U3004 ( .B1(n12123), .B2(n8557), .C1(n12120), .C2(n8101), .A(n1458), .ZN(n1451) );
  OAI22_X1 U3005 ( .A1(n11164), .A2(n12117), .B1(n11420), .B2(n12114), .ZN(
        n1458) );
  AOI221_X1 U3006 ( .B1(n12075), .B2(n8512), .C1(n12072), .C2(n8056), .A(n1466), .ZN(n1459) );
  OAI22_X1 U3007 ( .A1(n11165), .A2(n12069), .B1(n11421), .B2(n12066), .ZN(
        n1466) );
  AOI221_X1 U3008 ( .B1(n12135), .B2(n8558), .C1(n12132), .C2(n8102), .A(n1438), .ZN(n1433) );
  OAI22_X1 U3009 ( .A1(n11166), .A2(n12129), .B1(n11422), .B2(n12126), .ZN(
        n1438) );
  AOI221_X1 U3010 ( .B1(n12159), .B2(n8406), .C1(n12156), .C2(n7950), .A(n1436), .ZN(n1435) );
  OAI22_X1 U3011 ( .A1(n11167), .A2(n12153), .B1(n11423), .B2(n12150), .ZN(
        n1436) );
  AOI221_X1 U3012 ( .B1(n12147), .B2(n8456), .C1(n12144), .C2(n8000), .A(n1437), .ZN(n1434) );
  OAI22_X1 U3013 ( .A1(n11168), .A2(n12141), .B1(n11424), .B2(n12138), .ZN(
        n1437) );
  AOI221_X1 U3014 ( .B1(n12123), .B2(n8559), .C1(n12120), .C2(n8103), .A(n1439), .ZN(n1432) );
  OAI22_X1 U3015 ( .A1(n11169), .A2(n12117), .B1(n11425), .B2(n12114), .ZN(
        n1439) );
  AOI221_X1 U3016 ( .B1(n12075), .B2(n8513), .C1(n12072), .C2(n8057), .A(n1447), .ZN(n1440) );
  OAI22_X1 U3017 ( .A1(n11170), .A2(n12069), .B1(n11426), .B2(n12066), .ZN(
        n1447) );
  AOI221_X1 U3018 ( .B1(n12135), .B2(n8560), .C1(n12132), .C2(n8104), .A(n1419), .ZN(n1414) );
  OAI22_X1 U3019 ( .A1(n11171), .A2(n12129), .B1(n11427), .B2(n12126), .ZN(
        n1419) );
  AOI221_X1 U3020 ( .B1(n12159), .B2(n8408), .C1(n12156), .C2(n7952), .A(n1417), .ZN(n1416) );
  OAI22_X1 U3021 ( .A1(n11172), .A2(n12153), .B1(n11428), .B2(n12150), .ZN(
        n1417) );
  AOI221_X1 U3022 ( .B1(n12147), .B2(n8458), .C1(n12144), .C2(n8002), .A(n1418), .ZN(n1415) );
  OAI22_X1 U3023 ( .A1(n11173), .A2(n12141), .B1(n11429), .B2(n12138), .ZN(
        n1418) );
  AOI221_X1 U3024 ( .B1(n12123), .B2(n8561), .C1(n12120), .C2(n8105), .A(n1420), .ZN(n1413) );
  OAI22_X1 U3025 ( .A1(n11174), .A2(n12117), .B1(n11430), .B2(n12114), .ZN(
        n1420) );
  AOI221_X1 U3026 ( .B1(n12075), .B2(n8514), .C1(n12072), .C2(n8058), .A(n1428), .ZN(n1421) );
  OAI22_X1 U3027 ( .A1(n11175), .A2(n12069), .B1(n11431), .B2(n12066), .ZN(
        n1428) );
  AOI221_X1 U3028 ( .B1(n12135), .B2(n11519), .C1(n12132), .C2(n8106), .A(
        n1400), .ZN(n1395) );
  OAI22_X1 U3029 ( .A1(n11176), .A2(n12129), .B1(n11432), .B2(n12126), .ZN(
        n1400) );
  AOI221_X1 U3030 ( .B1(n12159), .B2(n11520), .C1(n12156), .C2(n7954), .A(
        n1398), .ZN(n1397) );
  OAI22_X1 U3031 ( .A1(n11177), .A2(n12153), .B1(n11433), .B2(n12150), .ZN(
        n1398) );
  AOI221_X1 U3032 ( .B1(n12123), .B2(n11521), .C1(n12120), .C2(n8107), .A(
        n1401), .ZN(n1394) );
  OAI22_X1 U3033 ( .A1(n11178), .A2(n12117), .B1(n11434), .B2(n12114), .ZN(
        n1401) );
  AOI221_X1 U3034 ( .B1(n12075), .B2(n8515), .C1(n12072), .C2(n8059), .A(n1409), .ZN(n1402) );
  OAI22_X1 U3035 ( .A1(n11179), .A2(n12069), .B1(n11435), .B2(n12066), .ZN(
        n1409) );
  AOI221_X1 U3036 ( .B1(n12135), .B2(n11522), .C1(n12132), .C2(n8108), .A(
        n1381), .ZN(n1376) );
  OAI22_X1 U3037 ( .A1(n11180), .A2(n12129), .B1(n11436), .B2(n12126), .ZN(
        n1381) );
  AOI221_X1 U3038 ( .B1(n12159), .B2(n11523), .C1(n12156), .C2(n7956), .A(
        n1379), .ZN(n1378) );
  OAI22_X1 U3039 ( .A1(n11181), .A2(n12153), .B1(n11437), .B2(n12150), .ZN(
        n1379) );
  AOI221_X1 U3040 ( .B1(n12123), .B2(n8565), .C1(n12120), .C2(n8109), .A(n1382), .ZN(n1375) );
  OAI22_X1 U3041 ( .A1(n11182), .A2(n12117), .B1(n11438), .B2(n12114), .ZN(
        n1382) );
  AOI221_X1 U3042 ( .B1(n12075), .B2(n8516), .C1(n12072), .C2(n8060), .A(n1390), .ZN(n1383) );
  OAI22_X1 U3043 ( .A1(n11183), .A2(n12069), .B1(n11439), .B2(n12066), .ZN(
        n1390) );
  AOI221_X1 U3044 ( .B1(n12136), .B2(n11524), .C1(n12133), .C2(n8110), .A(
        n1362), .ZN(n1357) );
  OAI22_X1 U3045 ( .A1(n11184), .A2(n12129), .B1(n11440), .B2(n12126), .ZN(
        n1362) );
  AOI221_X1 U3046 ( .B1(n12160), .B2(n11525), .C1(n12157), .C2(n7958), .A(
        n1360), .ZN(n1359) );
  OAI22_X1 U3047 ( .A1(n11185), .A2(n12153), .B1(n11441), .B2(n12150), .ZN(
        n1360) );
  AOI221_X1 U3048 ( .B1(n12124), .B2(n8567), .C1(n12121), .C2(n8111), .A(n1363), .ZN(n1356) );
  OAI22_X1 U3049 ( .A1(n11186), .A2(n12117), .B1(n11442), .B2(n12114), .ZN(
        n1363) );
  AOI221_X1 U3050 ( .B1(n12076), .B2(n8517), .C1(n12073), .C2(n8061), .A(n1371), .ZN(n1364) );
  OAI22_X1 U3051 ( .A1(n11187), .A2(n12069), .B1(n11443), .B2(n12066), .ZN(
        n1371) );
  AOI221_X1 U3052 ( .B1(n12136), .B2(n11526), .C1(n12133), .C2(n8112), .A(
        n1343), .ZN(n1338) );
  OAI22_X1 U3053 ( .A1(n11188), .A2(n12129), .B1(n11444), .B2(n12126), .ZN(
        n1343) );
  AOI221_X1 U3054 ( .B1(n12160), .B2(n11527), .C1(n12157), .C2(n7960), .A(
        n1341), .ZN(n1340) );
  OAI22_X1 U3055 ( .A1(n11189), .A2(n12153), .B1(n11445), .B2(n12150), .ZN(
        n1341) );
  AOI221_X1 U3056 ( .B1(n12124), .B2(n8569), .C1(n12121), .C2(n8113), .A(n1344), .ZN(n1337) );
  OAI22_X1 U3057 ( .A1(n11190), .A2(n12117), .B1(n11446), .B2(n12114), .ZN(
        n1344) );
  AOI221_X1 U3058 ( .B1(n12076), .B2(n8518), .C1(n12073), .C2(n8062), .A(n1352), .ZN(n1345) );
  OAI22_X1 U3059 ( .A1(n11191), .A2(n12069), .B1(n11447), .B2(n12066), .ZN(
        n1352) );
  NOR3_X1 U3060 ( .A1(n1808), .A2(n12567), .A3(n1809), .ZN(n1807) );
  XNOR2_X1 U3061 ( .A(n12564), .B(ADD_RD1[0]), .ZN(n1808) );
  XNOR2_X1 U3062 ( .A(n12566), .B(ADD_RD1[4]), .ZN(n1809) );
  AND2_X1 U3063 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[1]), .ZN(n1783) );
  NAND2_X1 U3064 ( .A1(n12559), .A2(n2466), .ZN(n1811) );
  NAND2_X1 U3065 ( .A1(RD2), .A2(EN), .ZN(n2466) );
  NAND2_X1 U3066 ( .A1(n12559), .A2(n1803), .ZN(n1148) );
  NAND2_X1 U3067 ( .A1(RD1), .A2(EN), .ZN(n1803) );
  INV_X1 U3068 ( .A(ADD_WR[0]), .ZN(n12564) );
  INV_X1 U3069 ( .A(ADD_RD1[3]), .ZN(n12572) );
  INV_X1 U3070 ( .A(ADD_RD1[0]), .ZN(n12571) );
  INV_X1 U3071 ( .A(ADD_WR[1]), .ZN(n12563) );
  INV_X1 U3072 ( .A(ADD_WR[2]), .ZN(n12565) );
  NAND4_X1 U3073 ( .A1(n1804), .A2(n1805), .A3(n1806), .A4(n1807), .ZN(n1774)
         );
  XNOR2_X1 U3074 ( .A(ADD_RD1[1]), .B(ADD_WR[1]), .ZN(n1804) );
  XNOR2_X1 U3075 ( .A(ADD_WR[3]), .B(ADD_RD1[3]), .ZN(n1805) );
  XNOR2_X1 U3076 ( .A(ADD_RD1[2]), .B(ADD_WR[2]), .ZN(n1806) );
  AND3_X1 U3077 ( .A1(ADD_RD1[4]), .A2(n12572), .A3(ADD_RD1[0]), .ZN(n1789) );
  AND3_X1 U3078 ( .A1(ADD_RD1[4]), .A2(n12571), .A3(ADD_RD1[3]), .ZN(n1780) );
  AND3_X1 U3079 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(ADD_RD1[3]), .ZN(n1782) );
  AND3_X1 U3080 ( .A1(n12571), .A2(n12572), .A3(ADD_RD1[4]), .ZN(n1788) );
  INV_X1 U3081 ( .A(ADD_RD1[1]), .ZN(n12573) );
  INV_X1 U3082 ( .A(WR), .ZN(n12567) );
  NAND2_X1 U3083 ( .A1(DATAIN[24]), .A2(n12554), .ZN(n1096) );
  NAND2_X1 U3084 ( .A1(DATAIN[3]), .A2(n12556), .ZN(n1075) );
  NAND2_X1 U3085 ( .A1(DATAIN[9]), .A2(n12555), .ZN(n1081) );
  NAND2_X1 U3086 ( .A1(DATAIN[10]), .A2(n12555), .ZN(n1082) );
  NAND2_X1 U3087 ( .A1(DATAIN[17]), .A2(n12555), .ZN(n1089) );
  NAND2_X1 U3088 ( .A1(DATAIN[20]), .A2(n12554), .ZN(n1092) );
  NAND2_X1 U3089 ( .A1(DATAIN[0]), .A2(n12555), .ZN(n1071) );
  NAND2_X1 U3090 ( .A1(DATAIN[1]), .A2(n12556), .ZN(n1073) );
  INV_X1 U3091 ( .A(n12177), .ZN(n12170) );
  INV_X1 U3092 ( .A(n12195), .ZN(n12188) );
  CLKBUF_X1 U3093 ( .A(RST), .Z(n12554) );
  CLKBUF_X1 U3094 ( .A(RST), .Z(n12555) );
  CLKBUF_X1 U3095 ( .A(RST), .Z(n12556) );
  CLKBUF_X1 U3096 ( .A(RST), .Z(n12557) );
  CLKBUF_X1 U3097 ( .A(RST), .Z(n12558) );
  CLKBUF_X1 U3098 ( .A(RST), .Z(n12559) );
endmodule


module REGISTER_GENERIC_WIDTH32_10 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296;

  DFF_X1 \DOUT_reg[31]  ( .D(n68), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[30]  ( .D(n69), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[29]  ( .D(n70), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[28]  ( .D(n71), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[27]  ( .D(n72), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n73), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[25]  ( .D(n74), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[24]  ( .D(n75), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[22]  ( .D(n77), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[21]  ( .D(n78), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[20]  ( .D(n79), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n80), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n81), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n83), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n84), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n89), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n90), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n91), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n92), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n93), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n94), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n95), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n96), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n97), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n98), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n260) );
  BUF_X1 U4 ( .A(n35), .Z(n259) );
  BUF_X1 U5 ( .A(n35), .Z(n258) );
  NAND2_X1 U6 ( .A1(RST), .A2(n261), .ZN(n35) );
  BUF_X1 U7 ( .A(n34), .Z(n263) );
  BUF_X1 U8 ( .A(n34), .Z(n261) );
  BUF_X1 U9 ( .A(n34), .Z(n262) );
  OAI22_X1 U10 ( .A1(n36), .A2(n263), .B1(n260), .B2(n295), .ZN(n99) );
  INV_X1 U11 ( .A(DIN[0]), .ZN(n295) );
  OAI22_X1 U12 ( .A1(n37), .A2(n263), .B1(n260), .B2(n294), .ZN(n98) );
  INV_X1 U13 ( .A(DIN[1]), .ZN(n294) );
  OAI22_X1 U14 ( .A1(n38), .A2(n263), .B1(n260), .B2(n293), .ZN(n97) );
  INV_X1 U15 ( .A(DIN[2]), .ZN(n293) );
  OAI22_X1 U16 ( .A1(n39), .A2(n263), .B1(n260), .B2(n292), .ZN(n96) );
  INV_X1 U17 ( .A(DIN[3]), .ZN(n292) );
  OAI22_X1 U18 ( .A1(n40), .A2(n263), .B1(n260), .B2(n291), .ZN(n95) );
  INV_X1 U19 ( .A(DIN[4]), .ZN(n291) );
  OAI22_X1 U20 ( .A1(n41), .A2(n263), .B1(n260), .B2(n290), .ZN(n94) );
  INV_X1 U21 ( .A(DIN[5]), .ZN(n290) );
  OAI22_X1 U22 ( .A1(n42), .A2(n263), .B1(n260), .B2(n289), .ZN(n93) );
  INV_X1 U23 ( .A(DIN[6]), .ZN(n289) );
  OAI22_X1 U24 ( .A1(n43), .A2(n263), .B1(n260), .B2(n288), .ZN(n92) );
  INV_X1 U25 ( .A(DIN[7]), .ZN(n288) );
  OAI22_X1 U26 ( .A1(n44), .A2(n263), .B1(n260), .B2(n287), .ZN(n91) );
  INV_X1 U27 ( .A(DIN[8]), .ZN(n287) );
  OAI22_X1 U28 ( .A1(n45), .A2(n262), .B1(n260), .B2(n286), .ZN(n90) );
  INV_X1 U29 ( .A(DIN[9]), .ZN(n286) );
  OAI22_X1 U30 ( .A1(n46), .A2(n262), .B1(n259), .B2(n285), .ZN(n89) );
  INV_X1 U31 ( .A(DIN[10]), .ZN(n285) );
  OAI22_X1 U32 ( .A1(n47), .A2(n262), .B1(n259), .B2(n284), .ZN(n88) );
  INV_X1 U33 ( .A(DIN[11]), .ZN(n284) );
  OAI22_X1 U34 ( .A1(n48), .A2(n262), .B1(n259), .B2(n283), .ZN(n87) );
  INV_X1 U35 ( .A(DIN[12]), .ZN(n283) );
  OAI22_X1 U36 ( .A1(n49), .A2(n262), .B1(n259), .B2(n282), .ZN(n86) );
  INV_X1 U37 ( .A(DIN[13]), .ZN(n282) );
  OAI22_X1 U38 ( .A1(n50), .A2(n262), .B1(n259), .B2(n281), .ZN(n85) );
  INV_X1 U39 ( .A(DIN[14]), .ZN(n281) );
  OAI22_X1 U40 ( .A1(n51), .A2(n262), .B1(n259), .B2(n280), .ZN(n84) );
  INV_X1 U41 ( .A(DIN[15]), .ZN(n280) );
  OAI22_X1 U42 ( .A1(n52), .A2(n262), .B1(n259), .B2(n279), .ZN(n83) );
  INV_X1 U43 ( .A(DIN[16]), .ZN(n279) );
  OAI22_X1 U44 ( .A1(n53), .A2(n262), .B1(n259), .B2(n278), .ZN(n82) );
  INV_X1 U45 ( .A(DIN[17]), .ZN(n278) );
  OAI22_X1 U46 ( .A1(n54), .A2(n262), .B1(n259), .B2(n277), .ZN(n81) );
  INV_X1 U47 ( .A(DIN[18]), .ZN(n277) );
  OAI22_X1 U48 ( .A1(n55), .A2(n262), .B1(n259), .B2(n276), .ZN(n80) );
  INV_X1 U49 ( .A(DIN[19]), .ZN(n276) );
  OAI22_X1 U50 ( .A1(n56), .A2(n262), .B1(n259), .B2(n275), .ZN(n79) );
  INV_X1 U51 ( .A(DIN[20]), .ZN(n275) );
  OAI22_X1 U52 ( .A1(n57), .A2(n261), .B1(n258), .B2(n274), .ZN(n78) );
  INV_X1 U53 ( .A(DIN[21]), .ZN(n274) );
  OAI22_X1 U54 ( .A1(n58), .A2(n261), .B1(n258), .B2(n273), .ZN(n77) );
  INV_X1 U55 ( .A(DIN[22]), .ZN(n273) );
  OAI22_X1 U56 ( .A1(n59), .A2(n261), .B1(n258), .B2(n272), .ZN(n76) );
  INV_X1 U57 ( .A(DIN[23]), .ZN(n272) );
  OAI22_X1 U58 ( .A1(n60), .A2(n261), .B1(n258), .B2(n271), .ZN(n75) );
  INV_X1 U59 ( .A(DIN[24]), .ZN(n271) );
  OAI22_X1 U60 ( .A1(n61), .A2(n261), .B1(n258), .B2(n270), .ZN(n74) );
  INV_X1 U61 ( .A(DIN[25]), .ZN(n270) );
  OAI22_X1 U62 ( .A1(n62), .A2(n261), .B1(n258), .B2(n269), .ZN(n73) );
  INV_X1 U63 ( .A(DIN[26]), .ZN(n269) );
  OAI22_X1 U64 ( .A1(n63), .A2(n261), .B1(n258), .B2(n268), .ZN(n72) );
  INV_X1 U65 ( .A(DIN[27]), .ZN(n268) );
  OAI22_X1 U66 ( .A1(n64), .A2(n261), .B1(n258), .B2(n267), .ZN(n71) );
  INV_X1 U67 ( .A(DIN[28]), .ZN(n267) );
  OAI22_X1 U68 ( .A1(n65), .A2(n261), .B1(n258), .B2(n266), .ZN(n70) );
  INV_X1 U69 ( .A(DIN[29]), .ZN(n266) );
  OAI22_X1 U70 ( .A1(n66), .A2(n261), .B1(n258), .B2(n265), .ZN(n69) );
  INV_X1 U71 ( .A(DIN[30]), .ZN(n265) );
  OAI22_X1 U72 ( .A1(n67), .A2(n261), .B1(n258), .B2(n264), .ZN(n68) );
  INV_X1 U73 ( .A(DIN[31]), .ZN(n264) );
  NAND2_X1 U74 ( .A1(n296), .A2(RST), .ZN(n34) );
  INV_X1 U75 ( .A(EN), .ZN(n296) );
endmodule


module REGISTER_GENERIC_WIDTH32_9 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298;

  DFF_X1 \DOUT_reg[31]  ( .D(n68), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[30]  ( .D(n69), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[29]  ( .D(n70), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[28]  ( .D(n71), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[27]  ( .D(n72), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n73), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[25]  ( .D(n74), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[24]  ( .D(n75), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[22]  ( .D(n77), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[21]  ( .D(n78), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[20]  ( .D(n79), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n80), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n81), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n83), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n84), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n89), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n90), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n91), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n92), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n93), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n94), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n95), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n96), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n97), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n98), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n262) );
  BUF_X1 U4 ( .A(n35), .Z(n261) );
  BUF_X1 U5 ( .A(n35), .Z(n260) );
  NAND2_X1 U6 ( .A1(RST), .A2(n263), .ZN(n35) );
  BUF_X1 U7 ( .A(n34), .Z(n265) );
  BUF_X1 U8 ( .A(n34), .Z(n263) );
  BUF_X1 U9 ( .A(n34), .Z(n264) );
  OAI22_X1 U10 ( .A1(n36), .A2(n265), .B1(n262), .B2(n297), .ZN(n99) );
  INV_X1 U11 ( .A(DIN[0]), .ZN(n297) );
  OAI22_X1 U12 ( .A1(n37), .A2(n265), .B1(n262), .B2(n296), .ZN(n98) );
  INV_X1 U13 ( .A(DIN[1]), .ZN(n296) );
  OAI22_X1 U14 ( .A1(n38), .A2(n265), .B1(n262), .B2(n295), .ZN(n97) );
  INV_X1 U15 ( .A(DIN[2]), .ZN(n295) );
  OAI22_X1 U16 ( .A1(n39), .A2(n265), .B1(n262), .B2(n294), .ZN(n96) );
  INV_X1 U17 ( .A(DIN[3]), .ZN(n294) );
  OAI22_X1 U18 ( .A1(n40), .A2(n265), .B1(n262), .B2(n293), .ZN(n95) );
  INV_X1 U19 ( .A(DIN[4]), .ZN(n293) );
  OAI22_X1 U20 ( .A1(n41), .A2(n265), .B1(n262), .B2(n292), .ZN(n94) );
  INV_X1 U21 ( .A(DIN[5]), .ZN(n292) );
  OAI22_X1 U22 ( .A1(n42), .A2(n265), .B1(n262), .B2(n291), .ZN(n93) );
  INV_X1 U23 ( .A(DIN[6]), .ZN(n291) );
  OAI22_X1 U24 ( .A1(n43), .A2(n265), .B1(n262), .B2(n290), .ZN(n92) );
  INV_X1 U25 ( .A(DIN[7]), .ZN(n290) );
  OAI22_X1 U26 ( .A1(n44), .A2(n265), .B1(n262), .B2(n289), .ZN(n91) );
  INV_X1 U27 ( .A(DIN[8]), .ZN(n289) );
  OAI22_X1 U28 ( .A1(n45), .A2(n264), .B1(n262), .B2(n288), .ZN(n90) );
  INV_X1 U29 ( .A(DIN[9]), .ZN(n288) );
  OAI22_X1 U30 ( .A1(n46), .A2(n264), .B1(n261), .B2(n287), .ZN(n89) );
  INV_X1 U31 ( .A(DIN[10]), .ZN(n287) );
  OAI22_X1 U32 ( .A1(n47), .A2(n264), .B1(n261), .B2(n286), .ZN(n88) );
  INV_X1 U33 ( .A(DIN[11]), .ZN(n286) );
  OAI22_X1 U34 ( .A1(n48), .A2(n264), .B1(n261), .B2(n285), .ZN(n87) );
  INV_X1 U35 ( .A(DIN[12]), .ZN(n285) );
  OAI22_X1 U36 ( .A1(n49), .A2(n264), .B1(n261), .B2(n284), .ZN(n86) );
  INV_X1 U37 ( .A(DIN[13]), .ZN(n284) );
  OAI22_X1 U38 ( .A1(n50), .A2(n264), .B1(n261), .B2(n283), .ZN(n85) );
  INV_X1 U39 ( .A(DIN[14]), .ZN(n283) );
  OAI22_X1 U40 ( .A1(n51), .A2(n264), .B1(n261), .B2(n282), .ZN(n84) );
  INV_X1 U41 ( .A(DIN[15]), .ZN(n282) );
  OAI22_X1 U42 ( .A1(n52), .A2(n264), .B1(n261), .B2(n281), .ZN(n83) );
  INV_X1 U43 ( .A(DIN[16]), .ZN(n281) );
  OAI22_X1 U44 ( .A1(n53), .A2(n264), .B1(n261), .B2(n280), .ZN(n82) );
  INV_X1 U45 ( .A(DIN[17]), .ZN(n280) );
  OAI22_X1 U46 ( .A1(n54), .A2(n264), .B1(n261), .B2(n279), .ZN(n81) );
  INV_X1 U47 ( .A(DIN[18]), .ZN(n279) );
  OAI22_X1 U48 ( .A1(n55), .A2(n264), .B1(n261), .B2(n278), .ZN(n80) );
  INV_X1 U49 ( .A(DIN[19]), .ZN(n278) );
  OAI22_X1 U50 ( .A1(n56), .A2(n264), .B1(n261), .B2(n277), .ZN(n79) );
  INV_X1 U51 ( .A(DIN[20]), .ZN(n277) );
  OAI22_X1 U52 ( .A1(n57), .A2(n263), .B1(n260), .B2(n276), .ZN(n78) );
  INV_X1 U53 ( .A(DIN[21]), .ZN(n276) );
  OAI22_X1 U54 ( .A1(n58), .A2(n263), .B1(n260), .B2(n275), .ZN(n77) );
  INV_X1 U55 ( .A(DIN[22]), .ZN(n275) );
  OAI22_X1 U56 ( .A1(n59), .A2(n263), .B1(n260), .B2(n274), .ZN(n76) );
  INV_X1 U57 ( .A(DIN[23]), .ZN(n274) );
  OAI22_X1 U58 ( .A1(n60), .A2(n263), .B1(n260), .B2(n273), .ZN(n75) );
  INV_X1 U59 ( .A(DIN[24]), .ZN(n273) );
  OAI22_X1 U60 ( .A1(n61), .A2(n263), .B1(n260), .B2(n272), .ZN(n74) );
  INV_X1 U61 ( .A(DIN[25]), .ZN(n272) );
  OAI22_X1 U62 ( .A1(n62), .A2(n263), .B1(n260), .B2(n271), .ZN(n73) );
  INV_X1 U63 ( .A(DIN[26]), .ZN(n271) );
  OAI22_X1 U64 ( .A1(n63), .A2(n263), .B1(n260), .B2(n270), .ZN(n72) );
  INV_X1 U65 ( .A(DIN[27]), .ZN(n270) );
  OAI22_X1 U66 ( .A1(n64), .A2(n263), .B1(n260), .B2(n269), .ZN(n71) );
  INV_X1 U67 ( .A(DIN[28]), .ZN(n269) );
  OAI22_X1 U68 ( .A1(n65), .A2(n263), .B1(n260), .B2(n268), .ZN(n70) );
  INV_X1 U69 ( .A(DIN[29]), .ZN(n268) );
  OAI22_X1 U70 ( .A1(n66), .A2(n263), .B1(n260), .B2(n267), .ZN(n69) );
  INV_X1 U71 ( .A(DIN[30]), .ZN(n267) );
  OAI22_X1 U72 ( .A1(n67), .A2(n263), .B1(n260), .B2(n266), .ZN(n68) );
  INV_X1 U73 ( .A(DIN[31]), .ZN(n266) );
  NAND2_X1 U74 ( .A1(n298), .A2(RST), .ZN(n34) );
  INV_X1 U75 ( .A(EN), .ZN(n298) );
endmodule


module SIGN_EXTEND_WIDTH_IN16_WIDTH_OUT32_0 ( A, S, Y );
  input [15:0] A;
  output [31:0] Y;
  input S;
  wire   N0;
  assign Y[15] = A[15];
  assign Y[14] = A[14];
  assign Y[13] = A[13];
  assign Y[12] = A[12];
  assign Y[11] = A[11];
  assign Y[10] = A[10];
  assign Y[9] = A[9];
  assign Y[8] = A[8];
  assign Y[7] = A[7];
  assign Y[6] = A[6];
  assign Y[5] = A[5];
  assign Y[4] = A[4];
  assign Y[3] = A[3];
  assign Y[2] = A[2];
  assign Y[1] = A[1];
  assign Y[0] = A[0];
  assign Y[16] = N0;
  assign Y[17] = N0;
  assign Y[18] = N0;
  assign Y[19] = N0;
  assign Y[20] = N0;
  assign Y[21] = N0;
  assign Y[22] = N0;
  assign Y[23] = N0;
  assign Y[24] = N0;
  assign Y[25] = N0;
  assign Y[26] = N0;
  assign Y[27] = N0;
  assign Y[28] = N0;
  assign Y[29] = N0;
  assign Y[30] = N0;
  assign Y[31] = N0;

  AND2_X1 U1 ( .A1(S), .A2(A[15]), .ZN(N0) );
endmodule


module SIGN_EXTEND_WIDTH_IN26_WIDTH_OUT32 ( A, S, Y );
  input [25:0] A;
  output [31:0] Y;
  input S;
  wire   N0;
  assign Y[25] = A[25];
  assign Y[24] = A[24];
  assign Y[23] = A[23];
  assign Y[22] = A[22];
  assign Y[21] = A[21];
  assign Y[20] = A[20];
  assign Y[19] = A[19];
  assign Y[18] = A[18];
  assign Y[17] = A[17];
  assign Y[16] = A[16];
  assign Y[15] = A[15];
  assign Y[14] = A[14];
  assign Y[13] = A[13];
  assign Y[12] = A[12];
  assign Y[11] = A[11];
  assign Y[10] = A[10];
  assign Y[9] = A[9];
  assign Y[8] = A[8];
  assign Y[7] = A[7];
  assign Y[6] = A[6];
  assign Y[5] = A[5];
  assign Y[4] = A[4];
  assign Y[3] = A[3];
  assign Y[2] = A[2];
  assign Y[1] = A[1];
  assign Y[0] = A[0];
  assign Y[26] = N0;
  assign Y[27] = N0;
  assign Y[28] = N0;
  assign Y[29] = N0;
  assign Y[30] = N0;
  assign Y[31] = N0;

  AND2_X1 U1 ( .A1(S), .A2(A[25]), .ZN(N0) );
endmodule


module MUX21_GENERIC_NBIT32_6 ( S1, S0, SEL, Y );
  input [31:0] S1;
  input [31:0] S0;
  output [31:0] Y;
  input SEL;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262;

  INV_X1 U1 ( .A(n262), .ZN(n252) );
  INV_X1 U2 ( .A(n262), .ZN(n253) );
  BUF_X1 U3 ( .A(n251), .Z(n260) );
  BUF_X1 U4 ( .A(n250), .Z(n259) );
  BUF_X1 U5 ( .A(n250), .Z(n257) );
  BUF_X1 U6 ( .A(n249), .Z(n256) );
  BUF_X1 U7 ( .A(n250), .Z(n258) );
  BUF_X1 U8 ( .A(n249), .Z(n255) );
  BUF_X1 U9 ( .A(n249), .Z(n254) );
  BUF_X1 U10 ( .A(n251), .Z(n262) );
  BUF_X1 U11 ( .A(n251), .Z(n261) );
  INV_X1 U12 ( .A(n64), .ZN(Y[1]) );
  AOI22_X1 U13 ( .A1(S0[1]), .A2(n252), .B1(S1[1]), .B2(n261), .ZN(n64) );
  INV_X1 U14 ( .A(n63), .ZN(Y[2]) );
  AOI22_X1 U15 ( .A1(S0[2]), .A2(n252), .B1(S1[2]), .B2(n261), .ZN(n63) );
  INV_X1 U16 ( .A(n62), .ZN(Y[3]) );
  AOI22_X1 U17 ( .A1(S0[3]), .A2(n252), .B1(S1[3]), .B2(n260), .ZN(n62) );
  INV_X1 U18 ( .A(n61), .ZN(Y[4]) );
  AOI22_X1 U19 ( .A1(S0[4]), .A2(n252), .B1(S1[4]), .B2(n260), .ZN(n61) );
  INV_X1 U20 ( .A(n60), .ZN(Y[5]) );
  AOI22_X1 U21 ( .A1(S0[5]), .A2(n252), .B1(S1[5]), .B2(n260), .ZN(n60) );
  INV_X1 U22 ( .A(n59), .ZN(Y[6]) );
  AOI22_X1 U23 ( .A1(S0[6]), .A2(n252), .B1(S1[6]), .B2(n260), .ZN(n59) );
  INV_X1 U24 ( .A(n58), .ZN(Y[7]) );
  AOI22_X1 U25 ( .A1(S0[7]), .A2(n252), .B1(S1[7]), .B2(n259), .ZN(n58) );
  INV_X1 U26 ( .A(n57), .ZN(Y[8]) );
  AOI22_X1 U27 ( .A1(S0[8]), .A2(n252), .B1(S1[8]), .B2(n259), .ZN(n57) );
  INV_X1 U28 ( .A(n56), .ZN(Y[9]) );
  AOI22_X1 U29 ( .A1(S0[9]), .A2(n252), .B1(S1[9]), .B2(n259), .ZN(n56) );
  INV_X1 U30 ( .A(n55), .ZN(Y[10]) );
  AOI22_X1 U31 ( .A1(S0[10]), .A2(n252), .B1(S1[10]), .B2(n259), .ZN(n55) );
  INV_X1 U32 ( .A(n65), .ZN(Y[0]) );
  AOI22_X1 U33 ( .A1(S0[0]), .A2(n252), .B1(S1[0]), .B2(n261), .ZN(n65) );
  INV_X1 U34 ( .A(n54), .ZN(Y[11]) );
  AOI22_X1 U35 ( .A1(S0[11]), .A2(n252), .B1(S1[11]), .B2(n258), .ZN(n54) );
  INV_X1 U36 ( .A(n53), .ZN(Y[12]) );
  AOI22_X1 U37 ( .A1(S0[12]), .A2(n253), .B1(S1[12]), .B2(n258), .ZN(n53) );
  INV_X1 U38 ( .A(n52), .ZN(Y[13]) );
  AOI22_X1 U39 ( .A1(S0[13]), .A2(n253), .B1(S1[13]), .B2(n258), .ZN(n52) );
  INV_X1 U40 ( .A(n51), .ZN(Y[14]) );
  AOI22_X1 U41 ( .A1(S0[14]), .A2(n253), .B1(S1[14]), .B2(n257), .ZN(n51) );
  INV_X1 U42 ( .A(n50), .ZN(Y[15]) );
  AOI22_X1 U43 ( .A1(S0[15]), .A2(n253), .B1(S1[15]), .B2(n257), .ZN(n50) );
  INV_X1 U44 ( .A(n49), .ZN(Y[16]) );
  AOI22_X1 U45 ( .A1(S0[16]), .A2(n253), .B1(S1[16]), .B2(n257), .ZN(n49) );
  INV_X1 U46 ( .A(n48), .ZN(Y[17]) );
  AOI22_X1 U47 ( .A1(S0[17]), .A2(n253), .B1(S1[17]), .B2(n257), .ZN(n48) );
  INV_X1 U48 ( .A(n47), .ZN(Y[18]) );
  AOI22_X1 U49 ( .A1(S0[18]), .A2(n253), .B1(S1[18]), .B2(n256), .ZN(n47) );
  INV_X1 U50 ( .A(n46), .ZN(Y[19]) );
  AOI22_X1 U51 ( .A1(S0[19]), .A2(n253), .B1(S1[19]), .B2(n256), .ZN(n46) );
  INV_X1 U52 ( .A(n45), .ZN(Y[20]) );
  AOI22_X1 U53 ( .A1(S0[20]), .A2(n253), .B1(S1[20]), .B2(n256), .ZN(n45) );
  INV_X1 U54 ( .A(n44), .ZN(Y[21]) );
  AOI22_X1 U55 ( .A1(S0[21]), .A2(n253), .B1(S1[21]), .B2(n256), .ZN(n44) );
  INV_X1 U56 ( .A(n43), .ZN(Y[22]) );
  AOI22_X1 U57 ( .A1(S0[22]), .A2(n253), .B1(S1[22]), .B2(n255), .ZN(n43) );
  INV_X1 U58 ( .A(n42), .ZN(Y[23]) );
  AOI22_X1 U59 ( .A1(S0[23]), .A2(n253), .B1(S1[23]), .B2(n258), .ZN(n42) );
  INV_X1 U60 ( .A(n41), .ZN(Y[24]) );
  AOI22_X1 U61 ( .A1(S0[24]), .A2(n253), .B1(S1[24]), .B2(n255), .ZN(n41) );
  INV_X1 U62 ( .A(n40), .ZN(Y[25]) );
  AOI22_X1 U63 ( .A1(S0[25]), .A2(n252), .B1(S1[25]), .B2(n255), .ZN(n40) );
  INV_X1 U64 ( .A(n39), .ZN(Y[26]) );
  AOI22_X1 U65 ( .A1(S0[26]), .A2(n253), .B1(S1[26]), .B2(n255), .ZN(n39) );
  INV_X1 U66 ( .A(n38), .ZN(Y[27]) );
  AOI22_X1 U67 ( .A1(S0[27]), .A2(n252), .B1(S1[27]), .B2(n254), .ZN(n38) );
  INV_X1 U68 ( .A(n37), .ZN(Y[28]) );
  AOI22_X1 U69 ( .A1(S0[28]), .A2(n253), .B1(S1[28]), .B2(n254), .ZN(n37) );
  INV_X1 U70 ( .A(n36), .ZN(Y[29]) );
  AOI22_X1 U71 ( .A1(S0[29]), .A2(n252), .B1(S1[29]), .B2(n254), .ZN(n36) );
  INV_X1 U72 ( .A(n35), .ZN(Y[30]) );
  AOI22_X1 U73 ( .A1(S0[30]), .A2(n253), .B1(S1[30]), .B2(n254), .ZN(n35) );
  BUF_X1 U74 ( .A(SEL), .Z(n251) );
  BUF_X1 U75 ( .A(SEL), .Z(n250) );
  BUF_X1 U76 ( .A(SEL), .Z(n249) );
  INV_X1 U77 ( .A(n34), .ZN(Y[31]) );
  AOI22_X1 U78 ( .A1(S0[31]), .A2(n252), .B1(n261), .B2(S1[31]), .ZN(n34) );
endmodule


module REGISTER_GENERIC_WIDTH32_8 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294;

  DFF_X1 \DOUT_reg[31]  ( .D(n84), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[30]  ( .D(n83), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[29]  ( .D(n82), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[28]  ( .D(n81), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[27]  ( .D(n80), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n79), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[25]  ( .D(n78), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[24]  ( .D(n77), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[22]  ( .D(n75), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[21]  ( .D(n74), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[20]  ( .D(n73), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n72), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n71), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n70), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n69), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n68), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n90), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n99), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n98), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n97), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n96), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n95), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n94), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n93), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n92), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n91), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n89), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n258) );
  BUF_X1 U4 ( .A(n35), .Z(n256) );
  BUF_X1 U5 ( .A(n35), .Z(n257) );
  NAND2_X1 U6 ( .A1(RST), .A2(n259), .ZN(n35) );
  BUF_X1 U7 ( .A(n34), .Z(n261) );
  BUF_X1 U8 ( .A(n34), .Z(n259) );
  BUF_X1 U9 ( .A(n34), .Z(n260) );
  OAI22_X1 U10 ( .A1(n37), .A2(n261), .B1(n258), .B2(n293), .ZN(n91) );
  INV_X1 U11 ( .A(DIN[1]), .ZN(n293) );
  OAI22_X1 U12 ( .A1(n38), .A2(n261), .B1(n258), .B2(n292), .ZN(n92) );
  INV_X1 U13 ( .A(DIN[2]), .ZN(n292) );
  OAI22_X1 U14 ( .A1(n39), .A2(n261), .B1(n258), .B2(n291), .ZN(n93) );
  INV_X1 U15 ( .A(DIN[3]), .ZN(n291) );
  OAI22_X1 U16 ( .A1(n40), .A2(n261), .B1(n258), .B2(n290), .ZN(n94) );
  INV_X1 U17 ( .A(DIN[4]), .ZN(n290) );
  OAI22_X1 U18 ( .A1(n41), .A2(n261), .B1(n258), .B2(n289), .ZN(n95) );
  INV_X1 U19 ( .A(DIN[5]), .ZN(n289) );
  OAI22_X1 U20 ( .A1(n42), .A2(n261), .B1(n258), .B2(n288), .ZN(n96) );
  INV_X1 U21 ( .A(DIN[6]), .ZN(n288) );
  OAI22_X1 U22 ( .A1(n43), .A2(n261), .B1(n258), .B2(n287), .ZN(n97) );
  INV_X1 U23 ( .A(DIN[7]), .ZN(n287) );
  OAI22_X1 U24 ( .A1(n44), .A2(n261), .B1(n258), .B2(n286), .ZN(n98) );
  INV_X1 U25 ( .A(DIN[8]), .ZN(n286) );
  OAI22_X1 U26 ( .A1(n45), .A2(n261), .B1(n258), .B2(n285), .ZN(n99) );
  INV_X1 U27 ( .A(DIN[9]), .ZN(n285) );
  OAI22_X1 U28 ( .A1(n46), .A2(n260), .B1(n258), .B2(n284), .ZN(n90) );
  INV_X1 U29 ( .A(DIN[10]), .ZN(n284) );
  OAI22_X1 U30 ( .A1(n36), .A2(n260), .B1(n257), .B2(n294), .ZN(n89) );
  INV_X1 U31 ( .A(DIN[0]), .ZN(n294) );
  OAI22_X1 U32 ( .A1(n47), .A2(n260), .B1(n257), .B2(n283), .ZN(n88) );
  INV_X1 U33 ( .A(DIN[11]), .ZN(n283) );
  OAI22_X1 U34 ( .A1(n48), .A2(n260), .B1(n257), .B2(n282), .ZN(n87) );
  INV_X1 U35 ( .A(DIN[12]), .ZN(n282) );
  OAI22_X1 U36 ( .A1(n49), .A2(n260), .B1(n257), .B2(n281), .ZN(n86) );
  INV_X1 U37 ( .A(DIN[13]), .ZN(n281) );
  OAI22_X1 U38 ( .A1(n50), .A2(n260), .B1(n257), .B2(n280), .ZN(n85) );
  INV_X1 U39 ( .A(DIN[14]), .ZN(n280) );
  OAI22_X1 U40 ( .A1(n51), .A2(n259), .B1(n256), .B2(n279), .ZN(n68) );
  INV_X1 U41 ( .A(DIN[15]), .ZN(n279) );
  OAI22_X1 U42 ( .A1(n52), .A2(n259), .B1(n256), .B2(n269), .ZN(n69) );
  INV_X1 U43 ( .A(DIN[16]), .ZN(n269) );
  OAI22_X1 U44 ( .A1(n53), .A2(n259), .B1(n256), .B2(n270), .ZN(n70) );
  INV_X1 U45 ( .A(DIN[17]), .ZN(n270) );
  OAI22_X1 U46 ( .A1(n54), .A2(n259), .B1(n256), .B2(n271), .ZN(n71) );
  INV_X1 U47 ( .A(DIN[18]), .ZN(n271) );
  OAI22_X1 U48 ( .A1(n55), .A2(n259), .B1(n256), .B2(n272), .ZN(n72) );
  INV_X1 U49 ( .A(DIN[19]), .ZN(n272) );
  OAI22_X1 U50 ( .A1(n56), .A2(n259), .B1(n256), .B2(n273), .ZN(n73) );
  INV_X1 U51 ( .A(DIN[20]), .ZN(n273) );
  OAI22_X1 U52 ( .A1(n57), .A2(n259), .B1(n256), .B2(n274), .ZN(n74) );
  INV_X1 U53 ( .A(DIN[21]), .ZN(n274) );
  OAI22_X1 U54 ( .A1(n58), .A2(n259), .B1(n256), .B2(n275), .ZN(n75) );
  INV_X1 U55 ( .A(DIN[22]), .ZN(n275) );
  OAI22_X1 U56 ( .A1(n59), .A2(n259), .B1(n256), .B2(n276), .ZN(n76) );
  INV_X1 U57 ( .A(DIN[23]), .ZN(n276) );
  OAI22_X1 U58 ( .A1(n60), .A2(n259), .B1(n256), .B2(n277), .ZN(n77) );
  INV_X1 U59 ( .A(DIN[24]), .ZN(n277) );
  OAI22_X1 U60 ( .A1(n61), .A2(n259), .B1(n256), .B2(n278), .ZN(n78) );
  INV_X1 U61 ( .A(DIN[25]), .ZN(n278) );
  OAI22_X1 U62 ( .A1(n62), .A2(n260), .B1(n257), .B2(n262), .ZN(n79) );
  INV_X1 U63 ( .A(DIN[26]), .ZN(n262) );
  OAI22_X1 U64 ( .A1(n63), .A2(n260), .B1(n257), .B2(n263), .ZN(n80) );
  INV_X1 U65 ( .A(DIN[27]), .ZN(n263) );
  OAI22_X1 U66 ( .A1(n64), .A2(n260), .B1(n257), .B2(n264), .ZN(n81) );
  INV_X1 U67 ( .A(DIN[28]), .ZN(n264) );
  OAI22_X1 U68 ( .A1(n65), .A2(n260), .B1(n257), .B2(n265), .ZN(n82) );
  INV_X1 U69 ( .A(DIN[29]), .ZN(n265) );
  OAI22_X1 U70 ( .A1(n66), .A2(n260), .B1(n257), .B2(n266), .ZN(n83) );
  INV_X1 U71 ( .A(DIN[30]), .ZN(n266) );
  NAND2_X1 U72 ( .A1(n268), .A2(RST), .ZN(n34) );
  INV_X1 U73 ( .A(EN), .ZN(n268) );
  OAI22_X1 U74 ( .A1(n67), .A2(n260), .B1(n257), .B2(n267), .ZN(n84) );
  INV_X1 U75 ( .A(DIN[31]), .ZN(n267) );
endmodule


module REGISTER_GENERIC_WIDTH5_0 ( CLK, RST, EN, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST, EN;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n2, n3, n4, n5, n6,
         n7, n8, n44;

  DFF_X1 \DOUT_reg[4]  ( .D(n14), .CK(CLK), .Q(DOUT[4]), .QN(n13) );
  DFF_X1 \DOUT_reg[3]  ( .D(n15), .CK(CLK), .Q(DOUT[3]), .QN(n12) );
  DFF_X1 \DOUT_reg[2]  ( .D(n16), .CK(CLK), .Q(DOUT[2]), .QN(n11) );
  DFF_X1 \DOUT_reg[1]  ( .D(n17), .CK(CLK), .Q(DOUT[1]), .QN(n10) );
  DFF_X1 \DOUT_reg[0]  ( .D(n18), .CK(CLK), .Q(DOUT[0]), .QN(n9) );
  AND2_X1 U3 ( .A1(RST), .A2(n2), .ZN(n4) );
  NAND2_X1 U4 ( .A1(n44), .A2(RST), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n44) );
  OAI21_X1 U6 ( .B1(n9), .B2(n2), .A(n3), .ZN(n18) );
  NAND2_X1 U7 ( .A1(DIN[0]), .A2(n4), .ZN(n3) );
  OAI21_X1 U8 ( .B1(n10), .B2(n2), .A(n5), .ZN(n17) );
  NAND2_X1 U9 ( .A1(DIN[1]), .A2(n4), .ZN(n5) );
  OAI21_X1 U10 ( .B1(n11), .B2(n2), .A(n6), .ZN(n16) );
  NAND2_X1 U11 ( .A1(DIN[2]), .A2(n4), .ZN(n6) );
  OAI21_X1 U12 ( .B1(n12), .B2(n2), .A(n7), .ZN(n15) );
  NAND2_X1 U13 ( .A1(DIN[3]), .A2(n4), .ZN(n7) );
  OAI21_X1 U14 ( .B1(n13), .B2(n2), .A(n8), .ZN(n14) );
  NAND2_X1 U15 ( .A1(DIN[4]), .A2(n4), .ZN(n8) );
endmodule


module REGISTER_GENERIC_WIDTH32_7 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298;

  DFF_X1 \DOUT_reg[31]  ( .D(n68), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[30]  ( .D(n69), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[29]  ( .D(n70), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[28]  ( .D(n71), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[27]  ( .D(n72), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n73), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[25]  ( .D(n74), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[24]  ( .D(n75), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[22]  ( .D(n77), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[21]  ( .D(n78), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[20]  ( .D(n79), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n80), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n81), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n83), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n84), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n89), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n90), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n91), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n92), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n93), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n94), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n95), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n96), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n97), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n98), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n262) );
  BUF_X1 U4 ( .A(n35), .Z(n261) );
  BUF_X1 U5 ( .A(n35), .Z(n260) );
  NAND2_X1 U6 ( .A1(RST), .A2(n263), .ZN(n35) );
  BUF_X1 U7 ( .A(n34), .Z(n265) );
  BUF_X1 U8 ( .A(n34), .Z(n263) );
  BUF_X1 U9 ( .A(n34), .Z(n264) );
  OAI22_X1 U10 ( .A1(n36), .A2(n265), .B1(n262), .B2(n296), .ZN(n99) );
  INV_X1 U11 ( .A(DIN[0]), .ZN(n296) );
  OAI22_X1 U12 ( .A1(n37), .A2(n265), .B1(n262), .B2(n295), .ZN(n98) );
  INV_X1 U13 ( .A(DIN[1]), .ZN(n295) );
  OAI22_X1 U14 ( .A1(n38), .A2(n265), .B1(n262), .B2(n294), .ZN(n97) );
  INV_X1 U15 ( .A(DIN[2]), .ZN(n294) );
  OAI22_X1 U16 ( .A1(n39), .A2(n265), .B1(n262), .B2(n293), .ZN(n96) );
  INV_X1 U17 ( .A(DIN[3]), .ZN(n293) );
  OAI22_X1 U18 ( .A1(n40), .A2(n265), .B1(n262), .B2(n292), .ZN(n95) );
  INV_X1 U19 ( .A(DIN[4]), .ZN(n292) );
  OAI22_X1 U20 ( .A1(n41), .A2(n265), .B1(n262), .B2(n291), .ZN(n94) );
  INV_X1 U21 ( .A(DIN[5]), .ZN(n291) );
  OAI22_X1 U22 ( .A1(n42), .A2(n265), .B1(n262), .B2(n290), .ZN(n93) );
  INV_X1 U23 ( .A(DIN[6]), .ZN(n290) );
  OAI22_X1 U24 ( .A1(n43), .A2(n265), .B1(n262), .B2(n289), .ZN(n92) );
  INV_X1 U25 ( .A(DIN[7]), .ZN(n289) );
  OAI22_X1 U26 ( .A1(n44), .A2(n265), .B1(n262), .B2(n288), .ZN(n91) );
  INV_X1 U27 ( .A(DIN[8]), .ZN(n288) );
  OAI22_X1 U28 ( .A1(n45), .A2(n264), .B1(n262), .B2(n287), .ZN(n90) );
  INV_X1 U29 ( .A(DIN[9]), .ZN(n287) );
  OAI22_X1 U30 ( .A1(n46), .A2(n264), .B1(n261), .B2(n286), .ZN(n89) );
  INV_X1 U31 ( .A(DIN[10]), .ZN(n286) );
  OAI22_X1 U32 ( .A1(n47), .A2(n264), .B1(n261), .B2(n285), .ZN(n88) );
  INV_X1 U33 ( .A(DIN[11]), .ZN(n285) );
  OAI22_X1 U34 ( .A1(n48), .A2(n264), .B1(n261), .B2(n284), .ZN(n87) );
  INV_X1 U35 ( .A(DIN[12]), .ZN(n284) );
  OAI22_X1 U36 ( .A1(n49), .A2(n264), .B1(n261), .B2(n283), .ZN(n86) );
  INV_X1 U37 ( .A(DIN[13]), .ZN(n283) );
  OAI22_X1 U38 ( .A1(n50), .A2(n264), .B1(n261), .B2(n282), .ZN(n85) );
  INV_X1 U39 ( .A(DIN[14]), .ZN(n282) );
  OAI22_X1 U40 ( .A1(n51), .A2(n264), .B1(n261), .B2(n281), .ZN(n84) );
  INV_X1 U41 ( .A(DIN[15]), .ZN(n281) );
  OAI22_X1 U42 ( .A1(n52), .A2(n264), .B1(n261), .B2(n280), .ZN(n83) );
  INV_X1 U43 ( .A(DIN[16]), .ZN(n280) );
  OAI22_X1 U44 ( .A1(n53), .A2(n264), .B1(n261), .B2(n279), .ZN(n82) );
  INV_X1 U45 ( .A(DIN[17]), .ZN(n279) );
  OAI22_X1 U46 ( .A1(n54), .A2(n264), .B1(n261), .B2(n278), .ZN(n81) );
  INV_X1 U47 ( .A(DIN[18]), .ZN(n278) );
  OAI22_X1 U48 ( .A1(n55), .A2(n264), .B1(n261), .B2(n277), .ZN(n80) );
  INV_X1 U49 ( .A(DIN[19]), .ZN(n277) );
  OAI22_X1 U50 ( .A1(n56), .A2(n264), .B1(n261), .B2(n276), .ZN(n79) );
  INV_X1 U51 ( .A(DIN[20]), .ZN(n276) );
  OAI22_X1 U52 ( .A1(n57), .A2(n263), .B1(n260), .B2(n275), .ZN(n78) );
  INV_X1 U53 ( .A(DIN[21]), .ZN(n275) );
  OAI22_X1 U54 ( .A1(n58), .A2(n263), .B1(n260), .B2(n274), .ZN(n77) );
  INV_X1 U55 ( .A(DIN[22]), .ZN(n274) );
  OAI22_X1 U56 ( .A1(n59), .A2(n263), .B1(n260), .B2(n273), .ZN(n76) );
  INV_X1 U57 ( .A(DIN[23]), .ZN(n273) );
  OAI22_X1 U58 ( .A1(n60), .A2(n263), .B1(n260), .B2(n272), .ZN(n75) );
  INV_X1 U59 ( .A(DIN[24]), .ZN(n272) );
  OAI22_X1 U60 ( .A1(n61), .A2(n263), .B1(n260), .B2(n271), .ZN(n74) );
  INV_X1 U61 ( .A(DIN[25]), .ZN(n271) );
  OAI22_X1 U62 ( .A1(n62), .A2(n263), .B1(n260), .B2(n270), .ZN(n73) );
  INV_X1 U63 ( .A(DIN[26]), .ZN(n270) );
  OAI22_X1 U64 ( .A1(n63), .A2(n263), .B1(n260), .B2(n269), .ZN(n72) );
  INV_X1 U65 ( .A(DIN[27]), .ZN(n269) );
  OAI22_X1 U66 ( .A1(n64), .A2(n263), .B1(n260), .B2(n268), .ZN(n71) );
  INV_X1 U67 ( .A(DIN[28]), .ZN(n268) );
  OAI22_X1 U68 ( .A1(n65), .A2(n263), .B1(n260), .B2(n267), .ZN(n70) );
  INV_X1 U69 ( .A(DIN[29]), .ZN(n267) );
  OAI22_X1 U70 ( .A1(n66), .A2(n263), .B1(n260), .B2(n266), .ZN(n69) );
  INV_X1 U71 ( .A(DIN[30]), .ZN(n266) );
  OAI22_X1 U72 ( .A1(n67), .A2(n263), .B1(n260), .B2(n297), .ZN(n68) );
  INV_X1 U73 ( .A(DIN[31]), .ZN(n297) );
  NAND2_X1 U74 ( .A1(n298), .A2(RST), .ZN(n34) );
  INV_X1 U75 ( .A(EN), .ZN(n298) );
endmodule


module MUX21_GENERIC_NBIT32_5 ( S1, S0, SEL, Y );
  input [31:0] S1;
  input [31:0] S0;
  output [31:0] Y;
  input SEL;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390;

  INV_X1 U1 ( .A(n390), .ZN(n380) );
  INV_X1 U2 ( .A(n390), .ZN(n381) );
  BUF_X1 U3 ( .A(n379), .Z(n388) );
  BUF_X1 U4 ( .A(n378), .Z(n387) );
  BUF_X1 U5 ( .A(n378), .Z(n385) );
  BUF_X1 U6 ( .A(n377), .Z(n384) );
  BUF_X1 U7 ( .A(n378), .Z(n386) );
  BUF_X1 U8 ( .A(n377), .Z(n383) );
  BUF_X1 U9 ( .A(n377), .Z(n382) );
  BUF_X1 U10 ( .A(n379), .Z(n390) );
  BUF_X1 U11 ( .A(n379), .Z(n389) );
  INV_X1 U12 ( .A(n34), .ZN(Y[31]) );
  AOI22_X1 U13 ( .A1(S0[31]), .A2(n380), .B1(n389), .B2(S1[31]), .ZN(n34) );
  INV_X1 U14 ( .A(n65), .ZN(Y[0]) );
  AOI22_X1 U15 ( .A1(S0[0]), .A2(n380), .B1(S1[0]), .B2(n389), .ZN(n65) );
  INV_X1 U16 ( .A(n64), .ZN(Y[1]) );
  AOI22_X1 U17 ( .A1(S0[1]), .A2(n380), .B1(S1[1]), .B2(n389), .ZN(n64) );
  INV_X1 U18 ( .A(n63), .ZN(Y[2]) );
  AOI22_X1 U19 ( .A1(S0[2]), .A2(n380), .B1(S1[2]), .B2(n389), .ZN(n63) );
  INV_X1 U20 ( .A(n62), .ZN(Y[3]) );
  AOI22_X1 U21 ( .A1(S0[3]), .A2(n380), .B1(S1[3]), .B2(n388), .ZN(n62) );
  INV_X1 U22 ( .A(n61), .ZN(Y[4]) );
  AOI22_X1 U23 ( .A1(S0[4]), .A2(n380), .B1(S1[4]), .B2(n388), .ZN(n61) );
  INV_X1 U24 ( .A(n60), .ZN(Y[5]) );
  AOI22_X1 U25 ( .A1(S0[5]), .A2(n380), .B1(S1[5]), .B2(n388), .ZN(n60) );
  INV_X1 U26 ( .A(n59), .ZN(Y[6]) );
  AOI22_X1 U27 ( .A1(S0[6]), .A2(n380), .B1(S1[6]), .B2(n388), .ZN(n59) );
  INV_X1 U28 ( .A(n58), .ZN(Y[7]) );
  AOI22_X1 U29 ( .A1(S0[7]), .A2(n380), .B1(S1[7]), .B2(n387), .ZN(n58) );
  INV_X1 U30 ( .A(n57), .ZN(Y[8]) );
  AOI22_X1 U31 ( .A1(S0[8]), .A2(n380), .B1(S1[8]), .B2(n387), .ZN(n57) );
  INV_X1 U32 ( .A(n56), .ZN(Y[9]) );
  AOI22_X1 U33 ( .A1(S0[9]), .A2(n380), .B1(S1[9]), .B2(n387), .ZN(n56) );
  INV_X1 U34 ( .A(n55), .ZN(Y[10]) );
  AOI22_X1 U35 ( .A1(S0[10]), .A2(n380), .B1(S1[10]), .B2(n387), .ZN(n55) );
  INV_X1 U36 ( .A(n54), .ZN(Y[11]) );
  AOI22_X1 U37 ( .A1(S0[11]), .A2(n380), .B1(S1[11]), .B2(n386), .ZN(n54) );
  INV_X1 U38 ( .A(n53), .ZN(Y[12]) );
  AOI22_X1 U39 ( .A1(S0[12]), .A2(n381), .B1(S1[12]), .B2(n386), .ZN(n53) );
  INV_X1 U40 ( .A(n52), .ZN(Y[13]) );
  AOI22_X1 U41 ( .A1(S0[13]), .A2(n381), .B1(S1[13]), .B2(n386), .ZN(n52) );
  INV_X1 U42 ( .A(n51), .ZN(Y[14]) );
  AOI22_X1 U43 ( .A1(S0[14]), .A2(n381), .B1(S1[14]), .B2(n385), .ZN(n51) );
  INV_X1 U44 ( .A(n50), .ZN(Y[15]) );
  AOI22_X1 U45 ( .A1(S0[15]), .A2(n381), .B1(S1[15]), .B2(n385), .ZN(n50) );
  INV_X1 U46 ( .A(n49), .ZN(Y[16]) );
  AOI22_X1 U47 ( .A1(S0[16]), .A2(n381), .B1(S1[16]), .B2(n385), .ZN(n49) );
  INV_X1 U48 ( .A(n48), .ZN(Y[17]) );
  AOI22_X1 U49 ( .A1(S0[17]), .A2(n381), .B1(S1[17]), .B2(n385), .ZN(n48) );
  INV_X1 U50 ( .A(n47), .ZN(Y[18]) );
  AOI22_X1 U51 ( .A1(S0[18]), .A2(n381), .B1(S1[18]), .B2(n384), .ZN(n47) );
  INV_X1 U52 ( .A(n46), .ZN(Y[19]) );
  AOI22_X1 U53 ( .A1(S0[19]), .A2(n381), .B1(S1[19]), .B2(n384), .ZN(n46) );
  INV_X1 U54 ( .A(n45), .ZN(Y[20]) );
  AOI22_X1 U55 ( .A1(S0[20]), .A2(n381), .B1(S1[20]), .B2(n384), .ZN(n45) );
  INV_X1 U56 ( .A(n44), .ZN(Y[21]) );
  AOI22_X1 U57 ( .A1(S0[21]), .A2(n381), .B1(S1[21]), .B2(n384), .ZN(n44) );
  INV_X1 U58 ( .A(n43), .ZN(Y[22]) );
  AOI22_X1 U59 ( .A1(S0[22]), .A2(n381), .B1(S1[22]), .B2(n383), .ZN(n43) );
  INV_X1 U60 ( .A(n42), .ZN(Y[23]) );
  AOI22_X1 U61 ( .A1(S0[23]), .A2(n381), .B1(S1[23]), .B2(n386), .ZN(n42) );
  INV_X1 U62 ( .A(n41), .ZN(Y[24]) );
  AOI22_X1 U63 ( .A1(S0[24]), .A2(n381), .B1(S1[24]), .B2(n383), .ZN(n41) );
  INV_X1 U64 ( .A(n40), .ZN(Y[25]) );
  AOI22_X1 U65 ( .A1(S0[25]), .A2(n380), .B1(S1[25]), .B2(n383), .ZN(n40) );
  INV_X1 U66 ( .A(n39), .ZN(Y[26]) );
  AOI22_X1 U67 ( .A1(S0[26]), .A2(n381), .B1(S1[26]), .B2(n383), .ZN(n39) );
  INV_X1 U68 ( .A(n38), .ZN(Y[27]) );
  AOI22_X1 U69 ( .A1(S0[27]), .A2(n380), .B1(S1[27]), .B2(n382), .ZN(n38) );
  INV_X1 U70 ( .A(n37), .ZN(Y[28]) );
  AOI22_X1 U71 ( .A1(S0[28]), .A2(n381), .B1(S1[28]), .B2(n382), .ZN(n37) );
  INV_X1 U72 ( .A(n36), .ZN(Y[29]) );
  AOI22_X1 U73 ( .A1(S0[29]), .A2(n380), .B1(S1[29]), .B2(n382), .ZN(n36) );
  INV_X1 U74 ( .A(n35), .ZN(Y[30]) );
  AOI22_X1 U75 ( .A1(S0[30]), .A2(n381), .B1(S1[30]), .B2(n382), .ZN(n35) );
  BUF_X1 U76 ( .A(SEL), .Z(n379) );
  BUF_X1 U77 ( .A(SEL), .Z(n378) );
  BUF_X1 U78 ( .A(SEL), .Z(n377) );
endmodule


module MUX21_GENERIC_NBIT32_4 ( S1, S0, SEL, Y );
  input [31:0] S1;
  input [31:0] S0;
  output [31:0] Y;
  input SEL;
  wire   n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454;

  INV_X1 U1 ( .A(n390), .ZN(n380) );
  INV_X1 U2 ( .A(n390), .ZN(n381) );
  BUF_X1 U3 ( .A(n379), .Z(n388) );
  BUF_X1 U4 ( .A(n378), .Z(n387) );
  BUF_X1 U5 ( .A(n378), .Z(n385) );
  BUF_X1 U6 ( .A(n377), .Z(n384) );
  BUF_X1 U7 ( .A(n378), .Z(n386) );
  BUF_X1 U8 ( .A(n377), .Z(n383) );
  BUF_X1 U9 ( .A(n377), .Z(n382) );
  BUF_X1 U10 ( .A(n379), .Z(n390) );
  BUF_X1 U11 ( .A(n379), .Z(n389) );
  INV_X1 U12 ( .A(n454), .ZN(Y[31]) );
  AOI22_X1 U13 ( .A1(S0[31]), .A2(n380), .B1(n389), .B2(S1[31]), .ZN(n454) );
  INV_X1 U14 ( .A(n423), .ZN(Y[0]) );
  AOI22_X1 U15 ( .A1(S0[0]), .A2(n380), .B1(S1[0]), .B2(n389), .ZN(n423) );
  INV_X1 U16 ( .A(n424), .ZN(Y[1]) );
  AOI22_X1 U17 ( .A1(S0[1]), .A2(n380), .B1(S1[1]), .B2(n389), .ZN(n424) );
  INV_X1 U18 ( .A(n425), .ZN(Y[2]) );
  AOI22_X1 U19 ( .A1(S0[2]), .A2(n380), .B1(S1[2]), .B2(n389), .ZN(n425) );
  INV_X1 U20 ( .A(n426), .ZN(Y[3]) );
  AOI22_X1 U21 ( .A1(S0[3]), .A2(n380), .B1(S1[3]), .B2(n388), .ZN(n426) );
  INV_X1 U22 ( .A(n427), .ZN(Y[4]) );
  AOI22_X1 U23 ( .A1(S0[4]), .A2(n380), .B1(S1[4]), .B2(n388), .ZN(n427) );
  INV_X1 U24 ( .A(n428), .ZN(Y[5]) );
  AOI22_X1 U25 ( .A1(S0[5]), .A2(n380), .B1(S1[5]), .B2(n388), .ZN(n428) );
  INV_X1 U26 ( .A(n429), .ZN(Y[6]) );
  AOI22_X1 U27 ( .A1(S0[6]), .A2(n380), .B1(S1[6]), .B2(n388), .ZN(n429) );
  INV_X1 U28 ( .A(n430), .ZN(Y[7]) );
  AOI22_X1 U29 ( .A1(S0[7]), .A2(n380), .B1(S1[7]), .B2(n387), .ZN(n430) );
  INV_X1 U30 ( .A(n431), .ZN(Y[8]) );
  AOI22_X1 U31 ( .A1(S0[8]), .A2(n380), .B1(S1[8]), .B2(n387), .ZN(n431) );
  INV_X1 U32 ( .A(n432), .ZN(Y[9]) );
  AOI22_X1 U33 ( .A1(S0[9]), .A2(n380), .B1(S1[9]), .B2(n387), .ZN(n432) );
  INV_X1 U34 ( .A(n433), .ZN(Y[10]) );
  AOI22_X1 U35 ( .A1(S0[10]), .A2(n380), .B1(S1[10]), .B2(n387), .ZN(n433) );
  INV_X1 U36 ( .A(n434), .ZN(Y[11]) );
  AOI22_X1 U37 ( .A1(S0[11]), .A2(n380), .B1(S1[11]), .B2(n386), .ZN(n434) );
  INV_X1 U38 ( .A(n435), .ZN(Y[12]) );
  AOI22_X1 U39 ( .A1(S0[12]), .A2(n381), .B1(S1[12]), .B2(n386), .ZN(n435) );
  INV_X1 U40 ( .A(n436), .ZN(Y[13]) );
  AOI22_X1 U41 ( .A1(S0[13]), .A2(n381), .B1(S1[13]), .B2(n386), .ZN(n436) );
  INV_X1 U42 ( .A(n437), .ZN(Y[14]) );
  AOI22_X1 U43 ( .A1(S0[14]), .A2(n381), .B1(S1[14]), .B2(n385), .ZN(n437) );
  INV_X1 U44 ( .A(n438), .ZN(Y[15]) );
  AOI22_X1 U45 ( .A1(S0[15]), .A2(n381), .B1(S1[15]), .B2(n385), .ZN(n438) );
  INV_X1 U46 ( .A(n439), .ZN(Y[16]) );
  AOI22_X1 U47 ( .A1(S0[16]), .A2(n381), .B1(S1[16]), .B2(n385), .ZN(n439) );
  INV_X1 U48 ( .A(n440), .ZN(Y[17]) );
  AOI22_X1 U49 ( .A1(S0[17]), .A2(n381), .B1(S1[17]), .B2(n385), .ZN(n440) );
  INV_X1 U50 ( .A(n441), .ZN(Y[18]) );
  AOI22_X1 U51 ( .A1(S0[18]), .A2(n381), .B1(S1[18]), .B2(n384), .ZN(n441) );
  INV_X1 U52 ( .A(n442), .ZN(Y[19]) );
  AOI22_X1 U53 ( .A1(S0[19]), .A2(n381), .B1(S1[19]), .B2(n384), .ZN(n442) );
  INV_X1 U54 ( .A(n443), .ZN(Y[20]) );
  AOI22_X1 U55 ( .A1(S0[20]), .A2(n381), .B1(S1[20]), .B2(n384), .ZN(n443) );
  INV_X1 U56 ( .A(n444), .ZN(Y[21]) );
  AOI22_X1 U57 ( .A1(S0[21]), .A2(n381), .B1(S1[21]), .B2(n384), .ZN(n444) );
  INV_X1 U58 ( .A(n445), .ZN(Y[22]) );
  AOI22_X1 U59 ( .A1(S0[22]), .A2(n381), .B1(S1[22]), .B2(n383), .ZN(n445) );
  INV_X1 U60 ( .A(n446), .ZN(Y[23]) );
  AOI22_X1 U61 ( .A1(S0[23]), .A2(n381), .B1(S1[23]), .B2(n386), .ZN(n446) );
  INV_X1 U62 ( .A(n447), .ZN(Y[24]) );
  AOI22_X1 U63 ( .A1(S0[24]), .A2(n381), .B1(S1[24]), .B2(n383), .ZN(n447) );
  INV_X1 U64 ( .A(n448), .ZN(Y[25]) );
  AOI22_X1 U65 ( .A1(S0[25]), .A2(n380), .B1(S1[25]), .B2(n383), .ZN(n448) );
  INV_X1 U66 ( .A(n449), .ZN(Y[26]) );
  AOI22_X1 U67 ( .A1(S0[26]), .A2(n381), .B1(S1[26]), .B2(n383), .ZN(n449) );
  INV_X1 U68 ( .A(n450), .ZN(Y[27]) );
  AOI22_X1 U69 ( .A1(S0[27]), .A2(n380), .B1(S1[27]), .B2(n382), .ZN(n450) );
  INV_X1 U70 ( .A(n451), .ZN(Y[28]) );
  AOI22_X1 U71 ( .A1(S0[28]), .A2(n381), .B1(S1[28]), .B2(n382), .ZN(n451) );
  INV_X1 U72 ( .A(n452), .ZN(Y[29]) );
  AOI22_X1 U73 ( .A1(S0[29]), .A2(n380), .B1(S1[29]), .B2(n382), .ZN(n452) );
  INV_X1 U74 ( .A(n453), .ZN(Y[30]) );
  AOI22_X1 U75 ( .A1(S0[30]), .A2(n381), .B1(S1[30]), .B2(n382), .ZN(n453) );
  BUF_X1 U76 ( .A(SEL), .Z(n379) );
  BUF_X1 U77 ( .A(SEL), .Z(n378) );
  BUF_X1 U78 ( .A(SEL), .Z(n377) );
endmodule


module MUX31_GENERIC_NBIT32_0 ( S2, S1, S0, SEL, Y );
  input [31:0] S2;
  input [31:0] S1;
  input [31:0] S0;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n390, n391;

  BUF_X1 U2 ( .A(n37), .Z(n352) );
  BUF_X1 U3 ( .A(n37), .Z(n353) );
  BUF_X1 U4 ( .A(n38), .Z(n349) );
  BUF_X1 U5 ( .A(n38), .Z(n350) );
  BUF_X1 U6 ( .A(n37), .Z(n354) );
  BUF_X1 U7 ( .A(n38), .Z(n351) );
  BUF_X1 U8 ( .A(n36), .Z(n355) );
  BUF_X1 U9 ( .A(n36), .Z(n356) );
  NOR3_X1 U10 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n391), .ZN(n37) );
  BUF_X1 U11 ( .A(n36), .Z(n357) );
  AND3_X1 U12 ( .A1(n390), .A2(n391), .A3(SEL[2]), .ZN(n38) );
  INV_X1 U13 ( .A(SEL[0]), .ZN(n390) );
  NOR3_X1 U14 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n390), .ZN(n36) );
  INV_X1 U15 ( .A(SEL[1]), .ZN(n391) );
  INV_X1 U16 ( .A(n35), .ZN(Y[31]) );
  AOI222_X1 U17 ( .A1(S0[31]), .A2(n357), .B1(S1[31]), .B2(n354), .C1(S2[31]), 
        .C2(n351), .ZN(n35) );
  INV_X1 U18 ( .A(n69), .ZN(Y[0]) );
  AOI222_X1 U19 ( .A1(S0[0]), .A2(n355), .B1(S1[0]), .B2(n352), .C1(S2[0]), 
        .C2(n349), .ZN(n69) );
  INV_X1 U20 ( .A(n68), .ZN(Y[1]) );
  AOI222_X1 U21 ( .A1(S0[1]), .A2(n355), .B1(S1[1]), .B2(n352), .C1(S2[1]), 
        .C2(n349), .ZN(n68) );
  INV_X1 U22 ( .A(n67), .ZN(Y[2]) );
  AOI222_X1 U23 ( .A1(S0[2]), .A2(n355), .B1(S1[2]), .B2(n352), .C1(S2[2]), 
        .C2(n349), .ZN(n67) );
  INV_X1 U24 ( .A(n66), .ZN(Y[3]) );
  AOI222_X1 U25 ( .A1(S0[3]), .A2(n355), .B1(S1[3]), .B2(n352), .C1(S2[3]), 
        .C2(n349), .ZN(n66) );
  INV_X1 U26 ( .A(n65), .ZN(Y[4]) );
  AOI222_X1 U27 ( .A1(S0[4]), .A2(n355), .B1(S1[4]), .B2(n352), .C1(S2[4]), 
        .C2(n349), .ZN(n65) );
  INV_X1 U28 ( .A(n64), .ZN(Y[5]) );
  AOI222_X1 U29 ( .A1(S0[5]), .A2(n355), .B1(S1[5]), .B2(n352), .C1(S2[5]), 
        .C2(n349), .ZN(n64) );
  INV_X1 U30 ( .A(n63), .ZN(Y[6]) );
  AOI222_X1 U31 ( .A1(S0[6]), .A2(n355), .B1(S1[6]), .B2(n352), .C1(S2[6]), 
        .C2(n349), .ZN(n63) );
  INV_X1 U32 ( .A(n62), .ZN(Y[7]) );
  AOI222_X1 U33 ( .A1(S0[7]), .A2(n355), .B1(S1[7]), .B2(n352), .C1(S2[7]), 
        .C2(n349), .ZN(n62) );
  INV_X1 U34 ( .A(n61), .ZN(Y[8]) );
  AOI222_X1 U35 ( .A1(S0[8]), .A2(n355), .B1(S1[8]), .B2(n352), .C1(S2[8]), 
        .C2(n349), .ZN(n61) );
  INV_X1 U36 ( .A(n60), .ZN(Y[9]) );
  AOI222_X1 U37 ( .A1(S0[9]), .A2(n355), .B1(S1[9]), .B2(n352), .C1(S2[9]), 
        .C2(n349), .ZN(n60) );
  INV_X1 U38 ( .A(n59), .ZN(Y[10]) );
  AOI222_X1 U39 ( .A1(S0[10]), .A2(n355), .B1(S1[10]), .B2(n352), .C1(S2[10]), 
        .C2(n349), .ZN(n59) );
  INV_X1 U40 ( .A(n58), .ZN(Y[11]) );
  AOI222_X1 U41 ( .A1(S0[11]), .A2(n356), .B1(S1[11]), .B2(n352), .C1(S2[11]), 
        .C2(n349), .ZN(n58) );
  INV_X1 U42 ( .A(n57), .ZN(Y[12]) );
  AOI222_X1 U43 ( .A1(S0[12]), .A2(n356), .B1(S1[12]), .B2(n353), .C1(S2[12]), 
        .C2(n350), .ZN(n57) );
  INV_X1 U44 ( .A(n56), .ZN(Y[13]) );
  AOI222_X1 U45 ( .A1(S0[13]), .A2(n356), .B1(S1[13]), .B2(n353), .C1(S2[13]), 
        .C2(n350), .ZN(n56) );
  INV_X1 U46 ( .A(n55), .ZN(Y[14]) );
  AOI222_X1 U47 ( .A1(S0[14]), .A2(n356), .B1(S1[14]), .B2(n353), .C1(S2[14]), 
        .C2(n350), .ZN(n55) );
  INV_X1 U48 ( .A(n54), .ZN(Y[15]) );
  AOI222_X1 U49 ( .A1(S0[15]), .A2(n356), .B1(S1[15]), .B2(n353), .C1(S2[15]), 
        .C2(n350), .ZN(n54) );
  INV_X1 U50 ( .A(n53), .ZN(Y[16]) );
  AOI222_X1 U51 ( .A1(S0[16]), .A2(n356), .B1(S1[16]), .B2(n353), .C1(S2[16]), 
        .C2(n350), .ZN(n53) );
  INV_X1 U52 ( .A(n52), .ZN(Y[17]) );
  AOI222_X1 U53 ( .A1(S0[17]), .A2(n356), .B1(S1[17]), .B2(n353), .C1(S2[17]), 
        .C2(n350), .ZN(n52) );
  INV_X1 U54 ( .A(n51), .ZN(Y[18]) );
  AOI222_X1 U55 ( .A1(S0[18]), .A2(n356), .B1(S1[18]), .B2(n353), .C1(S2[18]), 
        .C2(n350), .ZN(n51) );
  INV_X1 U56 ( .A(n50), .ZN(Y[19]) );
  AOI222_X1 U57 ( .A1(S0[19]), .A2(n356), .B1(S1[19]), .B2(n353), .C1(S2[19]), 
        .C2(n350), .ZN(n50) );
  INV_X1 U58 ( .A(n49), .ZN(Y[20]) );
  AOI222_X1 U59 ( .A1(S0[20]), .A2(n356), .B1(S1[20]), .B2(n353), .C1(S2[20]), 
        .C2(n350), .ZN(n49) );
  INV_X1 U60 ( .A(n48), .ZN(Y[21]) );
  AOI222_X1 U61 ( .A1(S0[21]), .A2(n356), .B1(S1[21]), .B2(n353), .C1(S2[21]), 
        .C2(n350), .ZN(n48) );
  INV_X1 U62 ( .A(n47), .ZN(Y[22]) );
  AOI222_X1 U63 ( .A1(S0[22]), .A2(n357), .B1(S1[22]), .B2(n353), .C1(S2[22]), 
        .C2(n350), .ZN(n47) );
  INV_X1 U64 ( .A(n46), .ZN(Y[23]) );
  AOI222_X1 U65 ( .A1(S0[23]), .A2(n357), .B1(S1[23]), .B2(n353), .C1(S2[23]), 
        .C2(n350), .ZN(n46) );
  INV_X1 U66 ( .A(n45), .ZN(Y[24]) );
  AOI222_X1 U67 ( .A1(S0[24]), .A2(n357), .B1(S1[24]), .B2(n354), .C1(S2[24]), 
        .C2(n351), .ZN(n45) );
  INV_X1 U68 ( .A(n44), .ZN(Y[25]) );
  AOI222_X1 U69 ( .A1(S0[25]), .A2(n357), .B1(S1[25]), .B2(n354), .C1(S2[25]), 
        .C2(n351), .ZN(n44) );
  INV_X1 U70 ( .A(n43), .ZN(Y[26]) );
  AOI222_X1 U71 ( .A1(S0[26]), .A2(n357), .B1(S1[26]), .B2(n354), .C1(S2[26]), 
        .C2(n351), .ZN(n43) );
  INV_X1 U72 ( .A(n42), .ZN(Y[27]) );
  AOI222_X1 U73 ( .A1(S0[27]), .A2(n357), .B1(S1[27]), .B2(n354), .C1(S2[27]), 
        .C2(n351), .ZN(n42) );
  INV_X1 U74 ( .A(n41), .ZN(Y[28]) );
  AOI222_X1 U75 ( .A1(S0[28]), .A2(n357), .B1(S1[28]), .B2(n354), .C1(S2[28]), 
        .C2(n351), .ZN(n41) );
  INV_X1 U76 ( .A(n40), .ZN(Y[29]) );
  AOI222_X1 U77 ( .A1(S0[29]), .A2(n357), .B1(S1[29]), .B2(n354), .C1(S2[29]), 
        .C2(n351), .ZN(n40) );
  INV_X1 U78 ( .A(n39), .ZN(Y[30]) );
  AOI222_X1 U79 ( .A1(S0[30]), .A2(n357), .B1(S1[30]), .B2(n354), .C1(S2[30]), 
        .C2(n351), .ZN(n39) );
endmodule


module MUX31_GENERIC_NBIT32_4 ( S2, S1, S0, SEL, Y );
  input [31:0] S2;
  input [31:0] S1;
  input [31:0] S0;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n425, n426;

  BUF_X1 U2 ( .A(n37), .Z(n387) );
  BUF_X1 U3 ( .A(n37), .Z(n388) );
  BUF_X1 U4 ( .A(n38), .Z(n384) );
  BUF_X1 U5 ( .A(n38), .Z(n385) );
  BUF_X1 U6 ( .A(n37), .Z(n389) );
  BUF_X1 U7 ( .A(n38), .Z(n386) );
  BUF_X1 U8 ( .A(n36), .Z(n390) );
  BUF_X1 U9 ( .A(n36), .Z(n391) );
  NOR3_X1 U10 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n426), .ZN(n37) );
  BUF_X1 U11 ( .A(n36), .Z(n392) );
  AND3_X1 U12 ( .A1(n425), .A2(n426), .A3(SEL[2]), .ZN(n38) );
  INV_X1 U13 ( .A(SEL[0]), .ZN(n425) );
  NOR3_X1 U14 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n425), .ZN(n36) );
  INV_X1 U15 ( .A(SEL[1]), .ZN(n426) );
  INV_X1 U16 ( .A(n35), .ZN(Y[31]) );
  AOI222_X1 U17 ( .A1(S0[31]), .A2(n392), .B1(S1[31]), .B2(n389), .C1(S2[31]), 
        .C2(n386), .ZN(n35) );
  INV_X1 U18 ( .A(n69), .ZN(Y[0]) );
  AOI222_X1 U19 ( .A1(S0[0]), .A2(n390), .B1(S1[0]), .B2(n387), .C1(S2[0]), 
        .C2(n384), .ZN(n69) );
  INV_X1 U20 ( .A(n68), .ZN(Y[1]) );
  AOI222_X1 U21 ( .A1(S0[1]), .A2(n390), .B1(S1[1]), .B2(n387), .C1(S2[1]), 
        .C2(n384), .ZN(n68) );
  INV_X1 U22 ( .A(n67), .ZN(Y[2]) );
  AOI222_X1 U23 ( .A1(S0[2]), .A2(n390), .B1(S1[2]), .B2(n387), .C1(S2[2]), 
        .C2(n384), .ZN(n67) );
  INV_X1 U24 ( .A(n66), .ZN(Y[3]) );
  AOI222_X1 U25 ( .A1(S0[3]), .A2(n390), .B1(S1[3]), .B2(n387), .C1(S2[3]), 
        .C2(n384), .ZN(n66) );
  INV_X1 U26 ( .A(n65), .ZN(Y[4]) );
  AOI222_X1 U27 ( .A1(S0[4]), .A2(n390), .B1(S1[4]), .B2(n387), .C1(S2[4]), 
        .C2(n384), .ZN(n65) );
  INV_X1 U28 ( .A(n64), .ZN(Y[5]) );
  AOI222_X1 U29 ( .A1(S0[5]), .A2(n390), .B1(S1[5]), .B2(n387), .C1(S2[5]), 
        .C2(n384), .ZN(n64) );
  INV_X1 U30 ( .A(n63), .ZN(Y[6]) );
  AOI222_X1 U31 ( .A1(S0[6]), .A2(n390), .B1(S1[6]), .B2(n387), .C1(S2[6]), 
        .C2(n384), .ZN(n63) );
  INV_X1 U32 ( .A(n62), .ZN(Y[7]) );
  AOI222_X1 U33 ( .A1(S0[7]), .A2(n390), .B1(S1[7]), .B2(n387), .C1(S2[7]), 
        .C2(n384), .ZN(n62) );
  INV_X1 U34 ( .A(n61), .ZN(Y[8]) );
  AOI222_X1 U35 ( .A1(S0[8]), .A2(n390), .B1(S1[8]), .B2(n387), .C1(S2[8]), 
        .C2(n384), .ZN(n61) );
  INV_X1 U36 ( .A(n60), .ZN(Y[9]) );
  AOI222_X1 U37 ( .A1(S0[9]), .A2(n390), .B1(S1[9]), .B2(n387), .C1(S2[9]), 
        .C2(n384), .ZN(n60) );
  INV_X1 U38 ( .A(n59), .ZN(Y[10]) );
  AOI222_X1 U39 ( .A1(S0[10]), .A2(n390), .B1(S1[10]), .B2(n387), .C1(S2[10]), 
        .C2(n384), .ZN(n59) );
  INV_X1 U40 ( .A(n58), .ZN(Y[11]) );
  AOI222_X1 U41 ( .A1(S0[11]), .A2(n391), .B1(S1[11]), .B2(n387), .C1(S2[11]), 
        .C2(n384), .ZN(n58) );
  INV_X1 U42 ( .A(n57), .ZN(Y[12]) );
  AOI222_X1 U43 ( .A1(S0[12]), .A2(n391), .B1(S1[12]), .B2(n388), .C1(S2[12]), 
        .C2(n385), .ZN(n57) );
  INV_X1 U44 ( .A(n56), .ZN(Y[13]) );
  AOI222_X1 U45 ( .A1(S0[13]), .A2(n391), .B1(S1[13]), .B2(n388), .C1(S2[13]), 
        .C2(n385), .ZN(n56) );
  INV_X1 U46 ( .A(n55), .ZN(Y[14]) );
  AOI222_X1 U47 ( .A1(S0[14]), .A2(n391), .B1(S1[14]), .B2(n388), .C1(S2[14]), 
        .C2(n385), .ZN(n55) );
  INV_X1 U48 ( .A(n54), .ZN(Y[15]) );
  AOI222_X1 U49 ( .A1(S0[15]), .A2(n391), .B1(S1[15]), .B2(n388), .C1(S2[15]), 
        .C2(n385), .ZN(n54) );
  INV_X1 U50 ( .A(n53), .ZN(Y[16]) );
  AOI222_X1 U51 ( .A1(S0[16]), .A2(n391), .B1(S1[16]), .B2(n388), .C1(S2[16]), 
        .C2(n385), .ZN(n53) );
  INV_X1 U52 ( .A(n52), .ZN(Y[17]) );
  AOI222_X1 U53 ( .A1(S0[17]), .A2(n391), .B1(S1[17]), .B2(n388), .C1(S2[17]), 
        .C2(n385), .ZN(n52) );
  INV_X1 U54 ( .A(n51), .ZN(Y[18]) );
  AOI222_X1 U55 ( .A1(S0[18]), .A2(n391), .B1(S1[18]), .B2(n388), .C1(S2[18]), 
        .C2(n385), .ZN(n51) );
  INV_X1 U56 ( .A(n50), .ZN(Y[19]) );
  AOI222_X1 U57 ( .A1(S0[19]), .A2(n391), .B1(S1[19]), .B2(n388), .C1(S2[19]), 
        .C2(n385), .ZN(n50) );
  INV_X1 U58 ( .A(n49), .ZN(Y[20]) );
  AOI222_X1 U59 ( .A1(S0[20]), .A2(n391), .B1(S1[20]), .B2(n388), .C1(S2[20]), 
        .C2(n385), .ZN(n49) );
  INV_X1 U60 ( .A(n48), .ZN(Y[21]) );
  AOI222_X1 U61 ( .A1(S0[21]), .A2(n391), .B1(S1[21]), .B2(n388), .C1(S2[21]), 
        .C2(n385), .ZN(n48) );
  INV_X1 U62 ( .A(n47), .ZN(Y[22]) );
  AOI222_X1 U63 ( .A1(S0[22]), .A2(n392), .B1(S1[22]), .B2(n388), .C1(S2[22]), 
        .C2(n385), .ZN(n47) );
  INV_X1 U64 ( .A(n46), .ZN(Y[23]) );
  AOI222_X1 U65 ( .A1(S0[23]), .A2(n392), .B1(S1[23]), .B2(n388), .C1(S2[23]), 
        .C2(n385), .ZN(n46) );
  INV_X1 U66 ( .A(n45), .ZN(Y[24]) );
  AOI222_X1 U67 ( .A1(S0[24]), .A2(n392), .B1(S1[24]), .B2(n389), .C1(S2[24]), 
        .C2(n386), .ZN(n45) );
  INV_X1 U68 ( .A(n44), .ZN(Y[25]) );
  AOI222_X1 U69 ( .A1(S0[25]), .A2(n392), .B1(S1[25]), .B2(n389), .C1(S2[25]), 
        .C2(n386), .ZN(n44) );
  INV_X1 U70 ( .A(n43), .ZN(Y[26]) );
  AOI222_X1 U71 ( .A1(S0[26]), .A2(n392), .B1(S1[26]), .B2(n389), .C1(S2[26]), 
        .C2(n386), .ZN(n43) );
  INV_X1 U72 ( .A(n42), .ZN(Y[27]) );
  AOI222_X1 U73 ( .A1(S0[27]), .A2(n392), .B1(S1[27]), .B2(n389), .C1(S2[27]), 
        .C2(n386), .ZN(n42) );
  INV_X1 U74 ( .A(n41), .ZN(Y[28]) );
  AOI222_X1 U75 ( .A1(S0[28]), .A2(n392), .B1(S1[28]), .B2(n389), .C1(S2[28]), 
        .C2(n386), .ZN(n41) );
  INV_X1 U76 ( .A(n40), .ZN(Y[29]) );
  AOI222_X1 U77 ( .A1(S0[29]), .A2(n392), .B1(S1[29]), .B2(n389), .C1(S2[29]), 
        .C2(n386), .ZN(n40) );
  INV_X1 U78 ( .A(n39), .ZN(Y[30]) );
  AOI222_X1 U79 ( .A1(S0[30]), .A2(n392), .B1(S1[30]), .B2(n389), .C1(S2[30]), 
        .C2(n386), .ZN(n39) );
endmodule


module PG_NETWORK_WIDTH32 ( A, B, Ci, P, G );
  input [31:0] A;
  input [31:0] B;
  output [31:0] P;
  output [31:0] G;
  input Ci;
  wire   n3, n4, n14;

  XOR2_X1 U36 ( .A(B[9]), .B(A[9]), .Z(P[9]) );
  XOR2_X1 U37 ( .A(B[8]), .B(A[8]), .Z(P[8]) );
  XOR2_X1 U38 ( .A(B[7]), .B(A[7]), .Z(P[7]) );
  XOR2_X1 U39 ( .A(B[6]), .B(A[6]), .Z(P[6]) );
  XOR2_X1 U40 ( .A(B[5]), .B(A[5]), .Z(P[5]) );
  XOR2_X1 U41 ( .A(B[4]), .B(A[4]), .Z(P[4]) );
  XOR2_X1 U42 ( .A(B[3]), .B(A[3]), .Z(P[3]) );
  XOR2_X1 U43 ( .A(B[31]), .B(A[31]), .Z(P[31]) );
  XOR2_X1 U44 ( .A(B[30]), .B(A[30]), .Z(P[30]) );
  XOR2_X1 U45 ( .A(B[2]), .B(A[2]), .Z(P[2]) );
  XOR2_X1 U46 ( .A(B[29]), .B(A[29]), .Z(P[29]) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(P[28]) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(P[27]) );
  XOR2_X1 U49 ( .A(B[26]), .B(A[26]), .Z(P[26]) );
  XOR2_X1 U50 ( .A(B[25]), .B(A[25]), .Z(P[25]) );
  XOR2_X1 U51 ( .A(B[24]), .B(A[24]), .Z(P[24]) );
  XOR2_X1 U52 ( .A(B[23]), .B(A[23]), .Z(P[23]) );
  XOR2_X1 U53 ( .A(B[22]), .B(A[22]), .Z(P[22]) );
  XOR2_X1 U54 ( .A(B[21]), .B(A[21]), .Z(P[21]) );
  XOR2_X1 U55 ( .A(B[20]), .B(A[20]), .Z(P[20]) );
  XOR2_X1 U56 ( .A(B[1]), .B(A[1]), .Z(P[1]) );
  XOR2_X1 U57 ( .A(B[19]), .B(A[19]), .Z(P[19]) );
  XOR2_X1 U58 ( .A(B[18]), .B(A[18]), .Z(P[18]) );
  XOR2_X1 U59 ( .A(B[17]), .B(A[17]), .Z(P[17]) );
  XOR2_X1 U60 ( .A(B[16]), .B(A[16]), .Z(P[16]) );
  XOR2_X1 U61 ( .A(B[15]), .B(A[15]), .Z(P[15]) );
  XOR2_X1 U62 ( .A(B[14]), .B(A[14]), .Z(P[14]) );
  XOR2_X1 U63 ( .A(B[13]), .B(A[13]), .Z(P[13]) );
  XOR2_X1 U64 ( .A(B[12]), .B(A[12]), .Z(P[12]) );
  XOR2_X1 U65 ( .A(B[11]), .B(A[11]), .Z(P[11]) );
  XOR2_X1 U66 ( .A(B[10]), .B(A[10]), .Z(P[10]) );
  XOR2_X1 U67 ( .A(B[0]), .B(A[0]), .Z(P[0]) );
  AND2_X1 U1 ( .A1(B[18]), .A2(A[18]), .ZN(G[18]) );
  AND2_X1 U2 ( .A1(B[19]), .A2(A[19]), .ZN(G[19]) );
  AND2_X1 U3 ( .A1(B[16]), .A2(A[16]), .ZN(G[16]) );
  AND2_X1 U4 ( .A1(B[17]), .A2(A[17]), .ZN(G[17]) );
  AND2_X1 U5 ( .A1(B[10]), .A2(A[10]), .ZN(G[10]) );
  AND2_X1 U6 ( .A1(B[11]), .A2(A[11]), .ZN(G[11]) );
  AND2_X1 U7 ( .A1(B[8]), .A2(A[8]), .ZN(G[8]) );
  AND2_X1 U8 ( .A1(B[9]), .A2(A[9]), .ZN(G[9]) );
  AND2_X1 U9 ( .A1(B[12]), .A2(A[12]), .ZN(G[12]) );
  AND2_X1 U10 ( .A1(B[13]), .A2(A[13]), .ZN(G[13]) );
  AND2_X1 U11 ( .A1(B[26]), .A2(A[26]), .ZN(G[26]) );
  AND2_X1 U12 ( .A1(B[27]), .A2(A[27]), .ZN(G[27]) );
  AND2_X1 U13 ( .A1(B[24]), .A2(A[24]), .ZN(G[24]) );
  AND2_X1 U14 ( .A1(B[25]), .A2(A[25]), .ZN(G[25]) );
  AND2_X1 U15 ( .A1(B[30]), .A2(A[30]), .ZN(G[30]) );
  AND2_X1 U16 ( .A1(B[31]), .A2(A[31]), .ZN(G[31]) );
  AND2_X1 U17 ( .A1(B[6]), .A2(A[6]), .ZN(G[6]) );
  AND2_X1 U18 ( .A1(B[7]), .A2(A[7]), .ZN(G[7]) );
  AND2_X1 U19 ( .A1(B[2]), .A2(A[2]), .ZN(G[2]) );
  AND2_X1 U20 ( .A1(B[3]), .A2(A[3]), .ZN(G[3]) );
  INV_X1 U21 ( .A(n3), .ZN(G[0]) );
  AND2_X1 U22 ( .A1(B[1]), .A2(A[1]), .ZN(G[1]) );
  AOI21_X1 U23 ( .B1(A[0]), .B2(B[0]), .A(n14), .ZN(n3) );
  INV_X1 U24 ( .A(n4), .ZN(n14) );
  OAI21_X1 U25 ( .B1(A[0]), .B2(B[0]), .A(Ci), .ZN(n4) );
  AND2_X1 U26 ( .A1(B[29]), .A2(A[29]), .ZN(G[29]) );
  AND2_X1 U27 ( .A1(B[5]), .A2(A[5]), .ZN(G[5]) );
  AND2_X1 U28 ( .A1(B[28]), .A2(A[28]), .ZN(G[28]) );
  AND2_X1 U29 ( .A1(B[4]), .A2(A[4]), .ZN(G[4]) );
  AND2_X1 U30 ( .A1(B[22]), .A2(A[22]), .ZN(G[22]) );
  AND2_X1 U31 ( .A1(B[23]), .A2(A[23]), .ZN(G[23]) );
  AND2_X1 U32 ( .A1(B[14]), .A2(A[14]), .ZN(G[14]) );
  AND2_X1 U33 ( .A1(B[15]), .A2(A[15]), .ZN(G[15]) );
  AND2_X1 U34 ( .A1(B[20]), .A2(A[20]), .ZN(G[20]) );
  AND2_X1 U35 ( .A1(B[21]), .A2(A[21]), .ZN(G[21]) );
endmodule


module BLOCKPG_0 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n2) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_28 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_27 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_26 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_25 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_24 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_23 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_22 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n2;

  AND2_X1 U1 ( .A1(pik_1), .A2(pik), .ZN(pij) );
  INV_X1 U2 ( .A(n2), .ZN(gij) );
  AOI21_X1 U3 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n2) );
endmodule


module BLOCKPG_21 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_20 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_19 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  AND2_X1 U1 ( .A1(pik_1), .A2(pik), .ZN(pij) );
  INV_X1 U2 ( .A(n12), .ZN(gij) );
  AOI21_X1 U3 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
endmodule


module BLOCKPG_18 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  AND2_X1 U1 ( .A1(pik_1), .A2(pik), .ZN(pij) );
  INV_X1 U2 ( .A(n12), .ZN(gij) );
  AOI21_X1 U3 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
endmodule


module BLOCKPG_17 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_16 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_15 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_14 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_13 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_12 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gij) );
  AND2_X1 U2 ( .A1(pik_1), .A2(pik), .ZN(pij) );
  AOI21_X1 U3 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n2) );
endmodule


module BLOCKPG_11 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_10 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_9 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_8 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_7 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_6 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n2;

  AOI21_X1 U1 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(gij) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKG_0 ( pik, gik, pik_1, gik_1, gij );
  input pik, gik, pik_1, gik_1;
  output gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(gij) );
  AOI21_X1 U2 ( .B1(pik), .B2(gik_1), .A(gik), .ZN(n2) );
endmodule


module BLOCKPG_5 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AND2_X1 U2 ( .A1(pik_1), .A2(pik), .ZN(pij) );
  AOI21_X1 U3 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
endmodule


module BLOCKPG_4 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKPG_3 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
  AND2_X1 U3 ( .A1(pik_1), .A2(pik), .ZN(pij) );
endmodule


module BLOCKG_6 ( pik, gik, pik_1, gik_1, gij );
  input pik, gik, pik_1, gik_1;
  output gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(pik), .B2(gik_1), .A(gik), .ZN(n12) );
endmodule


module BLOCKG_5 ( pik, gik, pik_1, gik_1, gij );
  input pik, gik, pik_1, gik_1;
  output gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(pik), .B2(gik_1), .A(gik), .ZN(n12) );
endmodule


module BLOCKPG_2 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AND2_X1 U2 ( .A1(pik_1), .A2(pik), .ZN(pij) );
  AOI21_X1 U3 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n12) );
endmodule


module BLOCKPG_1 ( pik, gik, pik_1, gik_1, pij, gij );
  input pik, gik, pik_1, gik_1;
  output pij, gij;
  wire   n2;

  AND2_X1 U1 ( .A1(pik_1), .A2(pik), .ZN(pij) );
  AOI21_X1 U2 ( .B1(gik_1), .B2(pik), .A(gik), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(gij) );
endmodule


module BLOCKG_4 ( pik, gik, pik_1, gik_1, gij );
  input pik, gik, pik_1, gik_1;
  output gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(pik), .B2(gik_1), .A(gik), .ZN(n12) );
endmodule


module BLOCKG_3 ( pik, gik, pik_1, gik_1, gij );
  input pik, gik, pik_1, gik_1;
  output gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(pik), .B2(gik_1), .A(gik), .ZN(n12) );
endmodule


module BLOCKG_2 ( pik, gik, pik_1, gik_1, gij );
  input pik, gik, pik_1, gik_1;
  output gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(pik), .B2(gik_1), .A(gik), .ZN(n12) );
endmodule


module BLOCKG_1 ( pik, gik, pik_1, gik_1, gij );
  input pik, gik, pik_1, gik_1;
  output gij;
  wire   n12;

  INV_X1 U1 ( .A(n12), .ZN(gij) );
  AOI21_X1 U2 ( .B1(pik), .B2(gik_1), .A(gik), .ZN(n12) );
endmodule


module SPARSE_TREE_WIDTH32_RADIX4 ( A, B, Ci, Co );
  input [31:0] A;
  input [31:0] B;
  output [8:0] Co;
  input Ci;
  wire   Ci, \s_G[5][31] , \s_G[5][30] , \s_G[5][29] , \s_G[5][28] ,
         \s_G[5][27] , \s_G[5][26] , \s_G[5][25] , \s_G[5][24] , \s_G[5][23] ,
         \s_G[5][22] , \s_G[5][21] , \s_G[5][20] , \s_G[5][19] , \s_G[5][18] ,
         \s_G[5][17] , \s_G[5][16] , \s_G[5][15] , \s_G[5][14] , \s_G[5][13] ,
         \s_G[5][12] , \s_G[5][11] , \s_G[5][10] , \s_G[5][9] , \s_G[5][8] ,
         \s_G[5][7] , \s_G[5][6] , \s_G[5][5] , \s_G[5][4] , \s_G[5][3] ,
         \s_G[5][2] , \s_G[5][1] , \s_G[5][0] , \s_G[4][15] , \s_G[4][14] ,
         \s_G[4][13] , \s_G[4][12] , \s_G[4][11] , \s_G[4][10] , \s_G[4][9] ,
         \s_G[4][8] , \s_G[4][7] , \s_G[4][6] , \s_G[4][5] , \s_G[4][4] ,
         \s_G[4][3] , \s_G[4][2] , \s_G[4][1] , \s_G[4][0] , \s_G[3][7] ,
         \s_G[3][6] , \s_G[3][5] , \s_G[3][4] , \s_G[3][3] , \s_G[3][2] ,
         \s_G[3][1] , \s_G[2][7] , \s_G[2][5] , \s_G[2][3] , \s_G[1][7] ,
         \s_G[1][6] , \s_P[5][31] , \s_P[5][30] , \s_P[5][29] , \s_P[5][28] ,
         \s_P[5][27] , \s_P[5][26] , \s_P[5][25] , \s_P[5][24] , \s_P[5][23] ,
         \s_P[5][22] , \s_P[5][21] , \s_P[5][20] , \s_P[5][19] , \s_P[5][18] ,
         \s_P[5][17] , \s_P[5][16] , \s_P[5][15] , \s_P[5][14] , \s_P[5][13] ,
         \s_P[5][12] , \s_P[5][11] , \s_P[5][10] , \s_P[5][9] , \s_P[5][8] ,
         \s_P[5][7] , \s_P[5][6] , \s_P[5][5] , \s_P[5][4] , \s_P[5][3] ,
         \s_P[5][2] , \s_P[5][1] , \s_P[5][0] , \s_P[4][15] , \s_P[4][14] ,
         \s_P[4][13] , \s_P[4][12] , \s_P[4][11] , \s_P[4][10] , \s_P[4][9] ,
         \s_P[4][8] , \s_P[4][7] , \s_P[4][6] , \s_P[4][5] , \s_P[4][4] ,
         \s_P[4][3] , \s_P[4][2] , \s_P[4][1] , \s_P[4][0] , \s_P[3][7] ,
         \s_P[3][6] , \s_P[3][5] , \s_P[3][4] , \s_P[3][3] , \s_P[3][2] ,
         \s_P[3][1] , \s_P[3][0] , \s_P[2][7] , \s_P[2][5] , \s_P[2][3] ,
         \s_P[1][7] , \s_P[1][6] ;
  assign Co[0] = Ci;

  PG_NETWORK_WIDTH32 PGNET ( .A(A), .B(B), .Ci(Ci), .P({\s_P[5][31] , 
        \s_P[5][30] , \s_P[5][29] , \s_P[5][28] , \s_P[5][27] , \s_P[5][26] , 
        \s_P[5][25] , \s_P[5][24] , \s_P[5][23] , \s_P[5][22] , \s_P[5][21] , 
        \s_P[5][20] , \s_P[5][19] , \s_P[5][18] , \s_P[5][17] , \s_P[5][16] , 
        \s_P[5][15] , \s_P[5][14] , \s_P[5][13] , \s_P[5][12] , \s_P[5][11] , 
        \s_P[5][10] , \s_P[5][9] , \s_P[5][8] , \s_P[5][7] , \s_P[5][6] , 
        \s_P[5][5] , \s_P[5][4] , \s_P[5][3] , \s_P[5][2] , \s_P[5][1] , 
        \s_P[5][0] }), .G({\s_G[5][31] , \s_G[5][30] , \s_G[5][29] , 
        \s_G[5][28] , \s_G[5][27] , \s_G[5][26] , \s_G[5][25] , \s_G[5][24] , 
        \s_G[5][23] , \s_G[5][22] , \s_G[5][21] , \s_G[5][20] , \s_G[5][19] , 
        \s_G[5][18] , \s_G[5][17] , \s_G[5][16] , \s_G[5][15] , \s_G[5][14] , 
        \s_G[5][13] , \s_G[5][12] , \s_G[5][11] , \s_G[5][10] , \s_G[5][9] , 
        \s_G[5][8] , \s_G[5][7] , \s_G[5][6] , \s_G[5][5] , \s_G[5][4] , 
        \s_G[5][3] , \s_G[5][2] , \s_G[5][1] , \s_G[5][0] }) );
  BLOCKPG_0 PGij_5_0 ( .pik(\s_P[5][1] ), .gik(\s_G[5][1] ), .pik_1(
        \s_P[5][0] ), .gik_1(\s_G[5][0] ), .pij(\s_P[4][0] ), .gij(\s_G[4][0] ) );
  BLOCKPG_28 PGij_5_1 ( .pik(\s_P[5][3] ), .gik(\s_G[5][3] ), .pik_1(
        \s_P[5][2] ), .gik_1(\s_G[5][2] ), .pij(\s_P[4][1] ), .gij(\s_G[4][1] ) );
  BLOCKPG_27 PGij_5_2 ( .pik(\s_P[5][5] ), .gik(\s_G[5][5] ), .pik_1(
        \s_P[5][4] ), .gik_1(\s_G[5][4] ), .pij(\s_P[4][2] ), .gij(\s_G[4][2] ) );
  BLOCKPG_26 PGij_5_3 ( .pik(\s_P[5][7] ), .gik(\s_G[5][7] ), .pik_1(
        \s_P[5][6] ), .gik_1(\s_G[5][6] ), .pij(\s_P[4][3] ), .gij(\s_G[4][3] ) );
  BLOCKPG_25 PGij_5_4 ( .pik(\s_P[5][9] ), .gik(\s_G[5][9] ), .pik_1(
        \s_P[5][8] ), .gik_1(\s_G[5][8] ), .pij(\s_P[4][4] ), .gij(\s_G[4][4] ) );
  BLOCKPG_24 PGij_5_5 ( .pik(\s_P[5][11] ), .gik(\s_G[5][11] ), .pik_1(
        \s_P[5][10] ), .gik_1(\s_G[5][10] ), .pij(\s_P[4][5] ), .gij(
        \s_G[4][5] ) );
  BLOCKPG_23 PGij_5_6 ( .pik(\s_P[5][13] ), .gik(\s_G[5][13] ), .pik_1(
        \s_P[5][12] ), .gik_1(\s_G[5][12] ), .pij(\s_P[4][6] ), .gij(
        \s_G[4][6] ) );
  BLOCKPG_22 PGij_5_7 ( .pik(\s_P[5][15] ), .gik(\s_G[5][15] ), .pik_1(
        \s_P[5][14] ), .gik_1(\s_G[5][14] ), .pij(\s_P[4][7] ), .gij(
        \s_G[4][7] ) );
  BLOCKPG_21 PGij_5_8 ( .pik(\s_P[5][17] ), .gik(\s_G[5][17] ), .pik_1(
        \s_P[5][16] ), .gik_1(\s_G[5][16] ), .pij(\s_P[4][8] ), .gij(
        \s_G[4][8] ) );
  BLOCKPG_20 PGij_5_9 ( .pik(\s_P[5][19] ), .gik(\s_G[5][19] ), .pik_1(
        \s_P[5][18] ), .gik_1(\s_G[5][18] ), .pij(\s_P[4][9] ), .gij(
        \s_G[4][9] ) );
  BLOCKPG_19 PGij_5_10 ( .pik(\s_P[5][21] ), .gik(\s_G[5][21] ), .pik_1(
        \s_P[5][20] ), .gik_1(\s_G[5][20] ), .pij(\s_P[4][10] ), .gij(
        \s_G[4][10] ) );
  BLOCKPG_18 PGij_5_11 ( .pik(\s_P[5][23] ), .gik(\s_G[5][23] ), .pik_1(
        \s_P[5][22] ), .gik_1(\s_G[5][22] ), .pij(\s_P[4][11] ), .gij(
        \s_G[4][11] ) );
  BLOCKPG_17 PGij_5_12 ( .pik(\s_P[5][25] ), .gik(\s_G[5][25] ), .pik_1(
        \s_P[5][24] ), .gik_1(\s_G[5][24] ), .pij(\s_P[4][12] ), .gij(
        \s_G[4][12] ) );
  BLOCKPG_16 PGij_5_13 ( .pik(\s_P[5][27] ), .gik(\s_G[5][27] ), .pik_1(
        \s_P[5][26] ), .gik_1(\s_G[5][26] ), .pij(\s_P[4][13] ), .gij(
        \s_G[4][13] ) );
  BLOCKPG_15 PGij_5_14 ( .pik(\s_P[5][29] ), .gik(\s_G[5][29] ), .pik_1(
        \s_P[5][28] ), .gik_1(\s_G[5][28] ), .pij(\s_P[4][14] ), .gij(
        \s_G[4][14] ) );
  BLOCKPG_14 PGij_5_15 ( .pik(\s_P[5][31] ), .gik(\s_G[5][31] ), .pik_1(
        \s_P[5][30] ), .gik_1(\s_G[5][30] ), .pij(\s_P[4][15] ), .gij(
        \s_G[4][15] ) );
  BLOCKPG_13 PGij_4_0 ( .pik(\s_P[4][1] ), .gik(\s_G[4][1] ), .pik_1(
        \s_P[4][0] ), .gik_1(\s_G[4][0] ), .pij(\s_P[3][0] ), .gij(Co[1]) );
  BLOCKPG_12 PGij_4_1 ( .pik(\s_P[4][3] ), .gik(\s_G[4][3] ), .pik_1(
        \s_P[4][2] ), .gik_1(\s_G[4][2] ), .pij(\s_P[3][1] ), .gij(\s_G[3][1] ) );
  BLOCKPG_11 PGij_4_2 ( .pik(\s_P[4][5] ), .gik(\s_G[4][5] ), .pik_1(
        \s_P[4][4] ), .gik_1(\s_G[4][4] ), .pij(\s_P[3][2] ), .gij(\s_G[3][2] ) );
  BLOCKPG_10 PGij_4_3 ( .pik(\s_P[4][7] ), .gik(\s_G[4][7] ), .pik_1(
        \s_P[4][6] ), .gik_1(\s_G[4][6] ), .pij(\s_P[3][3] ), .gij(\s_G[3][3] ) );
  BLOCKPG_9 PGij_4_4 ( .pik(\s_P[4][9] ), .gik(\s_G[4][9] ), .pik_1(
        \s_P[4][8] ), .gik_1(\s_G[4][8] ), .pij(\s_P[3][4] ), .gij(\s_G[3][4] ) );
  BLOCKPG_8 PGij_4_5 ( .pik(\s_P[4][11] ), .gik(\s_G[4][11] ), .pik_1(
        \s_P[4][10] ), .gik_1(\s_G[4][10] ), .pij(\s_P[3][5] ), .gij(
        \s_G[3][5] ) );
  BLOCKPG_7 PGij_4_6 ( .pik(\s_P[4][13] ), .gik(\s_G[4][13] ), .pik_1(
        \s_P[4][12] ), .gik_1(\s_G[4][12] ), .pij(\s_P[3][6] ), .gij(
        \s_G[3][6] ) );
  BLOCKPG_6 PGij_4_7 ( .pik(\s_P[4][15] ), .gik(\s_G[4][15] ), .pik_1(
        \s_P[4][14] ), .gik_1(\s_G[4][14] ), .pij(\s_P[3][7] ), .gij(
        \s_G[3][7] ) );
  BLOCKG_0 G_GEN_3_0_0 ( .pik(\s_P[3][1] ), .gik(\s_G[3][1] ), .pik_1(
        \s_P[3][0] ), .gik_1(Co[1]), .gij(Co[2]) );
  BLOCKPG_5 PG_GEN_3_1_0 ( .pik(\s_P[3][3] ), .gik(\s_G[3][3] ), .pik_1(
        \s_P[3][2] ), .gik_1(\s_G[3][2] ), .pij(\s_P[2][3] ), .gij(\s_G[2][3] ) );
  BLOCKPG_4 PG_GEN_3_2_0 ( .pik(\s_P[3][5] ), .gik(\s_G[3][5] ), .pik_1(
        \s_P[3][4] ), .gik_1(\s_G[3][4] ), .pij(\s_P[2][5] ), .gij(\s_G[2][5] ) );
  BLOCKPG_3 PG_GEN_3_3_0 ( .pik(\s_P[3][7] ), .gik(\s_G[3][7] ), .pik_1(
        \s_P[3][6] ), .gik_1(\s_G[3][6] ), .pij(\s_P[2][7] ), .gij(\s_G[2][7] ) );
  BLOCKG_6 G_GEN_2_0_0 ( .pik(\s_P[3][2] ), .gik(\s_G[3][2] ), .pik_1(1'b0), 
        .gik_1(Co[2]), .gij(Co[3]) );
  BLOCKG_5 G_GEN_2_0_1 ( .pik(\s_P[2][3] ), .gik(\s_G[2][3] ), .pik_1(1'b0), 
        .gik_1(Co[2]), .gij(Co[4]) );
  BLOCKPG_2 PG_GEN_2_1_0 ( .pik(\s_P[3][6] ), .gik(\s_G[3][6] ), .pik_1(
        \s_P[2][5] ), .gik_1(\s_G[2][5] ), .pij(\s_P[1][6] ), .gij(\s_G[1][6] ) );
  BLOCKPG_1 PG_GEN_2_1_1 ( .pik(\s_P[2][7] ), .gik(\s_G[2][7] ), .pik_1(
        \s_P[2][5] ), .gik_1(\s_G[2][5] ), .pij(\s_P[1][7] ), .gij(\s_G[1][7] ) );
  BLOCKG_4 G_GEN_1_0_0 ( .pik(\s_P[3][4] ), .gik(\s_G[3][4] ), .pik_1(1'b0), 
        .gik_1(Co[4]), .gij(Co[5]) );
  BLOCKG_3 G_GEN_1_0_1 ( .pik(\s_P[2][5] ), .gik(\s_G[2][5] ), .pik_1(1'b0), 
        .gik_1(Co[4]), .gij(Co[6]) );
  BLOCKG_2 G_GEN_1_0_2 ( .pik(\s_P[1][6] ), .gik(\s_G[1][6] ), .pik_1(1'b0), 
        .gik_1(Co[4]), .gij(Co[7]) );
  BLOCKG_1 G_GEN_1_0_3 ( .pik(\s_P[1][7] ), .gik(\s_G[1][7] ), .pik_1(1'b0), 
        .gik_1(Co[4]), .gij(Co[8]) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_64 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_0 ( S1, S0, SEL, Y );
  input [3:0] S1;
  input [3:0] S0;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n33;

  INV_X1 U1 ( .A(SEL), .ZN(n33) );
  INV_X1 U2 ( .A(n8), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(S0[1]), .A2(n33), .B1(S1[1]), .B2(SEL), .ZN(n8) );
  INV_X1 U4 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(S0[3]), .A2(n33), .B1(SEL), .B2(S1[3]), .ZN(n6) );
  INV_X1 U6 ( .A(n7), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(S0[2]), .A2(n33), .B1(S1[2]), .B2(SEL), .ZN(n7) );
  INV_X1 U8 ( .A(n9), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(S0[0]), .A2(n33), .B1(S1[0]), .B2(SEL), .ZN(n9) );
endmodule


module CSB_RADIX4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_WIDTH4_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_WIDTH4_15 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  MUX21_GENERIC_NBIT4_0 MUX21_SUM ( .S1(S1), .S0(S0), .SEL(Ci), .Y(S) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_7 ( S1, S0, SEL, Y );
  input [3:0] S1;
  input [3:0] S0;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n49;

  INV_X1 U1 ( .A(SEL), .ZN(n49) );
  INV_X1 U2 ( .A(n8), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(S0[1]), .A2(n49), .B1(S1[1]), .B2(SEL), .ZN(n8) );
  INV_X1 U4 ( .A(n7), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(S0[2]), .A2(n49), .B1(S1[2]), .B2(SEL), .ZN(n7) );
  INV_X1 U6 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(S0[3]), .A2(n49), .B1(SEL), .B2(S1[3]), .ZN(n6) );
  INV_X1 U8 ( .A(n9), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(S0[0]), .A2(n49), .B1(S1[0]), .B2(SEL), .ZN(n9) );
endmodule


module CSB_RADIX4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_WIDTH4_14 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_WIDTH4_13 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  MUX21_GENERIC_NBIT4_7 MUX21_SUM ( .S1(S1), .S0(S0), .SEL(Ci), .Y(S) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_6 ( S1, S0, SEL, Y );
  input [3:0] S1;
  input [3:0] S0;
  output [3:0] Y;
  input SEL;
  wire   n49, n50, n51, n52, n53;

  INV_X1 U1 ( .A(SEL), .ZN(n49) );
  INV_X1 U2 ( .A(n51), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(S0[1]), .A2(n49), .B1(S1[1]), .B2(SEL), .ZN(n51) );
  INV_X1 U4 ( .A(n52), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(S0[2]), .A2(n49), .B1(S1[2]), .B2(SEL), .ZN(n52) );
  INV_X1 U6 ( .A(n53), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(S0[3]), .A2(n49), .B1(SEL), .B2(S1[3]), .ZN(n53) );
  INV_X1 U8 ( .A(n50), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(S0[0]), .A2(n49), .B1(S1[0]), .B2(SEL), .ZN(n50) );
endmodule


module CSB_RADIX4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_WIDTH4_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_WIDTH4_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  MUX21_GENERIC_NBIT4_6 MUX21_SUM ( .S1(S1), .S0(S0), .SEL(Ci), .Y(S) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_5 ( S1, S0, SEL, Y );
  input [3:0] S1;
  input [3:0] S0;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n37;

  INV_X1 U1 ( .A(SEL), .ZN(n37) );
  INV_X1 U2 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(S0[3]), .A2(n37), .B1(SEL), .B2(S1[3]), .ZN(n6) );
  INV_X1 U4 ( .A(n8), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(S0[1]), .A2(n37), .B1(S1[1]), .B2(SEL), .ZN(n8) );
  INV_X1 U6 ( .A(n7), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(S0[2]), .A2(n37), .B1(S1[2]), .B2(SEL), .ZN(n7) );
  INV_X1 U8 ( .A(n9), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(S0[0]), .A2(n37), .B1(S1[0]), .B2(SEL), .ZN(n9) );
endmodule


module CSB_RADIX4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_WIDTH4_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_WIDTH4_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  MUX21_GENERIC_NBIT4_5 MUX21_SUM ( .S1(S1), .S0(S0), .SEL(Ci), .Y(S) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_4 ( S1, S0, SEL, Y );
  input [3:0] S1;
  input [3:0] S0;
  output [3:0] Y;
  input SEL;
  wire   n49, n50, n51, n52, n53;

  INV_X1 U1 ( .A(SEL), .ZN(n49) );
  INV_X1 U2 ( .A(n51), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(S0[1]), .A2(n49), .B1(S1[1]), .B2(SEL), .ZN(n51) );
  INV_X1 U4 ( .A(n52), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(S0[2]), .A2(n49), .B1(S1[2]), .B2(SEL), .ZN(n52) );
  INV_X1 U6 ( .A(n53), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(S0[3]), .A2(n49), .B1(SEL), .B2(S1[3]), .ZN(n53) );
  INV_X1 U8 ( .A(n50), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(S0[0]), .A2(n49), .B1(S1[0]), .B2(SEL), .ZN(n50) );
endmodule


module CSB_RADIX4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_WIDTH4_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_WIDTH4_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  MUX21_GENERIC_NBIT4_4 MUX21_SUM ( .S1(S1), .S0(S0), .SEL(Ci), .Y(S) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_3 ( S1, S0, SEL, Y );
  input [3:0] S1;
  input [3:0] S0;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n37;

  INV_X1 U1 ( .A(SEL), .ZN(n37) );
  INV_X1 U2 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(S0[3]), .A2(n37), .B1(SEL), .B2(S1[3]), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(S0[2]), .A2(n37), .B1(S1[2]), .B2(SEL), .ZN(n7) );
  INV_X1 U6 ( .A(n8), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(S0[1]), .A2(n37), .B1(S1[1]), .B2(SEL), .ZN(n8) );
  INV_X1 U8 ( .A(n9), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(S0[0]), .A2(n37), .B1(S1[0]), .B2(SEL), .ZN(n9) );
endmodule


module CSB_RADIX4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_WIDTH4_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_WIDTH4_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  MUX21_GENERIC_NBIT4_3 MUX21_SUM ( .S1(S1), .S0(S0), .SEL(Ci), .Y(S) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_2 ( S1, S0, SEL, Y );
  input [3:0] S1;
  input [3:0] S0;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n37;

  INV_X1 U1 ( .A(SEL), .ZN(n37) );
  INV_X1 U2 ( .A(n7), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(S0[2]), .A2(n37), .B1(S1[2]), .B2(SEL), .ZN(n7) );
  INV_X1 U4 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(S0[3]), .A2(n37), .B1(SEL), .B2(S1[3]), .ZN(n6) );
  INV_X1 U6 ( .A(n8), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(S0[1]), .A2(n37), .B1(S1[1]), .B2(SEL), .ZN(n8) );
  INV_X1 U8 ( .A(n9), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(S0[0]), .A2(n37), .B1(S1[0]), .B2(SEL), .ZN(n9) );
endmodule


module CSB_RADIX4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_WIDTH4_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_WIDTH4_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  MUX21_GENERIC_NBIT4_2 MUX21_SUM ( .S1(S1), .S0(S0), .SEL(Ci), .Y(S) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_WIDTH4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FA_i_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_1 ( S1, S0, SEL, Y );
  input [3:0] S1;
  input [3:0] S0;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n33;

  INV_X1 U1 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U2 ( .A1(S0[3]), .A2(n33), .B1(SEL), .B2(S1[3]), .ZN(n6) );
  INV_X1 U3 ( .A(n7), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(S0[2]), .A2(n33), .B1(S1[2]), .B2(SEL), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(S0[1]), .A2(n33), .B1(S1[1]), .B2(SEL), .ZN(n8) );
  INV_X1 U7 ( .A(n9), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(S0[0]), .A2(n33), .B1(S1[0]), .B2(SEL), .ZN(n9) );
  INV_X1 U9 ( .A(SEL), .ZN(n33) );
endmodule


module CSB_RADIX4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_WIDTH4_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_WIDTH4_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  MUX21_GENERIC_NBIT4_1 MUX21_SUM ( .S1(S1), .S0(S0), .SEL(Ci), .Y(S) );
endmodule


module SUM_GENERATOR_WIDTH32_RADIX4 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  CSB_RADIX4_0 CSBi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(S[31:28])
         );
  CSB_RADIX4_7 CSBi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(S[27:24])
         );
  CSB_RADIX4_6 CSBi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(S[23:20])
         );
  CSB_RADIX4_5 CSBi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(S[19:16])
         );
  CSB_RADIX4_4 CSBi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(S[15:12])
         );
  CSB_RADIX4_3 CSBi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  CSB_RADIX4_2 CSBi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  CSB_RADIX4_1 CSBi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
endmodule


module ADDER_SUBTRACTOR_WIDTH32_RADIX4 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;
  wire   n5;
  wire   [31:0] s_B;
  wire   [7:0] carry_ST;

  XOR2_X1 U1 ( .A(n5), .B(B[9]), .Z(s_B[9]) );
  XOR2_X1 U2 ( .A(n5), .B(B[8]), .Z(s_B[8]) );
  XOR2_X1 U3 ( .A(n5), .B(B[7]), .Z(s_B[7]) );
  XOR2_X1 U4 ( .A(n5), .B(B[6]), .Z(s_B[6]) );
  XOR2_X1 U5 ( .A(n5), .B(B[5]), .Z(s_B[5]) );
  XOR2_X1 U6 ( .A(n5), .B(B[4]), .Z(s_B[4]) );
  XOR2_X1 U7 ( .A(n5), .B(B[3]), .Z(s_B[3]) );
  XOR2_X1 U8 ( .A(n5), .B(B[31]), .Z(s_B[31]) );
  XOR2_X1 U9 ( .A(n5), .B(B[30]), .Z(s_B[30]) );
  XOR2_X1 U10 ( .A(n5), .B(B[2]), .Z(s_B[2]) );
  XOR2_X1 U11 ( .A(n5), .B(B[29]), .Z(s_B[29]) );
  XOR2_X1 U12 ( .A(n5), .B(B[28]), .Z(s_B[28]) );
  XOR2_X1 U13 ( .A(n5), .B(B[27]), .Z(s_B[27]) );
  XOR2_X1 U14 ( .A(n5), .B(B[26]), .Z(s_B[26]) );
  XOR2_X1 U15 ( .A(n5), .B(B[25]), .Z(s_B[25]) );
  XOR2_X1 U16 ( .A(n5), .B(B[24]), .Z(s_B[24]) );
  XOR2_X1 U17 ( .A(n5), .B(B[23]), .Z(s_B[23]) );
  XOR2_X1 U18 ( .A(n5), .B(B[22]), .Z(s_B[22]) );
  XOR2_X1 U19 ( .A(n5), .B(B[21]), .Z(s_B[21]) );
  XOR2_X1 U20 ( .A(n5), .B(B[20]), .Z(s_B[20]) );
  XOR2_X1 U21 ( .A(n5), .B(B[1]), .Z(s_B[1]) );
  XOR2_X1 U22 ( .A(n5), .B(B[19]), .Z(s_B[19]) );
  XOR2_X1 U23 ( .A(n5), .B(B[18]), .Z(s_B[18]) );
  XOR2_X1 U24 ( .A(n5), .B(B[17]), .Z(s_B[17]) );
  XOR2_X1 U25 ( .A(n5), .B(B[16]), .Z(s_B[16]) );
  XOR2_X1 U26 ( .A(n5), .B(B[15]), .Z(s_B[15]) );
  XOR2_X1 U27 ( .A(n5), .B(B[14]), .Z(s_B[14]) );
  XOR2_X1 U28 ( .A(n5), .B(B[13]), .Z(s_B[13]) );
  XOR2_X1 U29 ( .A(n5), .B(B[12]), .Z(s_B[12]) );
  XOR2_X1 U30 ( .A(n5), .B(B[11]), .Z(s_B[11]) );
  XOR2_X1 U31 ( .A(n5), .B(B[10]), .Z(s_B[10]) );
  XOR2_X1 U32 ( .A(n5), .B(B[0]), .Z(s_B[0]) );
  SPARSE_TREE_WIDTH32_RADIX4 SPARSETREE ( .A(A), .B(s_B), .Ci(n5), .Co({Co, 
        carry_ST}) );
  SUM_GENERATOR_WIDTH32_RADIX4 SUMGEN ( .A(A), .B(s_B), .Ci(carry_ST), .S(S)
         );
  BUF_X2 U33 ( .A(Ci), .Z(n5) );
endmodule


module ZERO_DETECTOR_WIDTH32_1 ( A, Y );
  input [31:0] A;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NOR4_X1 U1 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n5) );
  NOR4_X1 U2 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n6) );
  NOR4_X1 U3 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n10) );
  NOR4_X1 U4 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n9) );
  NOR4_X1 U5 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n4) );
  NOR4_X1 U6 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n8) );
  NOR4_X1 U7 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n3) );
  NOR2_X1 U8 ( .A1(n1), .A2(n2), .ZN(Y) );
  NAND4_X1 U9 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
  NAND4_X1 U10 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NOR4_X1 U11 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n7) );
endmodule


module IVX_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_255 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_254 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_253 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_252 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_251 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_250 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_249 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_248 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_247 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_246 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_245 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_244 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_243 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_242 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_241 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_240 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_239 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_238 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_237 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_236 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_235 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_234 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_233 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_232 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_231 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_230 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_229 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_228 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_227 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_226 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_225 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_224 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_223 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_222 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_221 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_220 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_219 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_218 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_217 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_216 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_215 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_214 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_213 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_212 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_211 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_210 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_209 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_208 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_207 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_206 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_205 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_204 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_203 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_202 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_201 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_200 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_199 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_198 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_197 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_196 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_195 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_194 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_193 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_192 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_351 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_0 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_0 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_192 IVX_E ( .A(D), .Y(E) );
  NAND2_351 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_350 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_191 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_349 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_127 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_350 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_191 IVX_E ( .A(D), .Y(E) );
  NAND2_349 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_348 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_190 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_347 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_126 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_348 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_190 IVX_E ( .A(D), .Y(E) );
  NAND2_347 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_346 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_189 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_345 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_125 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_346 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_189 IVX_E ( .A(D), .Y(E) );
  NAND2_345 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_344 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_188 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_343 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_124 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_344 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_188 IVX_E ( .A(D), .Y(E) );
  NAND2_343 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_342 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_187 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_341 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_123 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_342 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_187 IVX_E ( .A(D), .Y(E) );
  NAND2_341 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_340 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_186 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_339 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_122 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_340 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_186 IVX_E ( .A(D), .Y(E) );
  NAND2_339 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_338 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_185 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_337 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_121 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_338 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_185 IVX_E ( .A(D), .Y(E) );
  NAND2_337 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_336 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_184 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_335 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_120 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_336 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_184 IVX_E ( .A(D), .Y(E) );
  NAND2_335 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_334 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_183 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_333 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_119 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_334 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_183 IVX_E ( .A(D), .Y(E) );
  NAND2_333 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_332 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_182 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_331 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_118 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_332 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_182 IVX_E ( .A(D), .Y(E) );
  NAND2_331 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_330 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_181 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_329 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_117 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_330 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_181 IVX_E ( .A(D), .Y(E) );
  NAND2_329 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_328 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_180 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_327 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_116 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_328 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_180 IVX_E ( .A(D), .Y(E) );
  NAND2_327 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_326 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_179 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_325 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_115 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_326 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_179 IVX_E ( .A(D), .Y(E) );
  NAND2_325 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_324 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_178 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_323 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_114 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_324 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_178 IVX_E ( .A(D), .Y(E) );
  NAND2_323 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_322 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_177 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_321 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_113 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_322 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_177 IVX_E ( .A(D), .Y(E) );
  NAND2_321 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_320 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_176 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_319 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_112 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_320 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_176 IVX_E ( .A(D), .Y(E) );
  NAND2_319 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_318 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_175 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_317 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_111 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_318 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_175 IVX_E ( .A(D), .Y(E) );
  NAND2_317 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_316 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_174 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_315 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_110 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_316 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_174 IVX_E ( .A(D), .Y(E) );
  NAND2_315 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_314 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_173 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_313 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_109 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_314 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_173 IVX_E ( .A(D), .Y(E) );
  NAND2_313 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_312 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_172 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_311 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_108 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_312 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_172 IVX_E ( .A(D), .Y(E) );
  NAND2_311 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_310 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_171 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_309 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_107 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_310 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_171 IVX_E ( .A(D), .Y(E) );
  NAND2_309 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_308 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_170 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_307 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_106 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_308 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_170 IVX_E ( .A(D), .Y(E) );
  NAND2_307 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_306 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_169 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_305 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_105 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_306 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_169 IVX_E ( .A(D), .Y(E) );
  NAND2_305 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_304 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_168 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_303 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_104 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_304 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_168 IVX_E ( .A(D), .Y(E) );
  NAND2_303 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_302 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_167 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_301 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_103 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_302 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_167 IVX_E ( .A(D), .Y(E) );
  NAND2_301 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_300 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_166 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_299 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_102 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_300 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_166 IVX_E ( .A(D), .Y(E) );
  NAND2_299 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_298 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_165 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_297 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_101 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_298 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_165 IVX_E ( .A(D), .Y(E) );
  NAND2_297 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_296 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_164 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_295 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_100 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_296 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_164 IVX_E ( .A(D), .Y(E) );
  NAND2_295 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_294 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_163 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_293 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_99 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_294 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_163 IVX_E ( .A(D), .Y(E) );
  NAND2_293 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_292 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_162 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_291 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_98 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_292 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_162 IVX_E ( .A(D), .Y(E) );
  NAND2_291 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_290 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_161 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_289 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_97 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_290 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_161 IVX_E ( .A(D), .Y(E) );
  NAND2_289 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_288 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_160 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_287 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_96 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_288 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_160 IVX_E ( .A(D), .Y(E) );
  NAND2_287 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_286 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_159 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_285 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_95 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_286 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_159 IVX_E ( .A(D), .Y(E) );
  NAND2_285 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_284 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_158 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_283 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_94 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_284 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_158 IVX_E ( .A(D), .Y(E) );
  NAND2_283 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_282 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_157 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_281 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_93 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_282 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_157 IVX_E ( .A(D), .Y(E) );
  NAND2_281 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_280 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_156 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_279 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_92 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_280 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_156 IVX_E ( .A(D), .Y(E) );
  NAND2_279 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_278 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_155 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_277 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_91 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_278 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_155 IVX_E ( .A(D), .Y(E) );
  NAND2_277 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_276 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_154 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_275 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_90 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_276 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_154 IVX_E ( .A(D), .Y(E) );
  NAND2_275 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_274 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_153 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_273 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_89 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_274 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_153 IVX_E ( .A(D), .Y(E) );
  NAND2_273 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_272 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_152 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_271 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_88 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_272 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_152 IVX_E ( .A(D), .Y(E) );
  NAND2_271 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_270 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_151 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_269 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_87 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_270 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_151 IVX_E ( .A(D), .Y(E) );
  NAND2_269 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_268 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_150 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_267 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_86 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_268 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_150 IVX_E ( .A(D), .Y(E) );
  NAND2_267 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_266 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_149 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_265 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_85 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_266 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_149 IVX_E ( .A(D), .Y(E) );
  NAND2_265 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_264 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_148 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_263 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_84 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_264 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_148 IVX_E ( .A(D), .Y(E) );
  NAND2_263 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_262 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_147 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_261 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_83 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_262 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_147 IVX_E ( .A(D), .Y(E) );
  NAND2_261 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_260 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_146 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_259 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_82 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_260 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_146 IVX_E ( .A(D), .Y(E) );
  NAND2_259 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_258 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_145 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_257 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_81 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_258 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_145 IVX_E ( .A(D), .Y(E) );
  NAND2_257 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_256 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_144 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_255 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_80 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_256 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_144 IVX_E ( .A(D), .Y(E) );
  NAND2_255 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_254 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_143 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_253 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_79 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_254 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_143 IVX_E ( .A(D), .Y(E) );
  NAND2_253 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_252 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_142 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_251 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_78 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_252 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_142 IVX_E ( .A(D), .Y(E) );
  NAND2_251 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_250 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_141 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_249 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_77 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_250 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_141 IVX_E ( .A(D), .Y(E) );
  NAND2_249 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_248 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_140 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_247 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_76 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_248 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_140 IVX_E ( .A(D), .Y(E) );
  NAND2_247 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_246 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_139 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_245 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_75 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_246 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_139 IVX_E ( .A(D), .Y(E) );
  NAND2_245 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_244 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_138 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_243 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_74 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_244 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_138 IVX_E ( .A(D), .Y(E) );
  NAND2_243 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_242 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_137 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_241 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_73 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_242 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_137 IVX_E ( .A(D), .Y(E) );
  NAND2_241 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_240 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_136 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_239 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_72 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_240 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_136 IVX_E ( .A(D), .Y(E) );
  NAND2_239 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_238 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_135 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_237 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_71 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_238 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_135 IVX_E ( .A(D), .Y(E) );
  NAND2_237 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_236 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_134 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_235 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_70 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_236 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_134 IVX_E ( .A(D), .Y(E) );
  NAND2_235 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_234 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_133 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_233 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_69 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_234 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_133 IVX_E ( .A(D), .Y(E) );
  NAND2_233 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_232 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_132 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_231 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_68 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_232 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_132 IVX_E ( .A(D), .Y(E) );
  NAND2_231 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_230 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_131 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_229 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_67 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_230 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_131 IVX_E ( .A(D), .Y(E) );
  NAND2_229 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_228 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_130 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_227 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_66 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_228 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_130 IVX_E ( .A(D), .Y(E) );
  NAND2_227 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_226 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_129 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_225 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_65 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_226 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_129 IVX_E ( .A(D), .Y(E) );
  NAND2_225 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_224 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_128 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_223 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_64 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_224 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_128 IVX_E ( .A(D), .Y(E) );
  NAND2_223 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_222 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_127 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_221 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_63 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_222 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_127 IVX_E ( .A(D), .Y(E) );
  NAND2_221 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_220 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_126 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_219 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_62 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_220 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_126 IVX_E ( .A(D), .Y(E) );
  NAND2_219 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_218 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_125 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_217 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_61 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_218 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_125 IVX_E ( .A(D), .Y(E) );
  NAND2_217 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_216 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_124 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_215 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_60 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_216 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_124 IVX_E ( .A(D), .Y(E) );
  NAND2_215 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_214 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_123 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_213 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_59 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_214 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_123 IVX_E ( .A(D), .Y(E) );
  NAND2_213 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_212 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_122 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_211 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_58 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_212 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_122 IVX_E ( .A(D), .Y(E) );
  NAND2_211 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_210 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_121 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_209 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_57 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_210 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_121 IVX_E ( .A(D), .Y(E) );
  NAND2_209 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_208 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_120 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_207 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_56 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_208 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_120 IVX_E ( .A(D), .Y(E) );
  NAND2_207 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_206 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_119 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_205 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_55 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_206 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_119 IVX_E ( .A(D), .Y(E) );
  NAND2_205 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_204 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_118 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_203 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_54 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_204 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_118 IVX_E ( .A(D), .Y(E) );
  NAND2_203 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_202 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_117 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_201 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_53 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_202 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_117 IVX_E ( .A(D), .Y(E) );
  NAND2_201 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_200 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_116 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_199 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_52 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_200 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_116 IVX_E ( .A(D), .Y(E) );
  NAND2_199 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_198 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_115 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_197 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_51 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_198 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_115 IVX_E ( .A(D), .Y(E) );
  NAND2_197 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_196 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_114 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_195 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_50 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_196 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_114 IVX_E ( .A(D), .Y(E) );
  NAND2_195 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_194 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_113 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_193 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_49 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_194 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_113 IVX_E ( .A(D), .Y(E) );
  NAND2_193 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_192 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_112 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_48 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_192 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_112 IVX_E ( .A(D), .Y(E) );
  NAND2_191 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_111 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_47 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_190 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_111 IVX_E ( .A(D), .Y(E) );
  NAND2_189 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_110 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_46 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_188 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_110 IVX_E ( .A(D), .Y(E) );
  NAND2_187 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_109 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_45 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_186 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_109 IVX_E ( .A(D), .Y(E) );
  NAND2_185 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_108 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_44 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_184 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_108 IVX_E ( .A(D), .Y(E) );
  NAND2_183 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_107 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_43 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_182 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_107 IVX_E ( .A(D), .Y(E) );
  NAND2_181 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_106 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_42 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_180 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_106 IVX_E ( .A(D), .Y(E) );
  NAND2_179 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_105 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_41 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_178 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_105 IVX_E ( .A(D), .Y(E) );
  NAND2_177 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_104 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_40 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_176 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_104 IVX_E ( .A(D), .Y(E) );
  NAND2_175 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_103 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_39 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_174 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_103 IVX_E ( .A(D), .Y(E) );
  NAND2_173 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_102 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_38 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_172 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_102 IVX_E ( .A(D), .Y(E) );
  NAND2_171 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_101 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_37 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_170 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_101 IVX_E ( .A(D), .Y(E) );
  NAND2_169 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_100 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_36 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_168 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_100 IVX_E ( .A(D), .Y(E) );
  NAND2_167 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_99 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_35 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_166 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_99 IVX_E ( .A(D), .Y(E) );
  NAND2_165 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_98 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_34 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_164 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_98 IVX_E ( .A(D), .Y(E) );
  NAND2_163 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_97 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_33 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_162 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_97 IVX_E ( .A(D), .Y(E) );
  NAND2_161 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_96 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_32 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_160 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_96 IVX_E ( .A(D), .Y(E) );
  NAND2_159 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_95 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_31 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_158 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_95 IVX_E ( .A(D), .Y(E) );
  NAND2_157 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_94 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_30 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_156 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_94 IVX_E ( .A(D), .Y(E) );
  NAND2_155 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_93 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_29 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_154 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_93 IVX_E ( .A(D), .Y(E) );
  NAND2_153 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_92 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_28 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_152 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_92 IVX_E ( .A(D), .Y(E) );
  NAND2_151 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_91 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_27 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_150 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_91 IVX_E ( .A(D), .Y(E) );
  NAND2_149 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_90 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_26 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_148 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_90 IVX_E ( .A(D), .Y(E) );
  NAND2_147 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_89 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_25 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_146 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_89 IVX_E ( .A(D), .Y(E) );
  NAND2_145 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_88 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_24 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_144 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_88 IVX_E ( .A(D), .Y(E) );
  NAND2_143 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_87 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_23 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_142 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_87 IVX_E ( .A(D), .Y(E) );
  NAND2_141 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_86 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_22 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_140 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_86 IVX_E ( .A(D), .Y(E) );
  NAND2_139 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_85 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_21 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_138 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_85 IVX_E ( .A(D), .Y(E) );
  NAND2_137 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_84 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_20 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_136 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_84 IVX_E ( .A(D), .Y(E) );
  NAND2_135 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_83 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_19 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_134 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_83 IVX_E ( .A(D), .Y(E) );
  NAND2_133 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_82 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_18 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_132 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_82 IVX_E ( .A(D), .Y(E) );
  NAND2_131 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_81 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_17 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_130 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_81 IVX_E ( .A(D), .Y(E) );
  NAND2_129 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_80 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_16 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_128 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_80 IVX_E ( .A(D), .Y(E) );
  NAND2_127 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_79 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_15 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_126 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_79 IVX_E ( .A(D), .Y(E) );
  NAND2_125 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_78 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_14 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_124 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_78 IVX_E ( .A(D), .Y(E) );
  NAND2_123 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_77 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_13 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_122 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_77 IVX_E ( .A(D), .Y(E) );
  NAND2_121 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_76 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_12 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_120 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_76 IVX_E ( .A(D), .Y(E) );
  NAND2_119 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_75 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_11 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_118 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_75 IVX_E ( .A(D), .Y(E) );
  NAND2_117 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_74 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_10 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_116 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_74 IVX_E ( .A(D), .Y(E) );
  NAND2_115 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_73 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_9 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_114 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_73 IVX_E ( .A(D), .Y(E) );
  NAND2_113 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_72 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_8 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_112 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_72 IVX_E ( .A(D), .Y(E) );
  NAND2_111 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_71 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_7 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_110 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_71 IVX_E ( .A(D), .Y(E) );
  NAND2_109 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_70 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_6 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_108 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_70 IVX_E ( .A(D), .Y(E) );
  NAND2_107 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_69 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_5 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_106 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_69 IVX_E ( .A(D), .Y(E) );
  NAND2_105 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_68 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_4 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_104 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_68 IVX_E ( .A(D), .Y(E) );
  NAND2_103 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_67 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_3 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_102 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_67 IVX_E ( .A(D), .Y(E) );
  NAND2_101 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_66 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_99 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_2 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_100 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_66 IVX_E ( .A(D), .Y(E) );
  NAND2_99 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_98 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_65 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_97 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND3_1 ( A, B, C, Y );
  input A, B, C;
  output Y;
  wire   D, E;

  NAND2_98 NAND_D ( .A(A), .B(B), .Y(D) );
  IVX_65 IVX_E ( .A(D), .Y(E) );
  NAND2_97 NAND_Y ( .A(E), .B(C), .Y(Y) );
endmodule


module NAND2_96 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_95 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_64 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_94 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_0 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_96 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_95 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_64 IVX_G ( .A(E), .Y(G) );
  IVX_63 IVX_H ( .A(F), .Y(H) );
  NAND2_94 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_93 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_92 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_91 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_31 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_93 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_92 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_62 IVX_G ( .A(E), .Y(G) );
  IVX_61 IVX_H ( .A(F), .Y(H) );
  NAND2_91 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_90 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_89 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_88 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_30 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_90 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_89 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_60 IVX_G ( .A(E), .Y(G) );
  IVX_59 IVX_H ( .A(F), .Y(H) );
  NAND2_88 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_87 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_86 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_85 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_29 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_87 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_86 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_58 IVX_G ( .A(E), .Y(G) );
  IVX_57 IVX_H ( .A(F), .Y(H) );
  NAND2_85 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_84 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_83 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_82 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_28 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_84 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_83 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_56 IVX_G ( .A(E), .Y(G) );
  IVX_55 IVX_H ( .A(F), .Y(H) );
  NAND2_82 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_81 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_80 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_53 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_79 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_27 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_81 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_80 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_54 IVX_G ( .A(E), .Y(G) );
  IVX_53 IVX_H ( .A(F), .Y(H) );
  NAND2_79 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_78 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_77 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_76 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_26 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_78 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_77 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_52 IVX_G ( .A(E), .Y(G) );
  IVX_51 IVX_H ( .A(F), .Y(H) );
  NAND2_76 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_75 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_74 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_73 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_25 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_75 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_74 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_50 IVX_G ( .A(E), .Y(G) );
  IVX_49 IVX_H ( .A(F), .Y(H) );
  NAND2_73 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_72 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_71 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_70 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_24 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_72 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_71 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_48 IVX_G ( .A(E), .Y(G) );
  IVX_47 IVX_H ( .A(F), .Y(H) );
  NAND2_70 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_69 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_68 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_67 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_23 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_69 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_68 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_46 IVX_G ( .A(E), .Y(G) );
  IVX_45 IVX_H ( .A(F), .Y(H) );
  NAND2_67 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_66 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_65 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_43 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_64 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_22 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_66 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_65 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_44 IVX_G ( .A(E), .Y(G) );
  IVX_43 IVX_H ( .A(F), .Y(H) );
  NAND2_64 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_63 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_62 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_61 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_21 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_63 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_62 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_42 IVX_G ( .A(E), .Y(G) );
  IVX_41 IVX_H ( .A(F), .Y(H) );
  NAND2_61 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_60 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_59 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_58 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_20 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_60 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_59 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_40 IVX_G ( .A(E), .Y(G) );
  IVX_39 IVX_H ( .A(F), .Y(H) );
  NAND2_58 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_57 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_56 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_55 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_19 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_57 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_56 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_38 IVX_G ( .A(E), .Y(G) );
  IVX_37 IVX_H ( .A(F), .Y(H) );
  NAND2_55 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_54 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_53 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_36 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_35 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_52 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_18 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_54 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_53 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_36 IVX_G ( .A(E), .Y(G) );
  IVX_35 IVX_H ( .A(F), .Y(H) );
  NAND2_52 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_51 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_50 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_49 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_17 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_51 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_50 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_34 IVX_G ( .A(E), .Y(G) );
  IVX_33 IVX_H ( .A(F), .Y(H) );
  NAND2_49 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_48 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_47 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_46 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_16 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_48 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_47 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_32 IVX_G ( .A(E), .Y(G) );
  IVX_31 IVX_H ( .A(F), .Y(H) );
  NAND2_46 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_45 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_44 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_43 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_15 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_45 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_44 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_30 IVX_G ( .A(E), .Y(G) );
  IVX_29 IVX_H ( .A(F), .Y(H) );
  NAND2_43 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_42 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_41 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_40 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_14 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_42 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_41 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_28 IVX_G ( .A(E), .Y(G) );
  IVX_27 IVX_H ( .A(F), .Y(H) );
  NAND2_40 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_39 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_38 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_26 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_37 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_13 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_39 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_38 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_26 IVX_G ( .A(E), .Y(G) );
  IVX_25 IVX_H ( .A(F), .Y(H) );
  NAND2_37 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_36 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_35 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_34 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_12 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_36 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_35 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_24 IVX_G ( .A(E), .Y(G) );
  IVX_23 IVX_H ( .A(F), .Y(H) );
  NAND2_34 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_33 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_32 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_31 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_11 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_33 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_32 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_22 IVX_G ( .A(E), .Y(G) );
  IVX_21 IVX_H ( .A(F), .Y(H) );
  NAND2_31 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_30 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_29 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_28 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_10 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_30 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_29 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_20 IVX_G ( .A(E), .Y(G) );
  IVX_19 IVX_H ( .A(F), .Y(H) );
  NAND2_28 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_27 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_26 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_25 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_9 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_27 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_26 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_18 IVX_G ( .A(E), .Y(G) );
  IVX_17 IVX_H ( .A(F), .Y(H) );
  NAND2_25 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_24 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_23 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_22 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_8 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_24 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_23 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_16 IVX_G ( .A(E), .Y(G) );
  IVX_15 IVX_H ( .A(F), .Y(H) );
  NAND2_22 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_21 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_20 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_19 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_7 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_21 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_20 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_14 IVX_G ( .A(E), .Y(G) );
  IVX_13 IVX_H ( .A(F), .Y(H) );
  NAND2_19 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_18 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_17 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_16 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_6 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_18 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_17 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_12 IVX_G ( .A(E), .Y(G) );
  IVX_11 IVX_H ( .A(F), .Y(H) );
  NAND2_16 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_15 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_14 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_10 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_13 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_5 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_15 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_14 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_10 IVX_G ( .A(E), .Y(G) );
  IVX_9 IVX_H ( .A(F), .Y(H) );
  NAND2_13 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_12 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_11 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_10 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_4 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_12 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_11 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_8 IVX_G ( .A(E), .Y(G) );
  IVX_7 IVX_H ( .A(F), .Y(H) );
  NAND2_10 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_9 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_8 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_7 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_3 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_9 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_8 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_6 IVX_G ( .A(E), .Y(G) );
  IVX_5 IVX_H ( .A(F), .Y(H) );
  NAND2_7 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_6 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_5 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_4 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_2 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_6 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_5 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_4 IVX_G ( .A(E), .Y(G) );
  IVX_3 IVX_H ( .A(F), .Y(H) );
  NAND2_4 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module NAND2_3 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND2_2 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IVX_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IVX_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module NAND2_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND4_1 ( A, B, C, D, Y );
  input A, B, C, D;
  output Y;
  wire   E, F, G, H;

  NAND2_3 NAND_E ( .A(A), .B(B), .Y(E) );
  NAND2_2 NAND_F ( .A(C), .B(D), .Y(F) );
  IVX_2 IVX_G ( .A(E), .Y(G) );
  IVX_1 IVX_H ( .A(F), .Y(H) );
  NAND2_1 NAND_Y ( .A(G), .B(H), .Y(Y) );
endmodule


module LOGIC_WIDTH32 ( R1, R2, S0, S1, S2, S3, Y );
  input [31:0] R1;
  input [31:0] R2;
  output [31:0] Y;
  input S0, S1, S2, S3;
  wire   n37, n38, n39, n40, n41, n42, n43, n44, n45;
  wire   [31:0] negR1;
  wire   [31:0] negR2;
  wire   [31:0] L0;
  wire   [31:0] L1;
  wire   [31:0] L2;
  wire   [31:0] L3;

  IVX_0 IVX_i_0 ( .A(R1[0]), .Y(negR1[0]) );
  IVX_255 IVX_i_1 ( .A(R1[1]), .Y(negR1[1]) );
  IVX_254 IVX_i_2 ( .A(R1[2]), .Y(negR1[2]) );
  IVX_253 IVX_i_3 ( .A(R1[3]), .Y(negR1[3]) );
  IVX_252 IVX_i_4 ( .A(R1[4]), .Y(negR1[4]) );
  IVX_251 IVX_i_5 ( .A(R1[5]), .Y(negR1[5]) );
  IVX_250 IVX_i_6 ( .A(R1[6]), .Y(negR1[6]) );
  IVX_249 IVX_i_7 ( .A(R1[7]), .Y(negR1[7]) );
  IVX_248 IVX_i_8 ( .A(R1[8]), .Y(negR1[8]) );
  IVX_247 IVX_i_9 ( .A(R1[9]), .Y(negR1[9]) );
  IVX_246 IVX_i_10 ( .A(R1[10]), .Y(negR1[10]) );
  IVX_245 IVX_i_11 ( .A(R1[11]), .Y(negR1[11]) );
  IVX_244 IVX_i_12 ( .A(R1[12]), .Y(negR1[12]) );
  IVX_243 IVX_i_13 ( .A(R1[13]), .Y(negR1[13]) );
  IVX_242 IVX_i_14 ( .A(R1[14]), .Y(negR1[14]) );
  IVX_241 IVX_i_15 ( .A(R1[15]), .Y(negR1[15]) );
  IVX_240 IVX_i_16 ( .A(R1[16]), .Y(negR1[16]) );
  IVX_239 IVX_i_17 ( .A(R1[17]), .Y(negR1[17]) );
  IVX_238 IVX_i_18 ( .A(R1[18]), .Y(negR1[18]) );
  IVX_237 IVX_i_19 ( .A(R1[19]), .Y(negR1[19]) );
  IVX_236 IVX_i_20 ( .A(R1[20]), .Y(negR1[20]) );
  IVX_235 IVX_i_21 ( .A(R1[21]), .Y(negR1[21]) );
  IVX_234 IVX_i_22 ( .A(R1[22]), .Y(negR1[22]) );
  IVX_233 IVX_i_23 ( .A(R1[23]), .Y(negR1[23]) );
  IVX_232 IVX_i_24 ( .A(R1[24]), .Y(negR1[24]) );
  IVX_231 IVX_i_25 ( .A(R1[25]), .Y(negR1[25]) );
  IVX_230 IVX_i_26 ( .A(R1[26]), .Y(negR1[26]) );
  IVX_229 IVX_i_27 ( .A(R1[27]), .Y(negR1[27]) );
  IVX_228 IVX_i_28 ( .A(R1[28]), .Y(negR1[28]) );
  IVX_227 IVX_i_29 ( .A(R1[29]), .Y(negR1[29]) );
  IVX_226 IVX_i_30 ( .A(R1[30]), .Y(negR1[30]) );
  IVX_225 IVX_i_31 ( .A(R1[31]), .Y(negR1[31]) );
  IVX_224 IVX_i_0_0 ( .A(R2[0]), .Y(negR2[0]) );
  IVX_223 IVX_i_1_0 ( .A(R2[1]), .Y(negR2[1]) );
  IVX_222 IVX_i_2_0 ( .A(R2[2]), .Y(negR2[2]) );
  IVX_221 IVX_i_3_0 ( .A(R2[3]), .Y(negR2[3]) );
  IVX_220 IVX_i_4_0 ( .A(R2[4]), .Y(negR2[4]) );
  IVX_219 IVX_i_5_0 ( .A(R2[5]), .Y(negR2[5]) );
  IVX_218 IVX_i_6_0 ( .A(R2[6]), .Y(negR2[6]) );
  IVX_217 IVX_i_7_0 ( .A(R2[7]), .Y(negR2[7]) );
  IVX_216 IVX_i_8_0 ( .A(R2[8]), .Y(negR2[8]) );
  IVX_215 IVX_i_9_0 ( .A(R2[9]), .Y(negR2[9]) );
  IVX_214 IVX_i_10_0 ( .A(R2[10]), .Y(negR2[10]) );
  IVX_213 IVX_i_11_0 ( .A(R2[11]), .Y(negR2[11]) );
  IVX_212 IVX_i_12_0 ( .A(R2[12]), .Y(negR2[12]) );
  IVX_211 IVX_i_13_0 ( .A(R2[13]), .Y(negR2[13]) );
  IVX_210 IVX_i_14_0 ( .A(R2[14]), .Y(negR2[14]) );
  IVX_209 IVX_i_15_0 ( .A(R2[15]), .Y(negR2[15]) );
  IVX_208 IVX_i_16_0 ( .A(R2[16]), .Y(negR2[16]) );
  IVX_207 IVX_i_17_0 ( .A(R2[17]), .Y(negR2[17]) );
  IVX_206 IVX_i_18_0 ( .A(R2[18]), .Y(negR2[18]) );
  IVX_205 IVX_i_19_0 ( .A(R2[19]), .Y(negR2[19]) );
  IVX_204 IVX_i_20_0 ( .A(R2[20]), .Y(negR2[20]) );
  IVX_203 IVX_i_21_0 ( .A(R2[21]), .Y(negR2[21]) );
  IVX_202 IVX_i_22_0 ( .A(R2[22]), .Y(negR2[22]) );
  IVX_201 IVX_i_23_0 ( .A(R2[23]), .Y(negR2[23]) );
  IVX_200 IVX_i_24_0 ( .A(R2[24]), .Y(negR2[24]) );
  IVX_199 IVX_i_25_0 ( .A(R2[25]), .Y(negR2[25]) );
  IVX_198 IVX_i_26_0 ( .A(R2[26]), .Y(negR2[26]) );
  IVX_197 IVX_i_27_0 ( .A(R2[27]), .Y(negR2[27]) );
  IVX_196 IVX_i_28_0 ( .A(R2[28]), .Y(negR2[28]) );
  IVX_195 IVX_i_29_0 ( .A(R2[29]), .Y(negR2[29]) );
  IVX_194 IVX_i_30_0 ( .A(R2[30]), .Y(negR2[30]) );
  IVX_193 IVX_i_31_0 ( .A(R2[31]), .Y(negR2[31]) );
  NAND3_0 NAND3_0i_0 ( .A(negR1[0]), .B(negR2[0]), .C(S0), .Y(L0[0]) );
  NAND3_127 NAND3_0i_1 ( .A(negR1[1]), .B(negR2[1]), .C(S0), .Y(L0[1]) );
  NAND3_126 NAND3_0i_2 ( .A(negR1[2]), .B(negR2[2]), .C(S0), .Y(L0[2]) );
  NAND3_125 NAND3_0i_3 ( .A(negR1[3]), .B(negR2[3]), .C(S0), .Y(L0[3]) );
  NAND3_124 NAND3_0i_4 ( .A(negR1[4]), .B(negR2[4]), .C(S0), .Y(L0[4]) );
  NAND3_123 NAND3_0i_5 ( .A(negR1[5]), .B(negR2[5]), .C(S0), .Y(L0[5]) );
  NAND3_122 NAND3_0i_6 ( .A(negR1[6]), .B(negR2[6]), .C(S0), .Y(L0[6]) );
  NAND3_121 NAND3_0i_7 ( .A(negR1[7]), .B(negR2[7]), .C(S0), .Y(L0[7]) );
  NAND3_120 NAND3_0i_8 ( .A(negR1[8]), .B(negR2[8]), .C(S0), .Y(L0[8]) );
  NAND3_119 NAND3_0i_9 ( .A(negR1[9]), .B(negR2[9]), .C(S0), .Y(L0[9]) );
  NAND3_118 NAND3_0i_10 ( .A(negR1[10]), .B(negR2[10]), .C(S0), .Y(L0[10]) );
  NAND3_117 NAND3_0i_11 ( .A(negR1[11]), .B(negR2[11]), .C(S0), .Y(L0[11]) );
  NAND3_116 NAND3_0i_12 ( .A(negR1[12]), .B(negR2[12]), .C(S0), .Y(L0[12]) );
  NAND3_115 NAND3_0i_13 ( .A(negR1[13]), .B(negR2[13]), .C(S0), .Y(L0[13]) );
  NAND3_114 NAND3_0i_14 ( .A(negR1[14]), .B(negR2[14]), .C(S0), .Y(L0[14]) );
  NAND3_113 NAND3_0i_15 ( .A(negR1[15]), .B(negR2[15]), .C(S0), .Y(L0[15]) );
  NAND3_112 NAND3_0i_16 ( .A(negR1[16]), .B(negR2[16]), .C(S0), .Y(L0[16]) );
  NAND3_111 NAND3_0i_17 ( .A(negR1[17]), .B(negR2[17]), .C(S0), .Y(L0[17]) );
  NAND3_110 NAND3_0i_18 ( .A(negR1[18]), .B(negR2[18]), .C(S0), .Y(L0[18]) );
  NAND3_109 NAND3_0i_19 ( .A(negR1[19]), .B(negR2[19]), .C(S0), .Y(L0[19]) );
  NAND3_108 NAND3_0i_20 ( .A(negR1[20]), .B(negR2[20]), .C(S0), .Y(L0[20]) );
  NAND3_107 NAND3_0i_21 ( .A(negR1[21]), .B(negR2[21]), .C(S0), .Y(L0[21]) );
  NAND3_106 NAND3_0i_22 ( .A(negR1[22]), .B(negR2[22]), .C(S0), .Y(L0[22]) );
  NAND3_105 NAND3_0i_23 ( .A(negR1[23]), .B(negR2[23]), .C(S0), .Y(L0[23]) );
  NAND3_104 NAND3_0i_24 ( .A(negR1[24]), .B(negR2[24]), .C(S0), .Y(L0[24]) );
  NAND3_103 NAND3_0i_25 ( .A(negR1[25]), .B(negR2[25]), .C(S0), .Y(L0[25]) );
  NAND3_102 NAND3_0i_26 ( .A(negR1[26]), .B(negR2[26]), .C(S0), .Y(L0[26]) );
  NAND3_101 NAND3_0i_27 ( .A(negR1[27]), .B(negR2[27]), .C(S0), .Y(L0[27]) );
  NAND3_100 NAND3_0i_28 ( .A(negR1[28]), .B(negR2[28]), .C(S0), .Y(L0[28]) );
  NAND3_99 NAND3_0i_29 ( .A(negR1[29]), .B(negR2[29]), .C(S0), .Y(L0[29]) );
  NAND3_98 NAND3_0i_30 ( .A(negR1[30]), .B(negR2[30]), .C(S0), .Y(L0[30]) );
  NAND3_97 NAND3_0i_31 ( .A(negR1[31]), .B(negR2[31]), .C(S0), .Y(L0[31]) );
  NAND3_96 NAND3_1i_0 ( .A(negR1[0]), .B(R2[0]), .C(n37), .Y(L1[0]) );
  NAND3_95 NAND3_1i_1 ( .A(negR1[1]), .B(R2[1]), .C(n37), .Y(L1[1]) );
  NAND3_94 NAND3_1i_2 ( .A(negR1[2]), .B(R2[2]), .C(n37), .Y(L1[2]) );
  NAND3_93 NAND3_1i_3 ( .A(negR1[3]), .B(R2[3]), .C(n37), .Y(L1[3]) );
  NAND3_92 NAND3_1i_4 ( .A(negR1[4]), .B(R2[4]), .C(n37), .Y(L1[4]) );
  NAND3_91 NAND3_1i_5 ( .A(negR1[5]), .B(R2[5]), .C(n37), .Y(L1[5]) );
  NAND3_90 NAND3_1i_6 ( .A(negR1[6]), .B(R2[6]), .C(n37), .Y(L1[6]) );
  NAND3_89 NAND3_1i_7 ( .A(negR1[7]), .B(R2[7]), .C(n37), .Y(L1[7]) );
  NAND3_88 NAND3_1i_8 ( .A(negR1[8]), .B(R2[8]), .C(n37), .Y(L1[8]) );
  NAND3_87 NAND3_1i_9 ( .A(negR1[9]), .B(R2[9]), .C(n37), .Y(L1[9]) );
  NAND3_86 NAND3_1i_10 ( .A(negR1[10]), .B(R2[10]), .C(n37), .Y(L1[10]) );
  NAND3_85 NAND3_1i_11 ( .A(negR1[11]), .B(R2[11]), .C(n37), .Y(L1[11]) );
  NAND3_84 NAND3_1i_12 ( .A(negR1[12]), .B(R2[12]), .C(n38), .Y(L1[12]) );
  NAND3_83 NAND3_1i_13 ( .A(negR1[13]), .B(R2[13]), .C(n38), .Y(L1[13]) );
  NAND3_82 NAND3_1i_14 ( .A(negR1[14]), .B(R2[14]), .C(n38), .Y(L1[14]) );
  NAND3_81 NAND3_1i_15 ( .A(negR1[15]), .B(R2[15]), .C(n38), .Y(L1[15]) );
  NAND3_80 NAND3_1i_16 ( .A(negR1[16]), .B(R2[16]), .C(n38), .Y(L1[16]) );
  NAND3_79 NAND3_1i_17 ( .A(negR1[17]), .B(R2[17]), .C(n38), .Y(L1[17]) );
  NAND3_78 NAND3_1i_18 ( .A(negR1[18]), .B(R2[18]), .C(n38), .Y(L1[18]) );
  NAND3_77 NAND3_1i_19 ( .A(negR1[19]), .B(R2[19]), .C(n38), .Y(L1[19]) );
  NAND3_76 NAND3_1i_20 ( .A(negR1[20]), .B(R2[20]), .C(n38), .Y(L1[20]) );
  NAND3_75 NAND3_1i_21 ( .A(negR1[21]), .B(R2[21]), .C(n38), .Y(L1[21]) );
  NAND3_74 NAND3_1i_22 ( .A(negR1[22]), .B(R2[22]), .C(n38), .Y(L1[22]) );
  NAND3_73 NAND3_1i_23 ( .A(negR1[23]), .B(R2[23]), .C(n38), .Y(L1[23]) );
  NAND3_72 NAND3_1i_24 ( .A(negR1[24]), .B(R2[24]), .C(n39), .Y(L1[24]) );
  NAND3_71 NAND3_1i_25 ( .A(negR1[25]), .B(R2[25]), .C(n39), .Y(L1[25]) );
  NAND3_70 NAND3_1i_26 ( .A(negR1[26]), .B(R2[26]), .C(n39), .Y(L1[26]) );
  NAND3_69 NAND3_1i_27 ( .A(negR1[27]), .B(R2[27]), .C(n39), .Y(L1[27]) );
  NAND3_68 NAND3_1i_28 ( .A(negR1[28]), .B(R2[28]), .C(n39), .Y(L1[28]) );
  NAND3_67 NAND3_1i_29 ( .A(negR1[29]), .B(R2[29]), .C(n39), .Y(L1[29]) );
  NAND3_66 NAND3_1i_30 ( .A(negR1[30]), .B(R2[30]), .C(n39), .Y(L1[30]) );
  NAND3_65 NAND3_1i_31 ( .A(negR1[31]), .B(R2[31]), .C(n39), .Y(L1[31]) );
  NAND3_64 NAND3_2i_0 ( .A(R1[0]), .B(negR2[0]), .C(n40), .Y(L2[0]) );
  NAND3_63 NAND3_2i_1 ( .A(R1[1]), .B(negR2[1]), .C(n40), .Y(L2[1]) );
  NAND3_62 NAND3_2i_2 ( .A(R1[2]), .B(negR2[2]), .C(n40), .Y(L2[2]) );
  NAND3_61 NAND3_2i_3 ( .A(R1[3]), .B(negR2[3]), .C(n40), .Y(L2[3]) );
  NAND3_60 NAND3_2i_4 ( .A(R1[4]), .B(negR2[4]), .C(n40), .Y(L2[4]) );
  NAND3_59 NAND3_2i_5 ( .A(R1[5]), .B(negR2[5]), .C(n40), .Y(L2[5]) );
  NAND3_58 NAND3_2i_6 ( .A(R1[6]), .B(negR2[6]), .C(n40), .Y(L2[6]) );
  NAND3_57 NAND3_2i_7 ( .A(R1[7]), .B(negR2[7]), .C(n40), .Y(L2[7]) );
  NAND3_56 NAND3_2i_8 ( .A(R1[8]), .B(negR2[8]), .C(n40), .Y(L2[8]) );
  NAND3_55 NAND3_2i_9 ( .A(R1[9]), .B(negR2[9]), .C(n40), .Y(L2[9]) );
  NAND3_54 NAND3_2i_10 ( .A(R1[10]), .B(negR2[10]), .C(n40), .Y(L2[10]) );
  NAND3_53 NAND3_2i_11 ( .A(R1[11]), .B(negR2[11]), .C(n40), .Y(L2[11]) );
  NAND3_52 NAND3_2i_12 ( .A(R1[12]), .B(negR2[12]), .C(n41), .Y(L2[12]) );
  NAND3_51 NAND3_2i_13 ( .A(R1[13]), .B(negR2[13]), .C(n41), .Y(L2[13]) );
  NAND3_50 NAND3_2i_14 ( .A(R1[14]), .B(negR2[14]), .C(n41), .Y(L2[14]) );
  NAND3_49 NAND3_2i_15 ( .A(R1[15]), .B(negR2[15]), .C(n41), .Y(L2[15]) );
  NAND3_48 NAND3_2i_16 ( .A(R1[16]), .B(negR2[16]), .C(n41), .Y(L2[16]) );
  NAND3_47 NAND3_2i_17 ( .A(R1[17]), .B(negR2[17]), .C(n41), .Y(L2[17]) );
  NAND3_46 NAND3_2i_18 ( .A(R1[18]), .B(negR2[18]), .C(n41), .Y(L2[18]) );
  NAND3_45 NAND3_2i_19 ( .A(R1[19]), .B(negR2[19]), .C(n41), .Y(L2[19]) );
  NAND3_44 NAND3_2i_20 ( .A(R1[20]), .B(negR2[20]), .C(n41), .Y(L2[20]) );
  NAND3_43 NAND3_2i_21 ( .A(R1[21]), .B(negR2[21]), .C(n41), .Y(L2[21]) );
  NAND3_42 NAND3_2i_22 ( .A(R1[22]), .B(negR2[22]), .C(n41), .Y(L2[22]) );
  NAND3_41 NAND3_2i_23 ( .A(R1[23]), .B(negR2[23]), .C(n41), .Y(L2[23]) );
  NAND3_40 NAND3_2i_24 ( .A(R1[24]), .B(negR2[24]), .C(n42), .Y(L2[24]) );
  NAND3_39 NAND3_2i_25 ( .A(R1[25]), .B(negR2[25]), .C(n42), .Y(L2[25]) );
  NAND3_38 NAND3_2i_26 ( .A(R1[26]), .B(negR2[26]), .C(n42), .Y(L2[26]) );
  NAND3_37 NAND3_2i_27 ( .A(R1[27]), .B(negR2[27]), .C(n42), .Y(L2[27]) );
  NAND3_36 NAND3_2i_28 ( .A(R1[28]), .B(negR2[28]), .C(n42), .Y(L2[28]) );
  NAND3_35 NAND3_2i_29 ( .A(R1[29]), .B(negR2[29]), .C(n42), .Y(L2[29]) );
  NAND3_34 NAND3_2i_30 ( .A(R1[30]), .B(negR2[30]), .C(n42), .Y(L2[30]) );
  NAND3_33 NAND3_2i_31 ( .A(R1[31]), .B(negR2[31]), .C(n42), .Y(L2[31]) );
  NAND3_32 NAND3_3i_0 ( .A(R1[0]), .B(R2[0]), .C(n43), .Y(L3[0]) );
  NAND3_31 NAND3_3i_1 ( .A(R1[1]), .B(R2[1]), .C(n43), .Y(L3[1]) );
  NAND3_30 NAND3_3i_2 ( .A(R1[2]), .B(R2[2]), .C(n43), .Y(L3[2]) );
  NAND3_29 NAND3_3i_3 ( .A(R1[3]), .B(R2[3]), .C(n43), .Y(L3[3]) );
  NAND3_28 NAND3_3i_4 ( .A(R1[4]), .B(R2[4]), .C(n43), .Y(L3[4]) );
  NAND3_27 NAND3_3i_5 ( .A(R1[5]), .B(R2[5]), .C(n43), .Y(L3[5]) );
  NAND3_26 NAND3_3i_6 ( .A(R1[6]), .B(R2[6]), .C(n43), .Y(L3[6]) );
  NAND3_25 NAND3_3i_7 ( .A(R1[7]), .B(R2[7]), .C(n43), .Y(L3[7]) );
  NAND3_24 NAND3_3i_8 ( .A(R1[8]), .B(R2[8]), .C(n43), .Y(L3[8]) );
  NAND3_23 NAND3_3i_9 ( .A(R1[9]), .B(R2[9]), .C(n43), .Y(L3[9]) );
  NAND3_22 NAND3_3i_10 ( .A(R1[10]), .B(R2[10]), .C(n43), .Y(L3[10]) );
  NAND3_21 NAND3_3i_11 ( .A(R1[11]), .B(R2[11]), .C(n43), .Y(L3[11]) );
  NAND3_20 NAND3_3i_12 ( .A(R1[12]), .B(R2[12]), .C(n44), .Y(L3[12]) );
  NAND3_19 NAND3_3i_13 ( .A(R1[13]), .B(R2[13]), .C(n44), .Y(L3[13]) );
  NAND3_18 NAND3_3i_14 ( .A(R1[14]), .B(R2[14]), .C(n44), .Y(L3[14]) );
  NAND3_17 NAND3_3i_15 ( .A(R1[15]), .B(R2[15]), .C(n44), .Y(L3[15]) );
  NAND3_16 NAND3_3i_16 ( .A(R1[16]), .B(R2[16]), .C(n44), .Y(L3[16]) );
  NAND3_15 NAND3_3i_17 ( .A(R1[17]), .B(R2[17]), .C(n44), .Y(L3[17]) );
  NAND3_14 NAND3_3i_18 ( .A(R1[18]), .B(R2[18]), .C(n44), .Y(L3[18]) );
  NAND3_13 NAND3_3i_19 ( .A(R1[19]), .B(R2[19]), .C(n44), .Y(L3[19]) );
  NAND3_12 NAND3_3i_20 ( .A(R1[20]), .B(R2[20]), .C(n44), .Y(L3[20]) );
  NAND3_11 NAND3_3i_21 ( .A(R1[21]), .B(R2[21]), .C(n44), .Y(L3[21]) );
  NAND3_10 NAND3_3i_22 ( .A(R1[22]), .B(R2[22]), .C(n44), .Y(L3[22]) );
  NAND3_9 NAND3_3i_23 ( .A(R1[23]), .B(R2[23]), .C(n44), .Y(L3[23]) );
  NAND3_8 NAND3_3i_24 ( .A(R1[24]), .B(R2[24]), .C(n45), .Y(L3[24]) );
  NAND3_7 NAND3_3i_25 ( .A(R1[25]), .B(R2[25]), .C(n45), .Y(L3[25]) );
  NAND3_6 NAND3_3i_26 ( .A(R1[26]), .B(R2[26]), .C(n45), .Y(L3[26]) );
  NAND3_5 NAND3_3i_27 ( .A(R1[27]), .B(R2[27]), .C(n45), .Y(L3[27]) );
  NAND3_4 NAND3_3i_28 ( .A(R1[28]), .B(R2[28]), .C(n45), .Y(L3[28]) );
  NAND3_3 NAND3_3i_29 ( .A(R1[29]), .B(R2[29]), .C(n45), .Y(L3[29]) );
  NAND3_2 NAND3_3i_30 ( .A(R1[30]), .B(R2[30]), .C(n45), .Y(L3[30]) );
  NAND3_1 NAND3_3i_31 ( .A(R1[31]), .B(R2[31]), .C(n45), .Y(L3[31]) );
  NAND4_0 NAND4_i_0 ( .A(L0[0]), .B(L1[0]), .C(L2[0]), .D(L3[0]), .Y(Y[0]) );
  NAND4_31 NAND4_i_1 ( .A(L0[1]), .B(L1[1]), .C(L2[1]), .D(L3[1]), .Y(Y[1]) );
  NAND4_30 NAND4_i_2 ( .A(L0[2]), .B(L1[2]), .C(L2[2]), .D(L3[2]), .Y(Y[2]) );
  NAND4_29 NAND4_i_3 ( .A(L0[3]), .B(L1[3]), .C(L2[3]), .D(L3[3]), .Y(Y[3]) );
  NAND4_28 NAND4_i_4 ( .A(L0[4]), .B(L1[4]), .C(L2[4]), .D(L3[4]), .Y(Y[4]) );
  NAND4_27 NAND4_i_5 ( .A(L0[5]), .B(L1[5]), .C(L2[5]), .D(L3[5]), .Y(Y[5]) );
  NAND4_26 NAND4_i_6 ( .A(L0[6]), .B(L1[6]), .C(L2[6]), .D(L3[6]), .Y(Y[6]) );
  NAND4_25 NAND4_i_7 ( .A(L0[7]), .B(L1[7]), .C(L2[7]), .D(L3[7]), .Y(Y[7]) );
  NAND4_24 NAND4_i_8 ( .A(L0[8]), .B(L1[8]), .C(L2[8]), .D(L3[8]), .Y(Y[8]) );
  NAND4_23 NAND4_i_9 ( .A(L0[9]), .B(L1[9]), .C(L2[9]), .D(L3[9]), .Y(Y[9]) );
  NAND4_22 NAND4_i_10 ( .A(L0[10]), .B(L1[10]), .C(L2[10]), .D(L3[10]), .Y(
        Y[10]) );
  NAND4_21 NAND4_i_11 ( .A(L0[11]), .B(L1[11]), .C(L2[11]), .D(L3[11]), .Y(
        Y[11]) );
  NAND4_20 NAND4_i_12 ( .A(L0[12]), .B(L1[12]), .C(L2[12]), .D(L3[12]), .Y(
        Y[12]) );
  NAND4_19 NAND4_i_13 ( .A(L0[13]), .B(L1[13]), .C(L2[13]), .D(L3[13]), .Y(
        Y[13]) );
  NAND4_18 NAND4_i_14 ( .A(L0[14]), .B(L1[14]), .C(L2[14]), .D(L3[14]), .Y(
        Y[14]) );
  NAND4_17 NAND4_i_15 ( .A(L0[15]), .B(L1[15]), .C(L2[15]), .D(L3[15]), .Y(
        Y[15]) );
  NAND4_16 NAND4_i_16 ( .A(L0[16]), .B(L1[16]), .C(L2[16]), .D(L3[16]), .Y(
        Y[16]) );
  NAND4_15 NAND4_i_17 ( .A(L0[17]), .B(L1[17]), .C(L2[17]), .D(L3[17]), .Y(
        Y[17]) );
  NAND4_14 NAND4_i_18 ( .A(L0[18]), .B(L1[18]), .C(L2[18]), .D(L3[18]), .Y(
        Y[18]) );
  NAND4_13 NAND4_i_19 ( .A(L0[19]), .B(L1[19]), .C(L2[19]), .D(L3[19]), .Y(
        Y[19]) );
  NAND4_12 NAND4_i_20 ( .A(L0[20]), .B(L1[20]), .C(L2[20]), .D(L3[20]), .Y(
        Y[20]) );
  NAND4_11 NAND4_i_21 ( .A(L0[21]), .B(L1[21]), .C(L2[21]), .D(L3[21]), .Y(
        Y[21]) );
  NAND4_10 NAND4_i_22 ( .A(L0[22]), .B(L1[22]), .C(L2[22]), .D(L3[22]), .Y(
        Y[22]) );
  NAND4_9 NAND4_i_23 ( .A(L0[23]), .B(L1[23]), .C(L2[23]), .D(L3[23]), .Y(
        Y[23]) );
  NAND4_8 NAND4_i_24 ( .A(L0[24]), .B(L1[24]), .C(L2[24]), .D(L3[24]), .Y(
        Y[24]) );
  NAND4_7 NAND4_i_25 ( .A(L0[25]), .B(L1[25]), .C(L2[25]), .D(L3[25]), .Y(
        Y[25]) );
  NAND4_6 NAND4_i_26 ( .A(L0[26]), .B(L1[26]), .C(L2[26]), .D(L3[26]), .Y(
        Y[26]) );
  NAND4_5 NAND4_i_27 ( .A(L0[27]), .B(L1[27]), .C(L2[27]), .D(L3[27]), .Y(
        Y[27]) );
  NAND4_4 NAND4_i_28 ( .A(L0[28]), .B(L1[28]), .C(L2[28]), .D(L3[28]), .Y(
        Y[28]) );
  NAND4_3 NAND4_i_29 ( .A(L0[29]), .B(L1[29]), .C(L2[29]), .D(L3[29]), .Y(
        Y[29]) );
  NAND4_2 NAND4_i_30 ( .A(L0[30]), .B(L1[30]), .C(L2[30]), .D(L3[30]), .Y(
        Y[30]) );
  NAND4_1 NAND4_i_31 ( .A(L0[31]), .B(L1[31]), .C(L2[31]), .D(L3[31]), .Y(
        Y[31]) );
  BUF_X1 U1 ( .A(S1), .Z(n37) );
  BUF_X1 U2 ( .A(S2), .Z(n40) );
  BUF_X1 U3 ( .A(S3), .Z(n43) );
  BUF_X1 U4 ( .A(S1), .Z(n38) );
  BUF_X1 U5 ( .A(S2), .Z(n41) );
  BUF_X1 U6 ( .A(S3), .Z(n44) );
  BUF_X1 U7 ( .A(S1), .Z(n39) );
  BUF_X1 U8 ( .A(S2), .Z(n42) );
  BUF_X1 U9 ( .A(S3), .Z(n45) );
endmodule


module COMPARATOR ( Z, C, LE, LT, GE, GT, EQ, NE );
  input Z, C;
  output LE, LT, GE, GT, EQ, NE;
  wire   C, Z;
  assign GE = C;
  assign EQ = Z;

  INV_X1 U1 ( .A(Z), .ZN(NE) );
  INV_X1 U2 ( .A(LE), .ZN(GT) );
  INV_X1 U3 ( .A(C), .ZN(LT) );
  NAND2_X1 U4 ( .A1(C), .A2(NE), .ZN(LE) );
endmodule


module MASK_GENERATOR ( op, sel, mask00, mask08, mask16 );
  input [31:0] op;
  input [1:0] sel;
  output [38:0] mask00;
  output [38:0] mask08;
  output [38:0] mask16;
  wire   \mask08[30] , \mask08[29] , \mask08[28] , \mask08[27] , \mask08[26] ,
         \mask08[25] , \mask08[24] , \mask08[14] , \mask08[13] , \mask08[12] ,
         \mask08[11] , \mask08[10] , \mask08[9] , \mask08[8] , n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, \mask16[16] , n332, n334,
         n336, n338, n340, n342, n344, n346, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n366, n368, n370, n372, n374, n376, n379, n380, n381;
  assign mask16[38] = \mask08[30] ;
  assign mask08[30] = \mask08[30] ;
  assign mask16[37] = \mask08[29] ;
  assign mask08[29] = \mask08[29] ;
  assign mask16[36] = \mask08[28] ;
  assign mask08[28] = \mask08[28] ;
  assign mask16[35] = \mask08[27] ;
  assign mask08[27] = \mask08[27] ;
  assign mask16[34] = \mask08[26] ;
  assign mask08[26] = \mask08[26] ;
  assign mask16[33] = \mask08[25] ;
  assign mask08[25] = \mask08[25] ;
  assign mask16[32] = \mask08[24] ;
  assign mask08[24] = \mask08[24] ;
  assign mask16[6] = \mask08[14] ;
  assign mask08[14] = \mask08[14] ;
  assign mask16[5] = \mask08[13] ;
  assign mask08[13] = \mask08[13] ;
  assign mask16[4] = \mask08[12] ;
  assign mask08[12] = \mask08[12] ;
  assign mask16[3] = \mask08[11] ;
  assign mask08[11] = \mask08[11] ;
  assign mask16[2] = \mask08[10] ;
  assign mask08[10] = \mask08[10] ;
  assign mask16[1] = \mask08[9] ;
  assign mask08[9] = \mask08[9] ;
  assign mask16[0] = \mask08[8] ;
  assign mask08[8] = \mask08[8] ;
  assign mask16[17] = \mask16[16] ;
  assign mask16[18] = \mask16[16] ;
  assign mask16[20] = \mask16[16] ;
  assign mask16[21] = \mask16[16] ;
  assign mask16[22] = \mask16[16] ;
  assign mask16[19] = \mask16[16] ;
  assign mask16[16] = \mask16[16] ;

  NAND3_X1 U161 ( .A1(sel[1]), .A2(n381), .A3(op[31]), .ZN(n54) );
  NOR2_X1 U2 ( .A1(sel[0]), .A2(sel[1]), .ZN(n79) );
  BUF_X1 U3 ( .A(n322), .Z(n324) );
  BUF_X1 U4 ( .A(n322), .Z(n325) );
  BUF_X1 U5 ( .A(n323), .Z(n326) );
  BUF_X1 U6 ( .A(n323), .Z(n327) );
  INV_X1 U7 ( .A(n329), .ZN(n328) );
  INV_X1 U8 ( .A(\mask16[16] ), .ZN(n330) );
  BUF_X1 U9 ( .A(n380), .Z(n322) );
  INV_X1 U10 ( .A(mask16[7]), .ZN(n348) );
  BUF_X1 U11 ( .A(n380), .Z(n323) );
  INV_X1 U12 ( .A(\mask08[8] ), .ZN(n362) );
  INV_X1 U13 ( .A(\mask08[9] ), .ZN(n360) );
  INV_X1 U14 ( .A(\mask08[10] ), .ZN(n358) );
  INV_X1 U15 ( .A(\mask08[11] ), .ZN(n356) );
  INV_X1 U16 ( .A(\mask08[12] ), .ZN(n354) );
  INV_X1 U17 ( .A(\mask08[13] ), .ZN(n352) );
  INV_X1 U18 ( .A(\mask08[14] ), .ZN(n350) );
  NOR2_X1 U19 ( .A1(n361), .A2(n329), .ZN(\mask08[9] ) );
  NOR2_X1 U20 ( .A1(n355), .A2(n329), .ZN(\mask08[12] ) );
  NOR2_X1 U21 ( .A1(n353), .A2(n329), .ZN(\mask08[13] ) );
  NOR2_X1 U22 ( .A1(n351), .A2(n329), .ZN(\mask08[14] ) );
  NOR2_X1 U23 ( .A1(n363), .A2(n329), .ZN(\mask08[8] ) );
  NOR2_X1 U24 ( .A1(n359), .A2(n329), .ZN(\mask08[10] ) );
  NOR2_X1 U25 ( .A1(n357), .A2(n329), .ZN(\mask08[11] ) );
  OAI21_X1 U26 ( .B1(n370), .B2(n324), .A(n54), .ZN(\mask08[27] ) );
  OAI21_X1 U27 ( .B1(n368), .B2(n324), .A(n330), .ZN(\mask08[28] ) );
  OAI21_X1 U28 ( .B1(n374), .B2(n324), .A(n54), .ZN(\mask08[25] ) );
  OAI21_X1 U29 ( .B1(n376), .B2(n324), .A(n330), .ZN(\mask08[24] ) );
  OAI21_X1 U30 ( .B1(n372), .B2(n324), .A(n54), .ZN(\mask08[26] ) );
  OAI21_X1 U31 ( .B1(n366), .B2(n324), .A(n330), .ZN(\mask08[29] ) );
  OAI21_X1 U32 ( .B1(n364), .B2(n324), .A(n330), .ZN(\mask08[30] ) );
  NOR2_X1 U33 ( .A1(n349), .A2(n329), .ZN(mask16[7]) );
  INV_X1 U34 ( .A(n54), .ZN(\mask16[16] ) );
  INV_X1 U35 ( .A(n61), .ZN(mask16[8]) );
  NAND2_X1 U36 ( .A1(n69), .A2(n77), .ZN(mask00[8]) );
  INV_X1 U37 ( .A(n60), .ZN(mask16[9]) );
  NAND2_X1 U38 ( .A1(n68), .A2(n76), .ZN(mask00[9]) );
  INV_X1 U39 ( .A(n59), .ZN(mask16[10]) );
  NAND2_X1 U40 ( .A1(n67), .A2(n75), .ZN(mask00[10]) );
  INV_X1 U41 ( .A(n58), .ZN(mask16[11]) );
  NAND2_X1 U42 ( .A1(n66), .A2(n74), .ZN(mask00[11]) );
  INV_X1 U43 ( .A(n62), .ZN(mask08[7]) );
  OAI21_X1 U44 ( .B1(n329), .B2(n379), .A(n78), .ZN(mask00[7]) );
  OAI21_X1 U45 ( .B1(n326), .B2(n363), .A(n348), .ZN(mask00[23]) );
  OAI21_X1 U46 ( .B1(n349), .B2(n325), .A(n330), .ZN(mask08[38]) );
  OAI21_X1 U47 ( .B1(n327), .B2(n351), .A(n330), .ZN(mask08[37]) );
  INV_X1 U48 ( .A(n57), .ZN(mask16[12]) );
  NAND2_X1 U49 ( .A1(n65), .A2(n73), .ZN(mask00[12]) );
  INV_X1 U50 ( .A(n56), .ZN(mask16[13]) );
  NAND2_X1 U51 ( .A1(n64), .A2(n72), .ZN(mask00[13]) );
  INV_X1 U52 ( .A(n55), .ZN(mask16[14]) );
  NAND2_X1 U53 ( .A1(n63), .A2(n71), .ZN(mask00[14]) );
  NAND2_X1 U54 ( .A1(n54), .A2(n77), .ZN(mask16[24]) );
  OAI21_X1 U55 ( .B1(n326), .B2(n361), .A(n61), .ZN(mask00[24]) );
  NAND2_X1 U56 ( .A1(n54), .A2(n76), .ZN(mask16[25]) );
  OAI21_X1 U57 ( .B1(n326), .B2(n359), .A(n60), .ZN(mask00[25]) );
  NAND2_X1 U58 ( .A1(n54), .A2(n75), .ZN(mask16[26]) );
  OAI21_X1 U59 ( .B1(n326), .B2(n357), .A(n59), .ZN(mask00[26]) );
  NAND2_X1 U60 ( .A1(n54), .A2(n74), .ZN(mask16[27]) );
  OAI21_X1 U61 ( .B1(n326), .B2(n355), .A(n58), .ZN(mask00[27]) );
  NAND2_X1 U62 ( .A1(n54), .A2(n73), .ZN(mask16[28]) );
  OAI21_X1 U63 ( .B1(n326), .B2(n353), .A(n57), .ZN(mask00[28]) );
  NAND2_X1 U64 ( .A1(n54), .A2(n72), .ZN(mask16[29]) );
  OAI21_X1 U65 ( .B1(n326), .B2(n351), .A(n56), .ZN(mask00[29]) );
  NAND2_X1 U66 ( .A1(n54), .A2(n71), .ZN(mask16[30]) );
  OAI21_X1 U67 ( .B1(n349), .B2(n325), .A(n55), .ZN(mask00[30]) );
  INV_X1 U68 ( .A(n53), .ZN(mask16[15]) );
  NAND2_X1 U69 ( .A1(n348), .A2(n78), .ZN(mask08[15]) );
  NAND2_X1 U70 ( .A1(n59), .A2(n75), .ZN(mask08[18]) );
  OAI21_X1 U71 ( .B1(n372), .B2(n325), .A(n358), .ZN(mask00[18]) );
  NAND2_X1 U72 ( .A1(n58), .A2(n74), .ZN(mask08[19]) );
  OAI21_X1 U73 ( .B1(n370), .B2(n325), .A(n356), .ZN(mask00[19]) );
  NAND2_X1 U74 ( .A1(n57), .A2(n73), .ZN(mask08[20]) );
  OAI21_X1 U75 ( .B1(n368), .B2(n325), .A(n354), .ZN(mask00[20]) );
  NAND2_X1 U76 ( .A1(n56), .A2(n72), .ZN(mask08[21]) );
  OAI21_X1 U77 ( .B1(n366), .B2(n325), .A(n352), .ZN(mask00[21]) );
  NAND2_X1 U78 ( .A1(n55), .A2(n71), .ZN(mask08[22]) );
  OAI21_X1 U79 ( .B1(n364), .B2(n325), .A(n350), .ZN(mask00[22]) );
  NAND2_X1 U80 ( .A1(n53), .A2(n70), .ZN(mask08[23]) );
  NAND2_X1 U81 ( .A1(n54), .A2(n78), .ZN(mask16[23]) );
  OAI21_X1 U82 ( .B1(n326), .B2(n359), .A(n330), .ZN(mask08[33]) );
  NAND2_X1 U83 ( .A1(n61), .A2(n77), .ZN(mask08[16]) );
  OAI21_X1 U84 ( .B1(n376), .B2(n324), .A(n362), .ZN(mask00[16]) );
  NAND2_X1 U85 ( .A1(n60), .A2(n76), .ZN(mask08[17]) );
  OAI21_X1 U86 ( .B1(n374), .B2(n325), .A(n360), .ZN(mask00[17]) );
  OAI21_X1 U87 ( .B1(n327), .B2(n357), .A(n330), .ZN(mask08[34]) );
  NAND2_X1 U88 ( .A1(n54), .A2(n70), .ZN(mask16[31]) );
  OAI21_X1 U89 ( .B1(n326), .B2(n363), .A(n330), .ZN(mask08[31]) );
  OAI21_X1 U90 ( .B1(n326), .B2(n361), .A(n330), .ZN(mask08[32]) );
  OAI21_X1 U91 ( .B1(n344), .B2(n325), .A(n330), .ZN(mask00[32]) );
  OAI21_X1 U92 ( .B1(n326), .B2(n353), .A(n330), .ZN(mask08[36]) );
  OAI21_X1 U93 ( .B1(n336), .B2(n324), .A(n54), .ZN(mask00[36]) );
  OAI21_X1 U94 ( .B1(n326), .B2(n355), .A(n330), .ZN(mask08[35]) );
  OAI21_X1 U95 ( .B1(n338), .B2(n324), .A(n330), .ZN(mask00[35]) );
  INV_X1 U96 ( .A(n79), .ZN(n380) );
  NAND2_X1 U97 ( .A1(n62), .A2(n70), .ZN(mask00[15]) );
  INV_X1 U98 ( .A(n68), .ZN(mask08[1]) );
  AND2_X1 U99 ( .A1(n80), .A2(op[1]), .ZN(mask00[1]) );
  AOI21_X1 U100 ( .B1(sel[0]), .B2(sel[1]), .A(n79), .ZN(n80) );
  INV_X1 U101 ( .A(sel[0]), .ZN(n381) );
  NAND2_X1 U102 ( .A1(n79), .A2(op[8]), .ZN(n70) );
  INV_X1 U103 ( .A(n63), .ZN(mask08[6]) );
  AND2_X1 U104 ( .A1(n80), .A2(op[6]), .ZN(mask00[6]) );
  NAND2_X1 U105 ( .A1(op[24]), .A2(n328), .ZN(n61) );
  NAND2_X1 U106 ( .A1(op[25]), .A2(n328), .ZN(n60) );
  NAND2_X1 U107 ( .A1(op[26]), .A2(n328), .ZN(n59) );
  NAND2_X1 U108 ( .A1(op[27]), .A2(n328), .ZN(n58) );
  NAND2_X1 U109 ( .A1(op[28]), .A2(n328), .ZN(n57) );
  NAND2_X1 U110 ( .A1(op[29]), .A2(n328), .ZN(n56) );
  NAND2_X1 U111 ( .A1(op[30]), .A2(n328), .ZN(n55) );
  NAND2_X1 U112 ( .A1(op[31]), .A2(n328), .ZN(n53) );
  NAND2_X1 U113 ( .A1(op[1]), .A2(n79), .ZN(n77) );
  NAND2_X1 U114 ( .A1(op[2]), .A2(n79), .ZN(n76) );
  NAND2_X1 U115 ( .A1(op[3]), .A2(n79), .ZN(n75) );
  NAND2_X1 U116 ( .A1(op[4]), .A2(n79), .ZN(n74) );
  NAND2_X1 U117 ( .A1(op[5]), .A2(n79), .ZN(n73) );
  NAND2_X1 U118 ( .A1(op[6]), .A2(n79), .ZN(n72) );
  NAND2_X1 U119 ( .A1(op[7]), .A2(n79), .ZN(n71) );
  NAND2_X1 U120 ( .A1(op[0]), .A2(n79), .ZN(n78) );
  OAI21_X1 U121 ( .B1(n346), .B2(n325), .A(n53), .ZN(mask00[31]) );
  INV_X1 U122 ( .A(op[24]), .ZN(n346) );
  OAI21_X1 U123 ( .B1(n342), .B2(n325), .A(n54), .ZN(mask00[33]) );
  INV_X1 U124 ( .A(op[26]), .ZN(n342) );
  OAI21_X1 U125 ( .B1(n340), .B2(n325), .A(n330), .ZN(mask00[34]) );
  INV_X1 U126 ( .A(op[27]), .ZN(n340) );
  OAI21_X1 U127 ( .B1(n334), .B2(n324), .A(n54), .ZN(mask00[37]) );
  INV_X1 U128 ( .A(op[30]), .ZN(n334) );
  OAI21_X1 U129 ( .B1(n332), .B2(n324), .A(n330), .ZN(mask00[38]) );
  INV_X1 U130 ( .A(op[31]), .ZN(n332) );
  NAND2_X1 U131 ( .A1(op[13]), .A2(n328), .ZN(n64) );
  NAND2_X1 U132 ( .A1(op[15]), .A2(n328), .ZN(n62) );
  NAND2_X1 U133 ( .A1(op[8]), .A2(n328), .ZN(n69) );
  NAND2_X1 U134 ( .A1(op[11]), .A2(n328), .ZN(n66) );
  INV_X1 U135 ( .A(n65), .ZN(mask08[4]) );
  AND2_X1 U136 ( .A1(n80), .A2(op[4]), .ZN(mask00[4]) );
  INV_X1 U137 ( .A(n64), .ZN(mask08[5]) );
  AND2_X1 U138 ( .A1(n80), .A2(op[5]), .ZN(mask00[5]) );
  INV_X1 U139 ( .A(op[22]), .ZN(n351) );
  INV_X1 U140 ( .A(op[20]), .ZN(n355) );
  INV_X1 U141 ( .A(op[21]), .ZN(n353) );
  INV_X1 U142 ( .A(op[16]), .ZN(n363) );
  INV_X1 U143 ( .A(op[18]), .ZN(n359) );
  INV_X1 U144 ( .A(op[17]), .ZN(n361) );
  INV_X1 U145 ( .A(op[19]), .ZN(n357) );
  INV_X1 U146 ( .A(op[23]), .ZN(n349) );
  NAND2_X1 U147 ( .A1(op[9]), .A2(n80), .ZN(n68) );
  NAND2_X1 U148 ( .A1(op[12]), .A2(n80), .ZN(n65) );
  NAND2_X1 U149 ( .A1(op[14]), .A2(n80), .ZN(n63) );
  NAND2_X1 U150 ( .A1(op[10]), .A2(n80), .ZN(n67) );
  INV_X1 U151 ( .A(n66), .ZN(mask08[3]) );
  AND2_X1 U152 ( .A1(n80), .A2(op[3]), .ZN(mask00[3]) );
  INV_X1 U153 ( .A(n67), .ZN(mask08[2]) );
  AND2_X1 U154 ( .A1(n80), .A2(op[2]), .ZN(mask00[2]) );
  INV_X1 U155 ( .A(n69), .ZN(mask08[0]) );
  AND2_X1 U156 ( .A1(n80), .A2(op[0]), .ZN(mask00[0]) );
  INV_X1 U157 ( .A(op[14]), .ZN(n366) );
  INV_X1 U158 ( .A(op[15]), .ZN(n364) );
  INV_X1 U159 ( .A(op[12]), .ZN(n370) );
  INV_X1 U160 ( .A(op[13]), .ZN(n368) );
  INV_X1 U162 ( .A(op[10]), .ZN(n374) );
  INV_X1 U163 ( .A(op[9]), .ZN(n376) );
  INV_X1 U164 ( .A(op[11]), .ZN(n372) );
  INV_X1 U165 ( .A(op[7]), .ZN(n379) );
  INV_X1 U166 ( .A(op[28]), .ZN(n338) );
  INV_X1 U167 ( .A(op[29]), .ZN(n336) );
  INV_X1 U168 ( .A(op[25]), .ZN(n344) );
  INV_X1 U169 ( .A(n80), .ZN(n329) );
endmodule


module COARSE_SHIFT ( SEL, MASK00, MASK08, MASK16, Y );
  input [1:0] SEL;
  input [38:0] MASK00;
  input [38:0] MASK08;
  input [38:0] MASK16;
  output [38:0] Y;
  wire   n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n374;

  BUF_X1 U2 ( .A(n323), .Z(n326) );
  BUF_X1 U3 ( .A(n323), .Z(n325) );
  BUF_X1 U4 ( .A(n324), .Z(n327) );
  BUF_X1 U5 ( .A(n317), .Z(n320) );
  BUF_X1 U6 ( .A(n317), .Z(n319) );
  BUF_X1 U7 ( .A(n318), .Z(n321) );
  BUF_X1 U8 ( .A(n329), .Z(n332) );
  BUF_X1 U9 ( .A(n329), .Z(n331) );
  BUF_X1 U10 ( .A(n330), .Z(n333) );
  BUF_X1 U11 ( .A(n330), .Z(n334) );
  BUF_X1 U12 ( .A(n324), .Z(n328) );
  BUF_X1 U13 ( .A(n318), .Z(n322) );
  INV_X1 U14 ( .A(n75), .ZN(Y[1]) );
  INV_X1 U15 ( .A(n41), .ZN(Y[37]) );
  AOI222_X1 U16 ( .A1(MASK00[37]), .A2(n334), .B1(MASK16[37]), .B2(n328), .C1(
        MASK08[37]), .C2(n322), .ZN(n41) );
  INV_X1 U17 ( .A(n55), .ZN(Y[38]) );
  AOI222_X1 U18 ( .A1(MASK00[38]), .A2(n333), .B1(MASK16[38]), .B2(n327), .C1(
        MASK08[38]), .C2(n321), .ZN(n55) );
  INV_X1 U19 ( .A(n67), .ZN(Y[8]) );
  AOI222_X1 U20 ( .A1(MASK00[8]), .A2(n332), .B1(MASK16[8]), .B2(n326), .C1(
        MASK08[8]), .C2(n320), .ZN(n67) );
  INV_X1 U21 ( .A(n68), .ZN(Y[9]) );
  AOI222_X1 U22 ( .A1(MASK00[9]), .A2(n332), .B1(MASK16[9]), .B2(n326), .C1(
        MASK08[9]), .C2(n320), .ZN(n68) );
  INV_X1 U23 ( .A(n69), .ZN(Y[10]) );
  AOI222_X1 U24 ( .A1(MASK00[10]), .A2(n332), .B1(MASK16[10]), .B2(n326), .C1(
        MASK08[10]), .C2(n320), .ZN(n69) );
  INV_X1 U25 ( .A(n77), .ZN(Y[11]) );
  AOI222_X1 U26 ( .A1(MASK00[11]), .A2(n331), .B1(MASK16[11]), .B2(n325), .C1(
        MASK08[11]), .C2(n319), .ZN(n77) );
  INV_X1 U27 ( .A(n66), .ZN(Y[7]) );
  AOI222_X1 U28 ( .A1(MASK00[7]), .A2(n332), .B1(MASK16[7]), .B2(n326), .C1(
        MASK08[7]), .C2(n320), .ZN(n66) );
  INV_X1 U29 ( .A(n81), .ZN(Y[12]) );
  AOI222_X1 U30 ( .A1(MASK00[12]), .A2(n331), .B1(MASK16[12]), .B2(n325), .C1(
        MASK08[12]), .C2(n319), .ZN(n81) );
  INV_X1 U31 ( .A(n82), .ZN(Y[13]) );
  AOI222_X1 U32 ( .A1(MASK00[13]), .A2(n331), .B1(MASK16[13]), .B2(n325), .C1(
        MASK08[13]), .C2(n319), .ZN(n82) );
  INV_X1 U33 ( .A(n78), .ZN(Y[14]) );
  AOI222_X1 U34 ( .A1(MASK00[14]), .A2(n331), .B1(MASK16[14]), .B2(n325), .C1(
        MASK08[14]), .C2(n319), .ZN(n78) );
  INV_X1 U35 ( .A(n79), .ZN(Y[24]) );
  AOI222_X1 U36 ( .A1(MASK00[24]), .A2(n331), .B1(MASK16[24]), .B2(n325), .C1(
        MASK08[24]), .C2(n319), .ZN(n79) );
  INV_X1 U37 ( .A(n80), .ZN(Y[25]) );
  AOI222_X1 U38 ( .A1(MASK00[25]), .A2(n331), .B1(MASK16[25]), .B2(n325), .C1(
        MASK08[25]), .C2(n319), .ZN(n80) );
  INV_X1 U39 ( .A(n70), .ZN(Y[26]) );
  AOI222_X1 U40 ( .A1(MASK00[26]), .A2(n332), .B1(MASK16[26]), .B2(n326), .C1(
        MASK08[26]), .C2(n320), .ZN(n70) );
  INV_X1 U41 ( .A(n71), .ZN(Y[27]) );
  AOI222_X1 U42 ( .A1(MASK00[27]), .A2(n332), .B1(MASK16[27]), .B2(n325), .C1(
        MASK08[27]), .C2(n319), .ZN(n71) );
  INV_X1 U43 ( .A(n72), .ZN(Y[28]) );
  AOI222_X1 U44 ( .A1(MASK00[28]), .A2(n331), .B1(MASK16[28]), .B2(n325), .C1(
        MASK08[28]), .C2(n319), .ZN(n72) );
  INV_X1 U45 ( .A(n73), .ZN(Y[29]) );
  AOI222_X1 U46 ( .A1(MASK00[29]), .A2(n331), .B1(MASK16[29]), .B2(n325), .C1(
        MASK08[29]), .C2(n319), .ZN(n73) );
  INV_X1 U47 ( .A(n74), .ZN(Y[30]) );
  AOI222_X1 U48 ( .A1(MASK00[30]), .A2(n331), .B1(MASK16[30]), .B2(n325), .C1(
        MASK08[30]), .C2(n319), .ZN(n74) );
  INV_X1 U49 ( .A(n56), .ZN(Y[15]) );
  AOI222_X1 U50 ( .A1(MASK00[15]), .A2(n333), .B1(MASK16[15]), .B2(n327), .C1(
        MASK08[15]), .C2(n321), .ZN(n56) );
  INV_X1 U51 ( .A(n47), .ZN(Y[18]) );
  AOI222_X1 U52 ( .A1(MASK00[18]), .A2(n334), .B1(MASK16[18]), .B2(n327), .C1(
        MASK08[18]), .C2(n321), .ZN(n47) );
  INV_X1 U53 ( .A(n48), .ZN(Y[19]) );
  AOI222_X1 U54 ( .A1(MASK00[19]), .A2(n334), .B1(MASK16[19]), .B2(n327), .C1(
        MASK08[19]), .C2(n321), .ZN(n48) );
  INV_X1 U55 ( .A(n49), .ZN(Y[20]) );
  AOI222_X1 U56 ( .A1(MASK00[20]), .A2(n334), .B1(MASK16[20]), .B2(n327), .C1(
        MASK08[20]), .C2(n321), .ZN(n49) );
  INV_X1 U57 ( .A(n57), .ZN(Y[21]) );
  AOI222_X1 U58 ( .A1(MASK00[21]), .A2(n333), .B1(MASK16[21]), .B2(n327), .C1(
        MASK08[21]), .C2(n321), .ZN(n57) );
  INV_X1 U59 ( .A(n58), .ZN(Y[22]) );
  AOI222_X1 U60 ( .A1(MASK00[22]), .A2(n333), .B1(MASK16[22]), .B2(n327), .C1(
        MASK08[22]), .C2(n321), .ZN(n58) );
  INV_X1 U61 ( .A(n59), .ZN(Y[23]) );
  AOI222_X1 U62 ( .A1(MASK00[23]), .A2(n333), .B1(MASK16[23]), .B2(n326), .C1(
        MASK08[23]), .C2(n320), .ZN(n59) );
  INV_X1 U63 ( .A(n60), .ZN(Y[33]) );
  AOI222_X1 U64 ( .A1(MASK00[33]), .A2(n333), .B1(MASK16[33]), .B2(n326), .C1(
        MASK08[33]), .C2(n320), .ZN(n60) );
  INV_X1 U65 ( .A(n45), .ZN(Y[16]) );
  AOI222_X1 U66 ( .A1(MASK00[16]), .A2(n334), .B1(MASK16[16]), .B2(n328), .C1(
        MASK08[16]), .C2(n322), .ZN(n45) );
  INV_X1 U67 ( .A(n46), .ZN(Y[17]) );
  AOI222_X1 U68 ( .A1(MASK00[17]), .A2(n334), .B1(MASK16[17]), .B2(n328), .C1(
        MASK08[17]), .C2(n322), .ZN(n46) );
  INV_X1 U69 ( .A(n61), .ZN(Y[34]) );
  AOI222_X1 U70 ( .A1(MASK00[34]), .A2(n332), .B1(MASK16[34]), .B2(n326), .C1(
        MASK08[34]), .C2(n320), .ZN(n61) );
  INV_X1 U71 ( .A(n64), .ZN(Y[31]) );
  AOI222_X1 U72 ( .A1(MASK00[31]), .A2(n332), .B1(MASK16[31]), .B2(n326), .C1(
        MASK08[31]), .C2(n320), .ZN(n64) );
  INV_X1 U73 ( .A(n65), .ZN(Y[32]) );
  AOI222_X1 U74 ( .A1(MASK00[32]), .A2(n332), .B1(MASK16[32]), .B2(n326), .C1(
        MASK08[32]), .C2(n320), .ZN(n65) );
  INV_X1 U75 ( .A(n63), .ZN(Y[36]) );
  AOI222_X1 U76 ( .A1(MASK00[36]), .A2(n332), .B1(MASK16[36]), .B2(n326), .C1(
        MASK08[36]), .C2(n320), .ZN(n63) );
  INV_X1 U77 ( .A(n62), .ZN(Y[35]) );
  AOI222_X1 U78 ( .A1(MASK00[35]), .A2(n332), .B1(MASK16[35]), .B2(n326), .C1(
        MASK08[35]), .C2(n320), .ZN(n62) );
  BUF_X1 U79 ( .A(n42), .Z(n329) );
  BUF_X1 U80 ( .A(n43), .Z(n323) );
  BUF_X1 U81 ( .A(n44), .Z(n317) );
  BUF_X1 U82 ( .A(n42), .Z(n330) );
  BUF_X1 U83 ( .A(n43), .Z(n324) );
  BUF_X1 U84 ( .A(n44), .Z(n318) );
  AOI222_X1 U85 ( .A1(MASK00[1]), .A2(n331), .B1(MASK16[1]), .B2(n325), .C1(
        MASK08[1]), .C2(n319), .ZN(n75) );
  INV_X1 U86 ( .A(n50), .ZN(Y[6]) );
  AOI222_X1 U87 ( .A1(MASK00[6]), .A2(n333), .B1(MASK16[6]), .B2(n327), .C1(
        MASK08[6]), .C2(n321), .ZN(n50) );
  NOR2_X1 U88 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n42) );
  INV_X1 U89 ( .A(n51), .ZN(Y[4]) );
  AOI222_X1 U90 ( .A1(MASK00[4]), .A2(n333), .B1(MASK16[4]), .B2(n327), .C1(
        MASK08[4]), .C2(n321), .ZN(n51) );
  INV_X1 U91 ( .A(n52), .ZN(Y[5]) );
  AOI222_X1 U92 ( .A1(MASK00[5]), .A2(n333), .B1(MASK16[5]), .B2(n327), .C1(
        MASK08[5]), .C2(n321), .ZN(n52) );
  NOR2_X1 U93 ( .A1(n374), .A2(SEL[0]), .ZN(n43) );
  INV_X1 U94 ( .A(n54), .ZN(Y[3]) );
  AOI222_X1 U95 ( .A1(MASK00[3]), .A2(n333), .B1(MASK16[3]), .B2(n327), .C1(
        MASK08[3]), .C2(n321), .ZN(n54) );
  INV_X1 U96 ( .A(n53), .ZN(Y[2]) );
  AOI222_X1 U97 ( .A1(MASK00[2]), .A2(n333), .B1(MASK16[2]), .B2(n327), .C1(
        MASK08[2]), .C2(n321), .ZN(n53) );
  INV_X1 U98 ( .A(n76), .ZN(Y[0]) );
  AOI222_X1 U99 ( .A1(MASK00[0]), .A2(n331), .B1(MASK16[0]), .B2(n325), .C1(
        MASK08[0]), .C2(n319), .ZN(n76) );
  INV_X1 U100 ( .A(SEL[1]), .ZN(n374) );
  AND2_X1 U101 ( .A1(SEL[0]), .A2(n374), .ZN(n44) );
endmodule


module FINE_SHIFT ( op, sel, shifted );
  input [38:0] op;
  input [2:0] sel;
  output [31:0] shifted;
  wire   n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413;

  AND2_X1 U1 ( .A1(sel[2]), .A2(sel[1]), .ZN(n359) );
  INV_X1 U2 ( .A(n362), .ZN(n360) );
  INV_X1 U3 ( .A(n362), .ZN(n361) );
  INV_X1 U4 ( .A(n368), .ZN(n367) );
  INV_X1 U5 ( .A(n359), .ZN(n366) );
  INV_X1 U6 ( .A(n359), .ZN(n365) );
  INV_X1 U7 ( .A(n364), .ZN(n363) );
  OAI221_X1 U8 ( .B1(op[13]), .B2(n43), .C1(op[11]), .C2(n365), .A(n106), .ZN(
        n103) );
  AOI22_X1 U9 ( .A1(n46), .A2(n388), .B1(n360), .B2(n380), .ZN(n106) );
  OAI221_X1 U10 ( .B1(op[12]), .B2(n43), .C1(op[10]), .C2(n365), .A(n105), 
        .ZN(n40) );
  AOI22_X1 U11 ( .A1(n46), .A2(n389), .B1(n47), .B2(n402), .ZN(n105) );
  OAI221_X1 U12 ( .B1(op[14]), .B2(n43), .C1(op[12]), .C2(n366), .A(n104), 
        .ZN(n101) );
  AOI22_X1 U13 ( .A1(n46), .A2(n387), .B1(n361), .B2(n389), .ZN(n104) );
  OAI221_X1 U14 ( .B1(op[15]), .B2(n43), .C1(op[13]), .C2(n365), .A(n102), 
        .ZN(n99) );
  AOI22_X1 U15 ( .A1(n363), .A2(n386), .B1(n361), .B2(n388), .ZN(n102) );
  OAI221_X1 U16 ( .B1(op[16]), .B2(n43), .C1(op[14]), .C2(n366), .A(n100), 
        .ZN(n97) );
  AOI22_X1 U17 ( .A1(n363), .A2(n385), .B1(n361), .B2(n387), .ZN(n100) );
  OAI221_X1 U18 ( .B1(op[17]), .B2(n43), .C1(op[15]), .C2(n365), .A(n98), .ZN(
        n95) );
  AOI22_X1 U19 ( .A1(n363), .A2(n384), .B1(n361), .B2(n386), .ZN(n98) );
  OAI221_X1 U20 ( .B1(op[18]), .B2(n43), .C1(op[16]), .C2(n366), .A(n96), .ZN(
        n93) );
  AOI22_X1 U21 ( .A1(n363), .A2(n383), .B1(n361), .B2(n385), .ZN(n96) );
  OAI221_X1 U22 ( .B1(op[9]), .B2(n367), .C1(op[7]), .C2(n365), .A(n51), .ZN(
        n48) );
  AOI22_X1 U23 ( .A1(n46), .A2(n403), .B1(n360), .B2(n405), .ZN(n51) );
  INV_X1 U24 ( .A(op[11]), .ZN(n405) );
  OAI221_X1 U25 ( .B1(op[10]), .B2(n367), .C1(op[8]), .C2(n365), .A(n49), .ZN(
        n42) );
  AOI22_X1 U26 ( .A1(n46), .A2(n402), .B1(n360), .B2(n404), .ZN(n49) );
  OAI221_X1 U27 ( .B1(op[19]), .B2(n43), .C1(op[17]), .C2(n365), .A(n94), .ZN(
        n91) );
  AOI22_X1 U28 ( .A1(n363), .A2(n382), .B1(n361), .B2(n384), .ZN(n94) );
  OAI221_X1 U29 ( .B1(op[20]), .B2(n43), .C1(op[18]), .C2(n366), .A(n92), .ZN(
        n89) );
  AOI22_X1 U30 ( .A1(n363), .A2(n395), .B1(n361), .B2(n383), .ZN(n92) );
  OAI221_X1 U31 ( .B1(op[21]), .B2(n43), .C1(op[19]), .C2(n366), .A(n90), .ZN(
        n87) );
  AOI22_X1 U32 ( .A1(n363), .A2(n396), .B1(n361), .B2(n382), .ZN(n90) );
  OAI221_X1 U33 ( .B1(op[22]), .B2(n43), .C1(op[20]), .C2(n366), .A(n88), .ZN(
        n83) );
  AOI22_X1 U34 ( .A1(n363), .A2(n397), .B1(n361), .B2(n395), .ZN(n88) );
  OAI221_X1 U35 ( .B1(op[23]), .B2(n367), .C1(op[21]), .C2(n366), .A(n84), 
        .ZN(n81) );
  AOI22_X1 U36 ( .A1(n363), .A2(n398), .B1(n361), .B2(n396), .ZN(n84) );
  OAI221_X1 U37 ( .B1(op[24]), .B2(n43), .C1(op[22]), .C2(n366), .A(n82), .ZN(
        n79) );
  AOI22_X1 U38 ( .A1(n363), .A2(n399), .B1(n361), .B2(n397), .ZN(n82) );
  OAI221_X1 U39 ( .B1(op[25]), .B2(n367), .C1(op[23]), .C2(n366), .A(n80), 
        .ZN(n77) );
  AOI22_X1 U40 ( .A1(n46), .A2(n400), .B1(n361), .B2(n398), .ZN(n80) );
  OAI221_X1 U41 ( .B1(op[26]), .B2(n43), .C1(op[24]), .C2(n366), .A(n78), .ZN(
        n75) );
  AOI22_X1 U42 ( .A1(n46), .A2(n401), .B1(n360), .B2(n399), .ZN(n78) );
  OAI221_X1 U43 ( .B1(op[27]), .B2(n367), .C1(op[25]), .C2(n366), .A(n76), 
        .ZN(n73) );
  AOI22_X1 U44 ( .A1(n46), .A2(n381), .B1(n360), .B2(n400), .ZN(n76) );
  OAI221_X1 U45 ( .B1(op[28]), .B2(n43), .C1(op[26]), .C2(n366), .A(n74), .ZN(
        n71) );
  AOI22_X1 U46 ( .A1(n363), .A2(n390), .B1(n360), .B2(n401), .ZN(n74) );
  OAI221_X1 U47 ( .B1(op[29]), .B2(n367), .C1(op[27]), .C2(n365), .A(n72), 
        .ZN(n69) );
  AOI22_X1 U48 ( .A1(n363), .A2(n391), .B1(n360), .B2(n381), .ZN(n72) );
  OAI221_X1 U49 ( .B1(op[30]), .B2(n367), .C1(op[28]), .C2(n365), .A(n70), 
        .ZN(n67) );
  AOI22_X1 U50 ( .A1(n363), .A2(n392), .B1(n360), .B2(n390), .ZN(n70) );
  OAI221_X1 U51 ( .B1(op[31]), .B2(n367), .C1(op[29]), .C2(n365), .A(n68), 
        .ZN(n65) );
  AOI22_X1 U52 ( .A1(n363), .A2(n393), .B1(n360), .B2(n391), .ZN(n68) );
  INV_X1 U53 ( .A(op[35]), .ZN(n393) );
  OAI221_X1 U54 ( .B1(op[32]), .B2(n367), .C1(op[30]), .C2(n365), .A(n66), 
        .ZN(n61) );
  AOI22_X1 U55 ( .A1(n363), .A2(n394), .B1(n360), .B2(n392), .ZN(n66) );
  INV_X1 U56 ( .A(op[36]), .ZN(n394) );
  OAI221_X1 U57 ( .B1(op[11]), .B2(n367), .C1(op[9]), .C2(n365), .A(n45), .ZN(
        n41) );
  AOI22_X1 U58 ( .A1(n363), .A2(n380), .B1(n361), .B2(n403), .ZN(n45) );
  INV_X1 U59 ( .A(op[31]), .ZN(n381) );
  INV_X1 U60 ( .A(op[32]), .ZN(n390) );
  BUF_X1 U61 ( .A(n379), .Z(n370) );
  BUF_X1 U62 ( .A(n378), .Z(n371) );
  BUF_X1 U63 ( .A(n379), .Z(n377) );
  BUF_X1 U64 ( .A(n379), .Z(n376) );
  BUF_X1 U65 ( .A(n379), .Z(n375) );
  BUF_X1 U66 ( .A(n378), .Z(n373) );
  BUF_X1 U67 ( .A(n370), .Z(n374) );
  BUF_X1 U68 ( .A(n379), .Z(n372) );
  BUF_X1 U69 ( .A(n379), .Z(n378) );
  INV_X1 U70 ( .A(op[12]), .ZN(n404) );
  INV_X1 U71 ( .A(op[13]), .ZN(n403) );
  INV_X1 U72 ( .A(op[14]), .ZN(n402) );
  INV_X1 U73 ( .A(op[15]), .ZN(n380) );
  INV_X1 U74 ( .A(op[16]), .ZN(n389) );
  INV_X1 U75 ( .A(op[17]), .ZN(n388) );
  INV_X1 U76 ( .A(op[18]), .ZN(n387) );
  INV_X1 U77 ( .A(op[19]), .ZN(n386) );
  INV_X1 U78 ( .A(op[20]), .ZN(n385) );
  INV_X1 U79 ( .A(op[21]), .ZN(n384) );
  INV_X1 U80 ( .A(op[22]), .ZN(n383) );
  INV_X1 U81 ( .A(op[23]), .ZN(n382) );
  INV_X1 U82 ( .A(op[24]), .ZN(n395) );
  INV_X1 U83 ( .A(op[25]), .ZN(n396) );
  INV_X1 U84 ( .A(op[26]), .ZN(n397) );
  INV_X1 U85 ( .A(op[27]), .ZN(n398) );
  INV_X1 U86 ( .A(op[28]), .ZN(n399) );
  INV_X1 U87 ( .A(op[29]), .ZN(n400) );
  INV_X1 U88 ( .A(op[30]), .ZN(n401) );
  OAI22_X1 U89 ( .A1(n376), .A2(n93), .B1(n369), .B2(n91), .ZN(shifted[16]) );
  OAI22_X1 U90 ( .A1(n376), .A2(n91), .B1(sel[0]), .B2(n89), .ZN(shifted[17])
         );
  OAI22_X1 U91 ( .A1(n376), .A2(n89), .B1(n369), .B2(n87), .ZN(shifted[18]) );
  OAI22_X1 U92 ( .A1(n373), .A2(n69), .B1(sel[0]), .B2(n67), .ZN(shifted[27])
         );
  OAI22_X1 U93 ( .A1(n373), .A2(n67), .B1(n369), .B2(n65), .ZN(shifted[28]) );
  OAI22_X1 U94 ( .A1(n372), .A2(n65), .B1(sel[0]), .B2(n61), .ZN(shifted[29])
         );
  OAI22_X1 U95 ( .A1(n374), .A2(n61), .B1(n369), .B2(n58), .ZN(shifted[30]) );
  OAI22_X1 U96 ( .A1(n372), .A2(n58), .B1(n369), .B2(n59), .ZN(shifted[31]) );
  OAI22_X1 U97 ( .A1(n375), .A2(n87), .B1(n369), .B2(n83), .ZN(shifted[19]) );
  OAI22_X1 U98 ( .A1(n375), .A2(n83), .B1(n369), .B2(n81), .ZN(shifted[20]) );
  OAI22_X1 U99 ( .A1(n375), .A2(n81), .B1(n369), .B2(n79), .ZN(shifted[21]) );
  OAI22_X1 U100 ( .A1(n374), .A2(n79), .B1(n369), .B2(n77), .ZN(shifted[22])
         );
  OAI22_X1 U101 ( .A1(n374), .A2(n77), .B1(n369), .B2(n75), .ZN(shifted[23])
         );
  OAI22_X1 U102 ( .A1(n374), .A2(n75), .B1(n369), .B2(n73), .ZN(shifted[24])
         );
  OAI22_X1 U103 ( .A1(n373), .A2(n73), .B1(n369), .B2(n71), .ZN(shifted[25])
         );
  OAI22_X1 U104 ( .A1(n373), .A2(n71), .B1(n369), .B2(n69), .ZN(shifted[26])
         );
  OAI22_X1 U105 ( .A1(n375), .A2(n85), .B1(n369), .B2(n63), .ZN(shifted[1]) );
  OAI22_X1 U106 ( .A1(n372), .A2(n56), .B1(sel[0]), .B2(n54), .ZN(shifted[3])
         );
  OAI22_X1 U107 ( .A1(n371), .A2(n48), .B1(n369), .B2(n42), .ZN(shifted[7]) );
  OAI22_X1 U108 ( .A1(n377), .A2(n103), .B1(n369), .B2(n101), .ZN(shifted[11])
         );
  OAI22_X1 U109 ( .A1(n377), .A2(n99), .B1(sel[0]), .B2(n97), .ZN(shifted[13])
         );
  OAI22_X1 U110 ( .A1(n376), .A2(n95), .B1(n369), .B2(n93), .ZN(shifted[15])
         );
  OAI22_X1 U111 ( .A1(n371), .A2(n52), .B1(sel[0]), .B2(n50), .ZN(shifted[5])
         );
  OAI22_X1 U112 ( .A1(sel[0]), .A2(n40), .B1(n41), .B2(n370), .ZN(shifted[9])
         );
  OAI221_X1 U113 ( .B1(op[3]), .B2(n367), .C1(op[1]), .C2(n365), .A(n411), 
        .ZN(n85) );
  INV_X1 U114 ( .A(n109), .ZN(n411) );
  OAI22_X1 U115 ( .A1(n364), .A2(op[7]), .B1(n362), .B2(op[5]), .ZN(n109) );
  OAI221_X1 U116 ( .B1(op[4]), .B2(n43), .C1(op[2]), .C2(n366), .A(n410), .ZN(
        n63) );
  INV_X1 U117 ( .A(n86), .ZN(n410) );
  OAI22_X1 U118 ( .A1(n364), .A2(op[8]), .B1(n362), .B2(op[6]), .ZN(n86) );
  OAI221_X1 U119 ( .B1(op[5]), .B2(n367), .C1(op[3]), .C2(n365), .A(n409), 
        .ZN(n56) );
  INV_X1 U120 ( .A(n64), .ZN(n409) );
  OAI22_X1 U121 ( .A1(n364), .A2(op[9]), .B1(n362), .B2(op[7]), .ZN(n64) );
  OAI221_X1 U122 ( .B1(op[6]), .B2(n367), .C1(op[4]), .C2(n365), .A(n408), 
        .ZN(n54) );
  INV_X1 U123 ( .A(n57), .ZN(n408) );
  OAI22_X1 U124 ( .A1(n364), .A2(op[10]), .B1(n362), .B2(op[8]), .ZN(n57) );
  OAI221_X1 U125 ( .B1(op[7]), .B2(n367), .C1(op[5]), .C2(n365), .A(n406), 
        .ZN(n52) );
  INV_X1 U126 ( .A(n55), .ZN(n406) );
  OAI22_X1 U127 ( .A1(n364), .A2(op[11]), .B1(n362), .B2(op[9]), .ZN(n55) );
  OAI221_X1 U128 ( .B1(op[8]), .B2(n367), .C1(op[6]), .C2(n366), .A(n53), .ZN(
        n50) );
  AOI22_X1 U129 ( .A1(n363), .A2(n404), .B1(n360), .B2(n407), .ZN(n53) );
  INV_X1 U130 ( .A(op[10]), .ZN(n407) );
  OAI221_X1 U131 ( .B1(op[37]), .B2(n364), .C1(op[35]), .C2(n362), .A(n62), 
        .ZN(n58) );
  AOI22_X1 U132 ( .A1(n368), .A2(n391), .B1(n359), .B2(n381), .ZN(n62) );
  AOI221_X1 U133 ( .B1(op[38]), .B2(n46), .C1(op[36]), .C2(n360), .A(n60), 
        .ZN(n59) );
  OAI22_X1 U134 ( .A1(n366), .A2(n390), .B1(n367), .B2(n392), .ZN(n60) );
  NOR2_X1 U135 ( .A1(n413), .A2(sel[2]), .ZN(n47) );
  NOR2_X1 U136 ( .A1(sel[1]), .A2(sel[2]), .ZN(n46) );
  NAND2_X1 U137 ( .A1(sel[2]), .A2(n413), .ZN(n43) );
  INV_X1 U138 ( .A(sel[1]), .ZN(n413) );
  INV_X1 U139 ( .A(op[33]), .ZN(n391) );
  INV_X1 U140 ( .A(op[34]), .ZN(n392) );
  INV_X1 U141 ( .A(n108), .ZN(n412) );
  AOI22_X1 U142 ( .A1(n360), .A2(op[4]), .B1(n46), .B2(op[6]), .ZN(n108) );
  INV_X1 U143 ( .A(n369), .ZN(n379) );
  OAI22_X1 U144 ( .A1(n372), .A2(n63), .B1(n369), .B2(n56), .ZN(shifted[2]) );
  OAI22_X1 U145 ( .A1(n371), .A2(n54), .B1(sel[0]), .B2(n52), .ZN(shifted[4])
         );
  OAI22_X1 U146 ( .A1(n369), .A2(n103), .B1(n370), .B2(n40), .ZN(shifted[10])
         );
  OAI22_X1 U147 ( .A1(n377), .A2(n101), .B1(sel[0]), .B2(n99), .ZN(shifted[12]) );
  OAI22_X1 U148 ( .A1(n377), .A2(n97), .B1(n369), .B2(n95), .ZN(shifted[14])
         );
  OAI22_X1 U149 ( .A1(n371), .A2(n50), .B1(n369), .B2(n48), .ZN(shifted[6]) );
  OAI22_X1 U150 ( .A1(n370), .A2(n42), .B1(n369), .B2(n41), .ZN(shifted[8]) );
  OAI22_X1 U151 ( .A1(sel[0]), .A2(n85), .B1(n107), .B2(n370), .ZN(shifted[0])
         );
  AOI221_X1 U152 ( .B1(op[2]), .B2(n368), .C1(op[0]), .C2(n359), .A(n412), 
        .ZN(n107) );
  BUF_X1 U153 ( .A(sel[0]), .Z(n369) );
  INV_X1 U154 ( .A(n47), .ZN(n362) );
  INV_X1 U155 ( .A(n46), .ZN(n364) );
  INV_X1 U156 ( .A(n43), .ZN(n368) );
endmodule


module SHIFTER_WIDTH32 ( R1, R2, SEL, Y );
  input [31:0] R1;
  input [31:0] R2;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n2, n3, n4, n1;
  wire   [38:0] m0;
  wire   [38:0] m8;
  wire   [38:0] m16;
  wire   [38:0] y2;

  XOR2_X1 U2 ( .A(n1), .B(R2[0]), .Z(n4) );
  XOR2_X1 U3 ( .A(n1), .B(R2[1]), .Z(n3) );
  XOR2_X1 U4 ( .A(n1), .B(R2[2]), .Z(n2) );
  MASK_GENERATOR level_1 ( .op(R1), .sel(SEL), .mask00(m0), .mask08(m8), 
        .mask16(m16) );
  COARSE_SHIFT level_2 ( .SEL(R2[4:3]), .MASK00(m0), .MASK08(m8), .MASK16(m16), 
        .Y(y2) );
  FINE_SHIFT level_3 ( .op(y2), .sel({n2, n3, n4}), .shifted(Y) );
  OR2_X1 U1 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n1) );
endmodule


module BOOTH_ENCODER_WIDTH16_0 ( A, b, vp );
  input [15:0] A;
  input [2:0] b;
  output [16:0] vp;
  wire   \notA[0] , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184;
  assign \notA[0]  = A[0];

  XOR2_X1 U90 ( .A(n31), .B(A[9]), .Z(n21) );
  NAND3_X1 U91 ( .A1(n176), .A2(n165), .A3(n31), .ZN(n68) );
  NOR2_X2 U3 ( .A1(n71), .A2(b[2]), .ZN(n26) );
  NOR2_X2 U4 ( .A1(n70), .A2(b[2]), .ZN(n29) );
  INV_X1 U5 ( .A(n62), .ZN(n173) );
  INV_X1 U6 ( .A(n24), .ZN(n169) );
  OAI21_X1 U7 ( .B1(n64), .B2(n166), .A(n62), .ZN(n60) );
  OAI21_X1 U8 ( .B1(n173), .B2(n167), .A(n57), .ZN(n58) );
  NAND2_X1 U9 ( .A1(n173), .A2(n167), .ZN(n57) );
  INV_X1 U10 ( .A(n49), .ZN(n181) );
  INV_X1 U11 ( .A(n40), .ZN(n179) );
  NAND2_X1 U12 ( .A1(n64), .A2(n166), .ZN(n62) );
  OAI221_X1 U13 ( .B1(n22), .B2(n41), .C1(n169), .C2(n182), .A(n44), .ZN(vp[3]) );
  AOI22_X1 U14 ( .A1(A[2]), .A2(n26), .B1(A[3]), .B2(n29), .ZN(n44) );
  OAI221_X1 U15 ( .B1(n22), .B2(n36), .C1(n169), .C2(n41), .A(n42), .ZN(vp[4])
         );
  AOI22_X1 U16 ( .A1(A[3]), .A2(n26), .B1(A[4]), .B2(n29), .ZN(n42) );
  OAI221_X1 U17 ( .B1(n22), .B2(n180), .C1(n169), .C2(n36), .A(n37), .ZN(vp[5]) );
  AOI22_X1 U18 ( .A1(A[4]), .A2(n26), .B1(A[5]), .B2(n29), .ZN(n37) );
  OAI221_X1 U19 ( .B1(n22), .B2(n32), .C1(n169), .C2(n180), .A(n35), .ZN(vp[6]) );
  AOI22_X1 U20 ( .A1(A[5]), .A2(n26), .B1(A[6]), .B2(n29), .ZN(n35) );
  OAI221_X1 U21 ( .B1(n22), .B2(n27), .C1(n169), .C2(n32), .A(n33), .ZN(vp[7])
         );
  AOI22_X1 U22 ( .A1(A[6]), .A2(n26), .B1(A[7]), .B2(n29), .ZN(n33) );
  OAI221_X1 U23 ( .B1(n22), .B2(n66), .C1(n171), .C2(n176), .A(n168), .ZN(
        vp[10]) );
  INV_X1 U24 ( .A(n69), .ZN(n168) );
  OAI22_X1 U25 ( .A1(n165), .A2(n172), .B1(n21), .B2(n169), .ZN(n69) );
  OAI221_X1 U26 ( .B1(n22), .B2(n60), .C1(n169), .C2(n174), .A(n63), .ZN(
        vp[12]) );
  AOI22_X1 U27 ( .A1(A[11]), .A2(n26), .B1(A[12]), .B2(n29), .ZN(n63) );
  OAI221_X1 U28 ( .B1(n22), .B2(n58), .C1(n169), .C2(n60), .A(n61), .ZN(vp[13]) );
  AOI22_X1 U29 ( .A1(A[12]), .A2(n26), .B1(A[13]), .B2(n29), .ZN(n61) );
  OAI221_X1 U30 ( .B1(n22), .B2(n54), .C1(n169), .C2(n58), .A(n59), .ZN(vp[14]) );
  AOI22_X1 U31 ( .A1(A[13]), .A2(n26), .B1(A[14]), .B2(n29), .ZN(n59) );
  OAI221_X1 U32 ( .B1(n22), .B2(n52), .C1(n169), .C2(n54), .A(n55), .ZN(vp[15]) );
  AOI22_X1 U33 ( .A1(A[14]), .A2(n26), .B1(A[15]), .B2(n29), .ZN(n55) );
  OAI221_X1 U34 ( .B1(n21), .B2(n22), .C1(n165), .C2(n171), .A(n23), .ZN(vp[9]) );
  AOI22_X1 U35 ( .A1(n24), .A2(n25), .B1(n26), .B2(A[8]), .ZN(n23) );
  OAI221_X1 U36 ( .B1(n178), .B2(n22), .C1(n169), .C2(n27), .A(n28), .ZN(vp[8]) );
  INV_X1 U37 ( .A(n25), .ZN(n178) );
  AOI22_X1 U38 ( .A1(A[7]), .A2(n26), .B1(n29), .B2(A[8]), .ZN(n28) );
  NOR2_X1 U39 ( .A1(n51), .A2(n170), .ZN(n24) );
  INV_X1 U40 ( .A(n70), .ZN(n170) );
  OR2_X1 U41 ( .A1(n70), .A2(n51), .ZN(n22) );
  NOR2_X1 U42 ( .A1(n30), .A2(A[8]), .ZN(n31) );
  AOI21_X1 U43 ( .B1(n30), .B2(A[8]), .A(n31), .ZN(n25) );
  OAI221_X1 U44 ( .B1(n22), .B2(n174), .C1(n172), .C2(n176), .A(n65), .ZN(
        vp[11]) );
  AOI22_X1 U45 ( .A1(n175), .A2(n24), .B1(A[11]), .B2(n29), .ZN(n65) );
  INV_X1 U46 ( .A(n66), .ZN(n175) );
  NOR2_X1 U47 ( .A1(n68), .A2(A[11]), .ZN(n64) );
  XNOR2_X1 U48 ( .A(n181), .B(A[3]), .ZN(n41) );
  XNOR2_X1 U49 ( .A(n179), .B(A[6]), .ZN(n32) );
  XOR2_X1 U50 ( .A(n164), .B(A[15]), .Z(n52) );
  NOR2_X1 U51 ( .A1(n57), .A2(A[14]), .ZN(n164) );
  XNOR2_X1 U52 ( .A(n57), .B(A[14]), .ZN(n54) );
  NOR2_X1 U53 ( .A1(n48), .A2(A[2]), .ZN(n49) );
  NOR2_X1 U54 ( .A1(n39), .A2(A[5]), .ZN(n40) );
  AOI21_X1 U55 ( .B1(n171), .B2(n22), .A(n184), .ZN(vp[0]) );
  OAI21_X1 U56 ( .B1(n183), .B2(n184), .A(n48), .ZN(n45) );
  OAI21_X1 U57 ( .B1(n51), .B2(n52), .A(n53), .ZN(vp[16]) );
  OAI21_X1 U58 ( .B1(n26), .B2(n29), .A(A[15]), .ZN(n53) );
  INV_X1 U59 ( .A(n29), .ZN(n171) );
  NAND2_X1 U60 ( .A1(n183), .A2(n184), .ZN(n48) );
  INV_X1 U61 ( .A(n26), .ZN(n172) );
  NAND2_X1 U62 ( .A1(n39), .A2(n43), .ZN(n36) );
  OAI21_X1 U63 ( .B1(A[3]), .B2(n181), .A(A[4]), .ZN(n43) );
  NAND2_X1 U64 ( .A1(n30), .A2(n34), .ZN(n27) );
  OAI21_X1 U65 ( .B1(A[6]), .B2(n179), .A(A[7]), .ZN(n34) );
  OR3_X1 U66 ( .A1(A[3]), .A2(A[4]), .A3(n181), .ZN(n39) );
  OR3_X1 U67 ( .A1(A[6]), .A2(A[7]), .A3(n179), .ZN(n30) );
  INV_X1 U68 ( .A(n47), .ZN(n182) );
  AOI21_X1 U69 ( .B1(n48), .B2(A[2]), .A(n49), .ZN(n47) );
  INV_X1 U70 ( .A(n38), .ZN(n180) );
  AOI21_X1 U71 ( .B1(n39), .B2(A[5]), .A(n40), .ZN(n38) );
  INV_X1 U72 ( .A(n67), .ZN(n174) );
  AOI21_X1 U73 ( .B1(n68), .B2(A[11]), .A(n64), .ZN(n67) );
  OAI21_X1 U74 ( .B1(b[1]), .B2(b[0]), .A(n71), .ZN(n70) );
  OAI221_X1 U75 ( .B1(n22), .B2(n45), .C1(n171), .C2(n183), .A(n50), .ZN(vp[1]) );
  OAI21_X1 U76 ( .B1(n26), .B2(n24), .A(\notA[0] ), .ZN(n50) );
  OAI221_X1 U77 ( .B1(n22), .B2(n182), .C1(n169), .C2(n45), .A(n46), .ZN(vp[2]) );
  AOI22_X1 U78 ( .A1(A[1]), .A2(n26), .B1(A[2]), .B2(n29), .ZN(n46) );
  INV_X1 U79 ( .A(\notA[0] ), .ZN(n184) );
  INV_X1 U80 ( .A(A[1]), .ZN(n183) );
  INV_X1 U81 ( .A(A[10]), .ZN(n176) );
  NAND2_X1 U82 ( .A1(b[2]), .A2(n71), .ZN(n51) );
  NAND2_X1 U83 ( .A1(b[1]), .A2(b[0]), .ZN(n71) );
  NAND2_X1 U84 ( .A1(n68), .A2(n72), .ZN(n66) );
  OAI21_X1 U85 ( .B1(A[9]), .B2(n177), .A(A[10]), .ZN(n72) );
  INV_X1 U86 ( .A(n31), .ZN(n177) );
  INV_X1 U87 ( .A(A[9]), .ZN(n165) );
  INV_X1 U88 ( .A(A[12]), .ZN(n166) );
  INV_X1 U89 ( .A(A[13]), .ZN(n167) );
endmodule


module BOOTH_ENCODER_WIDTH16_7 ( A, b, vp );
  input [15:0] A;
  input [2:0] b;
  output [16:0] vp;
  wire   \notA[0] , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236;
  assign \notA[0]  = A[0];

  XOR2_X1 U90 ( .A(n31), .B(A[9]), .Z(n21) );
  NAND3_X1 U91 ( .A1(n223), .A2(n217), .A3(n31), .ZN(n68) );
  NOR2_X2 U3 ( .A1(n71), .A2(b[2]), .ZN(n26) );
  NOR2_X2 U4 ( .A1(n70), .A2(b[2]), .ZN(n29) );
  OR2_X1 U5 ( .A1(n70), .A2(n51), .ZN(n22) );
  INV_X1 U6 ( .A(n62), .ZN(n220) );
  INV_X1 U7 ( .A(n24), .ZN(n234) );
  OAI21_X1 U8 ( .B1(n64), .B2(n218), .A(n62), .ZN(n60) );
  OAI21_X1 U9 ( .B1(n220), .B2(n219), .A(n57), .ZN(n58) );
  NAND2_X1 U10 ( .A1(n220), .A2(n219), .ZN(n57) );
  INV_X1 U11 ( .A(n49), .ZN(n229) );
  INV_X1 U12 ( .A(n40), .ZN(n227) );
  NAND2_X1 U13 ( .A1(n64), .A2(n218), .ZN(n62) );
  OAI221_X1 U14 ( .B1(n22), .B2(n41), .C1(n234), .C2(n230), .A(n44), .ZN(vp[3]) );
  AOI22_X1 U15 ( .A1(A[2]), .A2(n26), .B1(A[3]), .B2(n29), .ZN(n44) );
  OAI221_X1 U16 ( .B1(n22), .B2(n36), .C1(n234), .C2(n41), .A(n42), .ZN(vp[4])
         );
  AOI22_X1 U17 ( .A1(A[3]), .A2(n26), .B1(A[4]), .B2(n29), .ZN(n42) );
  OAI221_X1 U18 ( .B1(n22), .B2(n228), .C1(n234), .C2(n36), .A(n37), .ZN(vp[5]) );
  AOI22_X1 U19 ( .A1(A[4]), .A2(n26), .B1(A[5]), .B2(n29), .ZN(n37) );
  OAI221_X1 U20 ( .B1(n22), .B2(n32), .C1(n234), .C2(n228), .A(n35), .ZN(vp[6]) );
  AOI22_X1 U21 ( .A1(A[5]), .A2(n26), .B1(A[6]), .B2(n29), .ZN(n35) );
  OAI221_X1 U22 ( .B1(n22), .B2(n27), .C1(n234), .C2(n32), .A(n33), .ZN(vp[7])
         );
  AOI22_X1 U23 ( .A1(A[6]), .A2(n26), .B1(A[7]), .B2(n29), .ZN(n33) );
  OAI221_X1 U24 ( .B1(n22), .B2(n66), .C1(n233), .C2(n223), .A(n224), .ZN(
        vp[10]) );
  INV_X1 U25 ( .A(n69), .ZN(n224) );
  OAI22_X1 U26 ( .A1(n217), .A2(n235), .B1(n21), .B2(n234), .ZN(n69) );
  OAI221_X1 U27 ( .B1(n22), .B2(n221), .C1(n235), .C2(n223), .A(n65), .ZN(
        vp[11]) );
  AOI22_X1 U28 ( .A1(n222), .A2(n24), .B1(A[11]), .B2(n29), .ZN(n65) );
  INV_X1 U29 ( .A(n66), .ZN(n222) );
  OAI221_X1 U30 ( .B1(n22), .B2(n60), .C1(n234), .C2(n221), .A(n63), .ZN(
        vp[12]) );
  AOI22_X1 U31 ( .A1(A[11]), .A2(n26), .B1(A[12]), .B2(n29), .ZN(n63) );
  OAI221_X1 U32 ( .B1(n22), .B2(n58), .C1(n234), .C2(n60), .A(n61), .ZN(vp[13]) );
  AOI22_X1 U33 ( .A1(A[12]), .A2(n26), .B1(A[13]), .B2(n29), .ZN(n61) );
  OAI221_X1 U34 ( .B1(n22), .B2(n54), .C1(n234), .C2(n58), .A(n59), .ZN(vp[14]) );
  AOI22_X1 U35 ( .A1(A[13]), .A2(n26), .B1(A[14]), .B2(n29), .ZN(n59) );
  OAI221_X1 U36 ( .B1(n22), .B2(n52), .C1(n234), .C2(n54), .A(n55), .ZN(vp[15]) );
  AOI22_X1 U37 ( .A1(A[14]), .A2(n26), .B1(A[15]), .B2(n29), .ZN(n55) );
  OAI221_X1 U38 ( .B1(n21), .B2(n22), .C1(n217), .C2(n233), .A(n23), .ZN(vp[9]) );
  AOI22_X1 U39 ( .A1(n24), .A2(n25), .B1(n26), .B2(A[8]), .ZN(n23) );
  OAI221_X1 U40 ( .B1(n226), .B2(n22), .C1(n234), .C2(n27), .A(n28), .ZN(vp[8]) );
  INV_X1 U41 ( .A(n25), .ZN(n226) );
  AOI22_X1 U42 ( .A1(A[7]), .A2(n26), .B1(n29), .B2(A[8]), .ZN(n28) );
  NOR2_X1 U43 ( .A1(n51), .A2(n236), .ZN(n24) );
  INV_X1 U44 ( .A(n70), .ZN(n236) );
  NOR2_X1 U45 ( .A1(n30), .A2(A[8]), .ZN(n31) );
  AOI21_X1 U46 ( .B1(n30), .B2(A[8]), .A(n31), .ZN(n25) );
  NOR2_X1 U47 ( .A1(n68), .A2(A[11]), .ZN(n64) );
  XNOR2_X1 U48 ( .A(n229), .B(A[3]), .ZN(n41) );
  XNOR2_X1 U49 ( .A(n227), .B(A[6]), .ZN(n32) );
  XOR2_X1 U50 ( .A(n216), .B(A[15]), .Z(n52) );
  NOR2_X1 U51 ( .A1(n57), .A2(A[14]), .ZN(n216) );
  XNOR2_X1 U52 ( .A(n57), .B(A[14]), .ZN(n54) );
  NOR2_X1 U53 ( .A1(n48), .A2(A[2]), .ZN(n49) );
  NOR2_X1 U54 ( .A1(n39), .A2(A[5]), .ZN(n40) );
  AOI21_X1 U55 ( .B1(n233), .B2(n22), .A(n232), .ZN(vp[0]) );
  OAI21_X1 U56 ( .B1(n231), .B2(n232), .A(n48), .ZN(n45) );
  OAI21_X1 U57 ( .B1(n51), .B2(n52), .A(n53), .ZN(vp[16]) );
  OAI21_X1 U58 ( .B1(n26), .B2(n29), .A(A[15]), .ZN(n53) );
  INV_X1 U59 ( .A(n29), .ZN(n233) );
  NAND2_X1 U60 ( .A1(n231), .A2(n232), .ZN(n48) );
  INV_X1 U61 ( .A(n26), .ZN(n235) );
  NAND2_X1 U62 ( .A1(n39), .A2(n43), .ZN(n36) );
  OAI21_X1 U63 ( .B1(A[3]), .B2(n229), .A(A[4]), .ZN(n43) );
  NAND2_X1 U64 ( .A1(n30), .A2(n34), .ZN(n27) );
  OAI21_X1 U65 ( .B1(A[6]), .B2(n227), .A(A[7]), .ZN(n34) );
  OR3_X1 U66 ( .A1(A[3]), .A2(A[4]), .A3(n229), .ZN(n39) );
  OR3_X1 U67 ( .A1(A[6]), .A2(A[7]), .A3(n227), .ZN(n30) );
  INV_X1 U68 ( .A(n47), .ZN(n230) );
  AOI21_X1 U69 ( .B1(n48), .B2(A[2]), .A(n49), .ZN(n47) );
  INV_X1 U70 ( .A(n38), .ZN(n228) );
  AOI21_X1 U71 ( .B1(n39), .B2(A[5]), .A(n40), .ZN(n38) );
  INV_X1 U72 ( .A(n67), .ZN(n221) );
  AOI21_X1 U73 ( .B1(n68), .B2(A[11]), .A(n64), .ZN(n67) );
  OAI21_X1 U74 ( .B1(b[1]), .B2(b[0]), .A(n71), .ZN(n70) );
  OAI221_X1 U75 ( .B1(n22), .B2(n45), .C1(n233), .C2(n231), .A(n50), .ZN(vp[1]) );
  OAI21_X1 U76 ( .B1(n26), .B2(n24), .A(\notA[0] ), .ZN(n50) );
  OAI221_X1 U77 ( .B1(n22), .B2(n230), .C1(n234), .C2(n45), .A(n46), .ZN(vp[2]) );
  AOI22_X1 U78 ( .A1(A[1]), .A2(n26), .B1(A[2]), .B2(n29), .ZN(n46) );
  INV_X1 U79 ( .A(\notA[0] ), .ZN(n232) );
  INV_X1 U80 ( .A(A[1]), .ZN(n231) );
  INV_X1 U81 ( .A(A[10]), .ZN(n223) );
  NAND2_X1 U82 ( .A1(b[1]), .A2(b[0]), .ZN(n71) );
  NAND2_X1 U83 ( .A1(b[2]), .A2(n71), .ZN(n51) );
  NAND2_X1 U84 ( .A1(n68), .A2(n72), .ZN(n66) );
  OAI21_X1 U85 ( .B1(A[9]), .B2(n225), .A(A[10]), .ZN(n72) );
  INV_X1 U86 ( .A(n31), .ZN(n225) );
  INV_X1 U87 ( .A(A[9]), .ZN(n217) );
  INV_X1 U88 ( .A(A[12]), .ZN(n218) );
  INV_X1 U89 ( .A(A[13]), .ZN(n219) );
endmodule


module BOOTH_ENCODER_WIDTH16_6 ( A, b, vp );
  input [15:0] A;
  input [2:0] b;
  output [16:0] vp;
  wire   \notA[0] , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336;
  assign \notA[0]  = A[0];

  XOR2_X1 U90 ( .A(n31), .B(A[9]), .Z(n21) );
  NAND3_X1 U91 ( .A1(n323), .A2(n317), .A3(n31), .ZN(n68) );
  NOR2_X2 U3 ( .A1(n71), .A2(b[2]), .ZN(n26) );
  NOR2_X2 U4 ( .A1(n70), .A2(b[2]), .ZN(n29) );
  OR2_X1 U5 ( .A1(n70), .A2(n51), .ZN(n22) );
  INV_X1 U6 ( .A(n62), .ZN(n320) );
  INV_X1 U7 ( .A(n24), .ZN(n334) );
  OAI21_X1 U8 ( .B1(n64), .B2(n318), .A(n62), .ZN(n60) );
  OAI21_X1 U9 ( .B1(n320), .B2(n319), .A(n57), .ZN(n58) );
  INV_X1 U10 ( .A(n49), .ZN(n329) );
  INV_X1 U11 ( .A(n40), .ZN(n327) );
  NAND2_X1 U12 ( .A1(n320), .A2(n319), .ZN(n57) );
  NAND2_X1 U13 ( .A1(n64), .A2(n318), .ZN(n62) );
  AOI21_X1 U14 ( .B1(n30), .B2(A[8]), .A(n31), .ZN(n25) );
  NOR2_X1 U15 ( .A1(n30), .A2(A[8]), .ZN(n31) );
  OAI221_X1 U16 ( .B1(n22), .B2(n54), .C1(n334), .C2(n58), .A(n59), .ZN(vp[14]) );
  AOI22_X1 U17 ( .A1(A[13]), .A2(n26), .B1(A[14]), .B2(n29), .ZN(n59) );
  OAI221_X1 U18 ( .B1(n22), .B2(n41), .C1(n334), .C2(n330), .A(n44), .ZN(vp[3]) );
  AOI22_X1 U19 ( .A1(A[2]), .A2(n26), .B1(A[3]), .B2(n29), .ZN(n44) );
  OAI221_X1 U20 ( .B1(n22), .B2(n36), .C1(n334), .C2(n41), .A(n42), .ZN(vp[4])
         );
  AOI22_X1 U21 ( .A1(A[3]), .A2(n26), .B1(A[4]), .B2(n29), .ZN(n42) );
  OAI221_X1 U22 ( .B1(n22), .B2(n328), .C1(n334), .C2(n36), .A(n37), .ZN(vp[5]) );
  AOI22_X1 U23 ( .A1(A[4]), .A2(n26), .B1(A[5]), .B2(n29), .ZN(n37) );
  OAI221_X1 U24 ( .B1(n22), .B2(n32), .C1(n334), .C2(n328), .A(n35), .ZN(vp[6]) );
  AOI22_X1 U25 ( .A1(A[5]), .A2(n26), .B1(A[6]), .B2(n29), .ZN(n35) );
  OAI221_X1 U26 ( .B1(n22), .B2(n27), .C1(n334), .C2(n32), .A(n33), .ZN(vp[7])
         );
  AOI22_X1 U27 ( .A1(A[6]), .A2(n26), .B1(A[7]), .B2(n29), .ZN(n33) );
  OAI221_X1 U28 ( .B1(n22), .B2(n66), .C1(n333), .C2(n323), .A(n324), .ZN(
        vp[10]) );
  INV_X1 U29 ( .A(n69), .ZN(n324) );
  OAI22_X1 U30 ( .A1(n317), .A2(n335), .B1(n21), .B2(n334), .ZN(n69) );
  OAI221_X1 U31 ( .B1(n22), .B2(n321), .C1(n335), .C2(n323), .A(n65), .ZN(
        vp[11]) );
  AOI22_X1 U32 ( .A1(n322), .A2(n24), .B1(A[11]), .B2(n29), .ZN(n65) );
  INV_X1 U33 ( .A(n66), .ZN(n322) );
  OAI221_X1 U34 ( .B1(n22), .B2(n60), .C1(n334), .C2(n321), .A(n63), .ZN(
        vp[12]) );
  AOI22_X1 U35 ( .A1(A[11]), .A2(n26), .B1(A[12]), .B2(n29), .ZN(n63) );
  OAI221_X1 U36 ( .B1(n22), .B2(n58), .C1(n334), .C2(n60), .A(n61), .ZN(vp[13]) );
  AOI22_X1 U37 ( .A1(A[12]), .A2(n26), .B1(A[13]), .B2(n29), .ZN(n61) );
  OAI221_X1 U38 ( .B1(n22), .B2(n52), .C1(n334), .C2(n54), .A(n55), .ZN(vp[15]) );
  AOI22_X1 U39 ( .A1(A[14]), .A2(n26), .B1(A[15]), .B2(n29), .ZN(n55) );
  OAI221_X1 U40 ( .B1(n21), .B2(n22), .C1(n317), .C2(n333), .A(n23), .ZN(vp[9]) );
  AOI22_X1 U41 ( .A1(n24), .A2(n25), .B1(n26), .B2(A[8]), .ZN(n23) );
  OAI221_X1 U42 ( .B1(n326), .B2(n22), .C1(n334), .C2(n27), .A(n28), .ZN(vp[8]) );
  INV_X1 U43 ( .A(n25), .ZN(n326) );
  AOI22_X1 U44 ( .A1(A[7]), .A2(n26), .B1(n29), .B2(A[8]), .ZN(n28) );
  NOR2_X1 U45 ( .A1(n51), .A2(n336), .ZN(n24) );
  INV_X1 U46 ( .A(n70), .ZN(n336) );
  NOR2_X1 U47 ( .A1(n68), .A2(A[11]), .ZN(n64) );
  XNOR2_X1 U48 ( .A(n57), .B(A[14]), .ZN(n54) );
  XNOR2_X1 U49 ( .A(n329), .B(A[3]), .ZN(n41) );
  XNOR2_X1 U50 ( .A(n327), .B(A[6]), .ZN(n32) );
  NOR2_X1 U51 ( .A1(n48), .A2(A[2]), .ZN(n49) );
  NOR2_X1 U52 ( .A1(n39), .A2(A[5]), .ZN(n40) );
  XOR2_X1 U53 ( .A(n316), .B(A[15]), .Z(n52) );
  NOR2_X1 U54 ( .A1(n57), .A2(A[14]), .ZN(n316) );
  AOI21_X1 U55 ( .B1(n333), .B2(n22), .A(n332), .ZN(vp[0]) );
  OAI21_X1 U56 ( .B1(n331), .B2(n332), .A(n48), .ZN(n45) );
  OAI21_X1 U57 ( .B1(n51), .B2(n52), .A(n53), .ZN(vp[16]) );
  OAI21_X1 U58 ( .B1(n26), .B2(n29), .A(A[15]), .ZN(n53) );
  INV_X1 U59 ( .A(n29), .ZN(n333) );
  NAND2_X1 U60 ( .A1(n331), .A2(n332), .ZN(n48) );
  INV_X1 U61 ( .A(n26), .ZN(n335) );
  NAND2_X1 U62 ( .A1(n39), .A2(n43), .ZN(n36) );
  OAI21_X1 U63 ( .B1(A[3]), .B2(n329), .A(A[4]), .ZN(n43) );
  NAND2_X1 U64 ( .A1(n30), .A2(n34), .ZN(n27) );
  OAI21_X1 U65 ( .B1(A[6]), .B2(n327), .A(A[7]), .ZN(n34) );
  OR3_X1 U66 ( .A1(A[3]), .A2(A[4]), .A3(n329), .ZN(n39) );
  OR3_X1 U67 ( .A1(A[6]), .A2(A[7]), .A3(n327), .ZN(n30) );
  INV_X1 U68 ( .A(n47), .ZN(n330) );
  AOI21_X1 U69 ( .B1(n48), .B2(A[2]), .A(n49), .ZN(n47) );
  INV_X1 U70 ( .A(n38), .ZN(n328) );
  AOI21_X1 U71 ( .B1(n39), .B2(A[5]), .A(n40), .ZN(n38) );
  INV_X1 U72 ( .A(n67), .ZN(n321) );
  AOI21_X1 U73 ( .B1(n68), .B2(A[11]), .A(n64), .ZN(n67) );
  OAI21_X1 U74 ( .B1(b[1]), .B2(b[0]), .A(n71), .ZN(n70) );
  OAI221_X1 U75 ( .B1(n22), .B2(n45), .C1(n333), .C2(n331), .A(n50), .ZN(vp[1]) );
  OAI21_X1 U76 ( .B1(n26), .B2(n24), .A(\notA[0] ), .ZN(n50) );
  OAI221_X1 U77 ( .B1(n22), .B2(n330), .C1(n334), .C2(n45), .A(n46), .ZN(vp[2]) );
  AOI22_X1 U78 ( .A1(A[1]), .A2(n26), .B1(A[2]), .B2(n29), .ZN(n46) );
  INV_X1 U79 ( .A(\notA[0] ), .ZN(n332) );
  INV_X1 U80 ( .A(A[1]), .ZN(n331) );
  INV_X1 U81 ( .A(A[10]), .ZN(n323) );
  NAND2_X1 U82 ( .A1(b[1]), .A2(b[0]), .ZN(n71) );
  NAND2_X1 U83 ( .A1(b[2]), .A2(n71), .ZN(n51) );
  NAND2_X1 U84 ( .A1(n68), .A2(n72), .ZN(n66) );
  OAI21_X1 U85 ( .B1(A[9]), .B2(n325), .A(A[10]), .ZN(n72) );
  INV_X1 U86 ( .A(n31), .ZN(n325) );
  INV_X1 U87 ( .A(A[9]), .ZN(n317) );
  INV_X1 U88 ( .A(A[12]), .ZN(n318) );
  INV_X1 U89 ( .A(A[13]), .ZN(n319) );
endmodule


module BOOTH_ENCODER_WIDTH16_5 ( A, b, vp );
  input [15:0] A;
  input [2:0] b;
  output [16:0] vp;
  wire   \notA[0] , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337;
  assign \notA[0]  = A[0];

  XOR2_X1 U90 ( .A(n31), .B(A[9]), .Z(n21) );
  NAND3_X1 U91 ( .A1(n324), .A2(n318), .A3(n31), .ZN(n68) );
  NOR2_X2 U3 ( .A1(n71), .A2(b[2]), .ZN(n26) );
  NOR2_X2 U4 ( .A1(n70), .A2(b[2]), .ZN(n29) );
  OR2_X1 U5 ( .A1(n70), .A2(n51), .ZN(n22) );
  INV_X1 U6 ( .A(n62), .ZN(n321) );
  INV_X1 U7 ( .A(n24), .ZN(n335) );
  OAI21_X1 U8 ( .B1(n64), .B2(n319), .A(n62), .ZN(n60) );
  OAI21_X1 U9 ( .B1(n321), .B2(n320), .A(n57), .ZN(n58) );
  INV_X1 U10 ( .A(n49), .ZN(n330) );
  INV_X1 U11 ( .A(n40), .ZN(n328) );
  NAND2_X1 U12 ( .A1(n321), .A2(n320), .ZN(n57) );
  NAND2_X1 U13 ( .A1(n64), .A2(n319), .ZN(n62) );
  AOI21_X1 U14 ( .B1(n30), .B2(A[8]), .A(n31), .ZN(n25) );
  NOR2_X1 U15 ( .A1(n30), .A2(A[8]), .ZN(n31) );
  OAI221_X1 U16 ( .B1(n22), .B2(n54), .C1(n335), .C2(n58), .A(n59), .ZN(vp[14]) );
  AOI22_X1 U17 ( .A1(A[13]), .A2(n26), .B1(A[14]), .B2(n29), .ZN(n59) );
  OAI221_X1 U18 ( .B1(n22), .B2(n41), .C1(n335), .C2(n331), .A(n44), .ZN(vp[3]) );
  AOI22_X1 U19 ( .A1(A[2]), .A2(n26), .B1(A[3]), .B2(n29), .ZN(n44) );
  OAI221_X1 U20 ( .B1(n22), .B2(n36), .C1(n335), .C2(n41), .A(n42), .ZN(vp[4])
         );
  AOI22_X1 U21 ( .A1(A[3]), .A2(n26), .B1(A[4]), .B2(n29), .ZN(n42) );
  OAI221_X1 U22 ( .B1(n22), .B2(n329), .C1(n335), .C2(n36), .A(n37), .ZN(vp[5]) );
  AOI22_X1 U23 ( .A1(A[4]), .A2(n26), .B1(A[5]), .B2(n29), .ZN(n37) );
  OAI221_X1 U24 ( .B1(n22), .B2(n32), .C1(n335), .C2(n329), .A(n35), .ZN(vp[6]) );
  AOI22_X1 U25 ( .A1(A[5]), .A2(n26), .B1(A[6]), .B2(n29), .ZN(n35) );
  OAI221_X1 U26 ( .B1(n22), .B2(n27), .C1(n335), .C2(n32), .A(n33), .ZN(vp[7])
         );
  AOI22_X1 U27 ( .A1(A[6]), .A2(n26), .B1(A[7]), .B2(n29), .ZN(n33) );
  OAI221_X1 U28 ( .B1(n22), .B2(n66), .C1(n334), .C2(n324), .A(n325), .ZN(
        vp[10]) );
  INV_X1 U29 ( .A(n69), .ZN(n325) );
  OAI22_X1 U30 ( .A1(n318), .A2(n336), .B1(n21), .B2(n335), .ZN(n69) );
  OAI221_X1 U31 ( .B1(n22), .B2(n322), .C1(n336), .C2(n324), .A(n65), .ZN(
        vp[11]) );
  AOI22_X1 U32 ( .A1(n323), .A2(n24), .B1(A[11]), .B2(n29), .ZN(n65) );
  INV_X1 U33 ( .A(n66), .ZN(n323) );
  OAI221_X1 U34 ( .B1(n22), .B2(n60), .C1(n335), .C2(n322), .A(n63), .ZN(
        vp[12]) );
  AOI22_X1 U35 ( .A1(A[11]), .A2(n26), .B1(A[12]), .B2(n29), .ZN(n63) );
  OAI221_X1 U36 ( .B1(n22), .B2(n58), .C1(n335), .C2(n60), .A(n61), .ZN(vp[13]) );
  AOI22_X1 U37 ( .A1(A[12]), .A2(n26), .B1(A[13]), .B2(n29), .ZN(n61) );
  OAI221_X1 U38 ( .B1(n22), .B2(n52), .C1(n335), .C2(n54), .A(n55), .ZN(vp[15]) );
  AOI22_X1 U39 ( .A1(A[14]), .A2(n26), .B1(A[15]), .B2(n29), .ZN(n55) );
  OAI221_X1 U40 ( .B1(n21), .B2(n22), .C1(n318), .C2(n334), .A(n23), .ZN(vp[9]) );
  AOI22_X1 U41 ( .A1(n24), .A2(n25), .B1(n26), .B2(A[8]), .ZN(n23) );
  OAI221_X1 U42 ( .B1(n327), .B2(n22), .C1(n335), .C2(n27), .A(n28), .ZN(vp[8]) );
  INV_X1 U43 ( .A(n25), .ZN(n327) );
  AOI22_X1 U44 ( .A1(A[7]), .A2(n26), .B1(n29), .B2(A[8]), .ZN(n28) );
  NOR2_X1 U45 ( .A1(n51), .A2(n337), .ZN(n24) );
  INV_X1 U46 ( .A(n70), .ZN(n337) );
  NOR2_X1 U47 ( .A1(n68), .A2(A[11]), .ZN(n64) );
  XNOR2_X1 U48 ( .A(n57), .B(A[14]), .ZN(n54) );
  XNOR2_X1 U49 ( .A(n330), .B(A[3]), .ZN(n41) );
  XNOR2_X1 U50 ( .A(n328), .B(A[6]), .ZN(n32) );
  NOR2_X1 U51 ( .A1(n48), .A2(A[2]), .ZN(n49) );
  NOR2_X1 U52 ( .A1(n39), .A2(A[5]), .ZN(n40) );
  XOR2_X1 U53 ( .A(n317), .B(A[15]), .Z(n52) );
  NOR2_X1 U54 ( .A1(n57), .A2(A[14]), .ZN(n317) );
  AOI21_X1 U55 ( .B1(n334), .B2(n22), .A(n333), .ZN(vp[0]) );
  OAI21_X1 U56 ( .B1(n332), .B2(n333), .A(n48), .ZN(n45) );
  OAI21_X1 U57 ( .B1(n51), .B2(n52), .A(n53), .ZN(vp[16]) );
  OAI21_X1 U58 ( .B1(n26), .B2(n29), .A(A[15]), .ZN(n53) );
  INV_X1 U59 ( .A(n29), .ZN(n334) );
  NAND2_X1 U60 ( .A1(n332), .A2(n333), .ZN(n48) );
  INV_X1 U61 ( .A(n26), .ZN(n336) );
  NAND2_X1 U62 ( .A1(n39), .A2(n43), .ZN(n36) );
  OAI21_X1 U63 ( .B1(A[3]), .B2(n330), .A(A[4]), .ZN(n43) );
  NAND2_X1 U64 ( .A1(n30), .A2(n34), .ZN(n27) );
  OAI21_X1 U65 ( .B1(A[6]), .B2(n328), .A(A[7]), .ZN(n34) );
  OR3_X1 U66 ( .A1(A[3]), .A2(A[4]), .A3(n330), .ZN(n39) );
  OR3_X1 U67 ( .A1(A[6]), .A2(A[7]), .A3(n328), .ZN(n30) );
  INV_X1 U68 ( .A(n47), .ZN(n331) );
  AOI21_X1 U69 ( .B1(n48), .B2(A[2]), .A(n49), .ZN(n47) );
  INV_X1 U70 ( .A(n38), .ZN(n329) );
  AOI21_X1 U71 ( .B1(n39), .B2(A[5]), .A(n40), .ZN(n38) );
  INV_X1 U72 ( .A(n67), .ZN(n322) );
  AOI21_X1 U73 ( .B1(n68), .B2(A[11]), .A(n64), .ZN(n67) );
  OAI21_X1 U74 ( .B1(b[1]), .B2(b[0]), .A(n71), .ZN(n70) );
  OAI221_X1 U75 ( .B1(n22), .B2(n45), .C1(n334), .C2(n332), .A(n50), .ZN(vp[1]) );
  OAI21_X1 U76 ( .B1(n26), .B2(n24), .A(\notA[0] ), .ZN(n50) );
  OAI221_X1 U77 ( .B1(n22), .B2(n331), .C1(n335), .C2(n45), .A(n46), .ZN(vp[2]) );
  AOI22_X1 U78 ( .A1(A[1]), .A2(n26), .B1(A[2]), .B2(n29), .ZN(n46) );
  INV_X1 U79 ( .A(\notA[0] ), .ZN(n333) );
  INV_X1 U80 ( .A(A[1]), .ZN(n332) );
  INV_X1 U81 ( .A(A[10]), .ZN(n324) );
  NAND2_X1 U82 ( .A1(b[1]), .A2(b[0]), .ZN(n71) );
  NAND2_X1 U83 ( .A1(b[2]), .A2(n71), .ZN(n51) );
  NAND2_X1 U84 ( .A1(n68), .A2(n72), .ZN(n66) );
  OAI21_X1 U85 ( .B1(A[9]), .B2(n326), .A(A[10]), .ZN(n72) );
  INV_X1 U86 ( .A(n31), .ZN(n326) );
  INV_X1 U87 ( .A(A[9]), .ZN(n318) );
  INV_X1 U88 ( .A(A[12]), .ZN(n319) );
  INV_X1 U89 ( .A(A[13]), .ZN(n320) );
endmodule


module BOOTH_ENCODER_WIDTH16_4 ( A, b, vp );
  input [15:0] A;
  input [2:0] b;
  output [16:0] vp;
  wire   \notA[0] , n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388;
  assign \notA[0]  = A[0];

  XOR2_X1 U90 ( .A(n378), .B(A[9]), .Z(n388) );
  NAND3_X1 U91 ( .A1(n324), .A2(n318), .A3(n378), .ZN(n342) );
  NOR2_X2 U3 ( .A1(n339), .A2(b[2]), .ZN(n383) );
  NOR2_X2 U4 ( .A1(n340), .A2(b[2]), .ZN(n380) );
  OR2_X1 U5 ( .A1(n340), .A2(n358), .ZN(n387) );
  INV_X1 U6 ( .A(n348), .ZN(n321) );
  INV_X1 U7 ( .A(n385), .ZN(n335) );
  OAI21_X1 U8 ( .B1(n346), .B2(n319), .A(n348), .ZN(n350) );
  OAI21_X1 U9 ( .B1(n321), .B2(n320), .A(n353), .ZN(n352) );
  INV_X1 U10 ( .A(n360), .ZN(n330) );
  INV_X1 U11 ( .A(n369), .ZN(n328) );
  NAND2_X1 U12 ( .A1(n321), .A2(n320), .ZN(n353) );
  NAND2_X1 U13 ( .A1(n346), .A2(n319), .ZN(n348) );
  AOI21_X1 U14 ( .B1(n379), .B2(A[8]), .A(n378), .ZN(n384) );
  NOR2_X1 U15 ( .A1(n379), .A2(A[8]), .ZN(n378) );
  OAI221_X1 U16 ( .B1(n387), .B2(n355), .C1(n335), .C2(n352), .A(n351), .ZN(
        vp[14]) );
  AOI22_X1 U17 ( .A1(A[13]), .A2(n383), .B1(A[14]), .B2(n380), .ZN(n351) );
  OAI221_X1 U18 ( .B1(n387), .B2(n368), .C1(n335), .C2(n331), .A(n365), .ZN(
        vp[3]) );
  AOI22_X1 U19 ( .A1(A[2]), .A2(n383), .B1(A[3]), .B2(n380), .ZN(n365) );
  OAI221_X1 U20 ( .B1(n387), .B2(n373), .C1(n335), .C2(n368), .A(n367), .ZN(
        vp[4]) );
  AOI22_X1 U21 ( .A1(A[3]), .A2(n383), .B1(A[4]), .B2(n380), .ZN(n367) );
  OAI221_X1 U22 ( .B1(n387), .B2(n329), .C1(n335), .C2(n373), .A(n372), .ZN(
        vp[5]) );
  AOI22_X1 U23 ( .A1(A[4]), .A2(n383), .B1(A[5]), .B2(n380), .ZN(n372) );
  OAI221_X1 U24 ( .B1(n387), .B2(n377), .C1(n335), .C2(n329), .A(n374), .ZN(
        vp[6]) );
  AOI22_X1 U25 ( .A1(A[5]), .A2(n383), .B1(A[6]), .B2(n380), .ZN(n374) );
  OAI221_X1 U26 ( .B1(n387), .B2(n382), .C1(n335), .C2(n377), .A(n376), .ZN(
        vp[7]) );
  AOI22_X1 U27 ( .A1(A[6]), .A2(n383), .B1(A[7]), .B2(n380), .ZN(n376) );
  OAI221_X1 U28 ( .B1(n387), .B2(n344), .C1(n334), .C2(n324), .A(n325), .ZN(
        vp[10]) );
  INV_X1 U29 ( .A(n341), .ZN(n325) );
  OAI22_X1 U30 ( .A1(n318), .A2(n336), .B1(n388), .B2(n335), .ZN(n341) );
  OAI221_X1 U31 ( .B1(n387), .B2(n322), .C1(n336), .C2(n324), .A(n345), .ZN(
        vp[11]) );
  AOI22_X1 U32 ( .A1(n323), .A2(n385), .B1(A[11]), .B2(n380), .ZN(n345) );
  INV_X1 U33 ( .A(n344), .ZN(n323) );
  OAI221_X1 U34 ( .B1(n387), .B2(n350), .C1(n335), .C2(n322), .A(n347), .ZN(
        vp[12]) );
  AOI22_X1 U35 ( .A1(A[11]), .A2(n383), .B1(A[12]), .B2(n380), .ZN(n347) );
  OAI221_X1 U36 ( .B1(n387), .B2(n352), .C1(n335), .C2(n350), .A(n349), .ZN(
        vp[13]) );
  AOI22_X1 U37 ( .A1(A[12]), .A2(n383), .B1(A[13]), .B2(n380), .ZN(n349) );
  OAI221_X1 U38 ( .B1(n387), .B2(n357), .C1(n335), .C2(n355), .A(n354), .ZN(
        vp[15]) );
  AOI22_X1 U39 ( .A1(A[14]), .A2(n383), .B1(A[15]), .B2(n380), .ZN(n354) );
  OAI221_X1 U40 ( .B1(n388), .B2(n387), .C1(n318), .C2(n334), .A(n386), .ZN(
        vp[9]) );
  AOI22_X1 U41 ( .A1(n385), .A2(n384), .B1(n383), .B2(A[8]), .ZN(n386) );
  OAI221_X1 U42 ( .B1(n327), .B2(n387), .C1(n335), .C2(n382), .A(n381), .ZN(
        vp[8]) );
  INV_X1 U43 ( .A(n384), .ZN(n327) );
  AOI22_X1 U44 ( .A1(A[7]), .A2(n383), .B1(n380), .B2(A[8]), .ZN(n381) );
  NOR2_X1 U45 ( .A1(n358), .A2(n337), .ZN(n385) );
  INV_X1 U46 ( .A(n340), .ZN(n337) );
  NOR2_X1 U47 ( .A1(n342), .A2(A[11]), .ZN(n346) );
  XNOR2_X1 U48 ( .A(n353), .B(A[14]), .ZN(n355) );
  XNOR2_X1 U49 ( .A(n330), .B(A[3]), .ZN(n368) );
  XNOR2_X1 U50 ( .A(n328), .B(A[6]), .ZN(n377) );
  NOR2_X1 U51 ( .A1(n361), .A2(A[2]), .ZN(n360) );
  NOR2_X1 U52 ( .A1(n370), .A2(A[5]), .ZN(n369) );
  XOR2_X1 U53 ( .A(n317), .B(A[15]), .Z(n357) );
  NOR2_X1 U54 ( .A1(n353), .A2(A[14]), .ZN(n317) );
  AOI21_X1 U55 ( .B1(n334), .B2(n387), .A(n333), .ZN(vp[0]) );
  OAI21_X1 U56 ( .B1(n332), .B2(n333), .A(n361), .ZN(n364) );
  OAI21_X1 U57 ( .B1(n358), .B2(n357), .A(n356), .ZN(vp[16]) );
  OAI21_X1 U58 ( .B1(n383), .B2(n380), .A(A[15]), .ZN(n356) );
  INV_X1 U59 ( .A(n380), .ZN(n334) );
  NAND2_X1 U60 ( .A1(n332), .A2(n333), .ZN(n361) );
  INV_X1 U61 ( .A(n383), .ZN(n336) );
  NAND2_X1 U62 ( .A1(n370), .A2(n366), .ZN(n373) );
  OAI21_X1 U63 ( .B1(A[3]), .B2(n330), .A(A[4]), .ZN(n366) );
  NAND2_X1 U64 ( .A1(n379), .A2(n375), .ZN(n382) );
  OAI21_X1 U65 ( .B1(A[6]), .B2(n328), .A(A[7]), .ZN(n375) );
  OR3_X1 U66 ( .A1(A[3]), .A2(A[4]), .A3(n330), .ZN(n370) );
  OR3_X1 U67 ( .A1(A[6]), .A2(A[7]), .A3(n328), .ZN(n379) );
  INV_X1 U68 ( .A(n362), .ZN(n331) );
  AOI21_X1 U69 ( .B1(n361), .B2(A[2]), .A(n360), .ZN(n362) );
  INV_X1 U70 ( .A(n371), .ZN(n329) );
  AOI21_X1 U71 ( .B1(n370), .B2(A[5]), .A(n369), .ZN(n371) );
  INV_X1 U72 ( .A(n343), .ZN(n322) );
  AOI21_X1 U73 ( .B1(n342), .B2(A[11]), .A(n346), .ZN(n343) );
  OAI21_X1 U74 ( .B1(b[1]), .B2(b[0]), .A(n339), .ZN(n340) );
  OAI221_X1 U75 ( .B1(n387), .B2(n364), .C1(n334), .C2(n332), .A(n359), .ZN(
        vp[1]) );
  OAI21_X1 U76 ( .B1(n383), .B2(n385), .A(\notA[0] ), .ZN(n359) );
  OAI221_X1 U77 ( .B1(n387), .B2(n331), .C1(n335), .C2(n364), .A(n363), .ZN(
        vp[2]) );
  AOI22_X1 U78 ( .A1(A[1]), .A2(n383), .B1(A[2]), .B2(n380), .ZN(n363) );
  INV_X1 U79 ( .A(\notA[0] ), .ZN(n333) );
  INV_X1 U80 ( .A(A[1]), .ZN(n332) );
  INV_X1 U81 ( .A(A[10]), .ZN(n324) );
  NAND2_X1 U82 ( .A1(b[1]), .A2(b[0]), .ZN(n339) );
  NAND2_X1 U83 ( .A1(b[2]), .A2(n339), .ZN(n358) );
  NAND2_X1 U84 ( .A1(n342), .A2(n338), .ZN(n344) );
  OAI21_X1 U85 ( .B1(A[9]), .B2(n326), .A(A[10]), .ZN(n338) );
  INV_X1 U86 ( .A(n378), .ZN(n326) );
  INV_X1 U87 ( .A(A[9]), .ZN(n318) );
  INV_X1 U88 ( .A(A[12]), .ZN(n319) );
  INV_X1 U89 ( .A(A[13]), .ZN(n320) );
endmodule


module BOOTH_ENCODER_WIDTH16_3 ( A, b, vp );
  input [15:0] A;
  input [2:0] b;
  output [16:0] vp;
  wire   \notA[0] , n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388;
  assign \notA[0]  = A[0];

  XOR2_X1 U90 ( .A(n378), .B(A[9]), .Z(n388) );
  NAND3_X1 U91 ( .A1(n324), .A2(n318), .A3(n378), .ZN(n342) );
  NOR2_X2 U3 ( .A1(n339), .A2(b[2]), .ZN(n383) );
  NOR2_X2 U4 ( .A1(n340), .A2(b[2]), .ZN(n380) );
  OR2_X1 U5 ( .A1(n340), .A2(n358), .ZN(n387) );
  INV_X1 U6 ( .A(n348), .ZN(n321) );
  INV_X1 U7 ( .A(n385), .ZN(n335) );
  OAI21_X1 U8 ( .B1(n346), .B2(n319), .A(n348), .ZN(n350) );
  OAI21_X1 U9 ( .B1(n321), .B2(n320), .A(n353), .ZN(n352) );
  INV_X1 U10 ( .A(n360), .ZN(n330) );
  INV_X1 U11 ( .A(n369), .ZN(n328) );
  NAND2_X1 U12 ( .A1(n321), .A2(n320), .ZN(n353) );
  NAND2_X1 U13 ( .A1(n346), .A2(n319), .ZN(n348) );
  AOI21_X1 U14 ( .B1(n379), .B2(A[8]), .A(n378), .ZN(n384) );
  NOR2_X1 U15 ( .A1(n379), .A2(A[8]), .ZN(n378) );
  OAI221_X1 U16 ( .B1(n387), .B2(n355), .C1(n335), .C2(n352), .A(n351), .ZN(
        vp[14]) );
  AOI22_X1 U17 ( .A1(A[13]), .A2(n383), .B1(A[14]), .B2(n380), .ZN(n351) );
  OAI221_X1 U18 ( .B1(n387), .B2(n368), .C1(n335), .C2(n331), .A(n365), .ZN(
        vp[3]) );
  AOI22_X1 U19 ( .A1(A[2]), .A2(n383), .B1(A[3]), .B2(n380), .ZN(n365) );
  OAI221_X1 U20 ( .B1(n387), .B2(n373), .C1(n335), .C2(n368), .A(n367), .ZN(
        vp[4]) );
  AOI22_X1 U21 ( .A1(A[3]), .A2(n383), .B1(A[4]), .B2(n380), .ZN(n367) );
  OAI221_X1 U22 ( .B1(n387), .B2(n329), .C1(n335), .C2(n373), .A(n372), .ZN(
        vp[5]) );
  AOI22_X1 U23 ( .A1(A[4]), .A2(n383), .B1(A[5]), .B2(n380), .ZN(n372) );
  OAI221_X1 U24 ( .B1(n387), .B2(n377), .C1(n335), .C2(n329), .A(n374), .ZN(
        vp[6]) );
  AOI22_X1 U25 ( .A1(A[5]), .A2(n383), .B1(A[6]), .B2(n380), .ZN(n374) );
  OAI221_X1 U26 ( .B1(n387), .B2(n382), .C1(n335), .C2(n377), .A(n376), .ZN(
        vp[7]) );
  AOI22_X1 U27 ( .A1(A[6]), .A2(n383), .B1(A[7]), .B2(n380), .ZN(n376) );
  OAI221_X1 U28 ( .B1(n387), .B2(n344), .C1(n334), .C2(n324), .A(n325), .ZN(
        vp[10]) );
  INV_X1 U29 ( .A(n341), .ZN(n325) );
  OAI22_X1 U30 ( .A1(n318), .A2(n336), .B1(n388), .B2(n335), .ZN(n341) );
  OAI221_X1 U31 ( .B1(n387), .B2(n322), .C1(n336), .C2(n324), .A(n345), .ZN(
        vp[11]) );
  AOI22_X1 U32 ( .A1(n323), .A2(n385), .B1(A[11]), .B2(n380), .ZN(n345) );
  INV_X1 U33 ( .A(n344), .ZN(n323) );
  OAI221_X1 U34 ( .B1(n387), .B2(n350), .C1(n335), .C2(n322), .A(n347), .ZN(
        vp[12]) );
  AOI22_X1 U35 ( .A1(A[11]), .A2(n383), .B1(A[12]), .B2(n380), .ZN(n347) );
  OAI221_X1 U36 ( .B1(n387), .B2(n352), .C1(n335), .C2(n350), .A(n349), .ZN(
        vp[13]) );
  AOI22_X1 U37 ( .A1(A[12]), .A2(n383), .B1(A[13]), .B2(n380), .ZN(n349) );
  OAI221_X1 U38 ( .B1(n387), .B2(n357), .C1(n335), .C2(n355), .A(n354), .ZN(
        vp[15]) );
  AOI22_X1 U39 ( .A1(A[14]), .A2(n383), .B1(A[15]), .B2(n380), .ZN(n354) );
  OAI221_X1 U40 ( .B1(n388), .B2(n387), .C1(n318), .C2(n334), .A(n386), .ZN(
        vp[9]) );
  AOI22_X1 U41 ( .A1(n385), .A2(n384), .B1(n383), .B2(A[8]), .ZN(n386) );
  OAI221_X1 U42 ( .B1(n327), .B2(n387), .C1(n335), .C2(n382), .A(n381), .ZN(
        vp[8]) );
  INV_X1 U43 ( .A(n384), .ZN(n327) );
  AOI22_X1 U44 ( .A1(A[7]), .A2(n383), .B1(n380), .B2(A[8]), .ZN(n381) );
  NOR2_X1 U45 ( .A1(n358), .A2(n337), .ZN(n385) );
  INV_X1 U46 ( .A(n340), .ZN(n337) );
  NOR2_X1 U47 ( .A1(n342), .A2(A[11]), .ZN(n346) );
  XNOR2_X1 U48 ( .A(n353), .B(A[14]), .ZN(n355) );
  XNOR2_X1 U49 ( .A(n330), .B(A[3]), .ZN(n368) );
  XNOR2_X1 U50 ( .A(n328), .B(A[6]), .ZN(n377) );
  NOR2_X1 U51 ( .A1(n361), .A2(A[2]), .ZN(n360) );
  NOR2_X1 U52 ( .A1(n370), .A2(A[5]), .ZN(n369) );
  XOR2_X1 U53 ( .A(n317), .B(A[15]), .Z(n357) );
  NOR2_X1 U54 ( .A1(n353), .A2(A[14]), .ZN(n317) );
  AOI21_X1 U55 ( .B1(n334), .B2(n387), .A(n333), .ZN(vp[0]) );
  OAI21_X1 U56 ( .B1(n332), .B2(n333), .A(n361), .ZN(n364) );
  OAI21_X1 U57 ( .B1(n358), .B2(n357), .A(n356), .ZN(vp[16]) );
  OAI21_X1 U58 ( .B1(n383), .B2(n380), .A(A[15]), .ZN(n356) );
  INV_X1 U59 ( .A(n380), .ZN(n334) );
  NAND2_X1 U60 ( .A1(n332), .A2(n333), .ZN(n361) );
  INV_X1 U61 ( .A(n383), .ZN(n336) );
  NAND2_X1 U62 ( .A1(n370), .A2(n366), .ZN(n373) );
  OAI21_X1 U63 ( .B1(A[3]), .B2(n330), .A(A[4]), .ZN(n366) );
  NAND2_X1 U64 ( .A1(n379), .A2(n375), .ZN(n382) );
  OAI21_X1 U65 ( .B1(A[6]), .B2(n328), .A(A[7]), .ZN(n375) );
  OR3_X1 U66 ( .A1(A[3]), .A2(A[4]), .A3(n330), .ZN(n370) );
  OR3_X1 U67 ( .A1(A[6]), .A2(A[7]), .A3(n328), .ZN(n379) );
  INV_X1 U68 ( .A(n362), .ZN(n331) );
  AOI21_X1 U69 ( .B1(n361), .B2(A[2]), .A(n360), .ZN(n362) );
  INV_X1 U70 ( .A(n371), .ZN(n329) );
  AOI21_X1 U71 ( .B1(n370), .B2(A[5]), .A(n369), .ZN(n371) );
  INV_X1 U72 ( .A(n343), .ZN(n322) );
  AOI21_X1 U73 ( .B1(n342), .B2(A[11]), .A(n346), .ZN(n343) );
  OAI21_X1 U74 ( .B1(b[1]), .B2(b[0]), .A(n339), .ZN(n340) );
  OAI221_X1 U75 ( .B1(n387), .B2(n364), .C1(n334), .C2(n332), .A(n359), .ZN(
        vp[1]) );
  OAI21_X1 U76 ( .B1(n383), .B2(n385), .A(\notA[0] ), .ZN(n359) );
  OAI221_X1 U77 ( .B1(n387), .B2(n331), .C1(n335), .C2(n364), .A(n363), .ZN(
        vp[2]) );
  AOI22_X1 U78 ( .A1(A[1]), .A2(n383), .B1(A[2]), .B2(n380), .ZN(n363) );
  INV_X1 U79 ( .A(\notA[0] ), .ZN(n333) );
  INV_X1 U80 ( .A(A[1]), .ZN(n332) );
  INV_X1 U81 ( .A(A[10]), .ZN(n324) );
  NAND2_X1 U82 ( .A1(b[1]), .A2(b[0]), .ZN(n339) );
  NAND2_X1 U83 ( .A1(b[2]), .A2(n339), .ZN(n358) );
  NAND2_X1 U84 ( .A1(n342), .A2(n338), .ZN(n344) );
  OAI21_X1 U85 ( .B1(A[9]), .B2(n326), .A(A[10]), .ZN(n338) );
  INV_X1 U86 ( .A(n378), .ZN(n326) );
  INV_X1 U87 ( .A(A[9]), .ZN(n318) );
  INV_X1 U88 ( .A(A[12]), .ZN(n319) );
  INV_X1 U89 ( .A(A[13]), .ZN(n320) );
endmodule


module BOOTH_ENCODER_WIDTH16_2 ( A, b, vp );
  input [15:0] A;
  input [2:0] b;
  output [16:0] vp;
  wire   \notA[0] , n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387;
  assign \notA[0]  = A[0];

  XOR2_X1 U90 ( .A(n377), .B(A[9]), .Z(n387) );
  NAND3_X1 U91 ( .A1(n323), .A2(n317), .A3(n377), .ZN(n341) );
  NOR2_X2 U3 ( .A1(n338), .A2(b[2]), .ZN(n382) );
  NOR2_X2 U4 ( .A1(n339), .A2(b[2]), .ZN(n379) );
  OR2_X1 U5 ( .A1(n339), .A2(n357), .ZN(n386) );
  INV_X1 U6 ( .A(n347), .ZN(n320) );
  INV_X1 U7 ( .A(n384), .ZN(n334) );
  OAI21_X1 U8 ( .B1(n345), .B2(n318), .A(n347), .ZN(n349) );
  OAI21_X1 U9 ( .B1(n320), .B2(n319), .A(n352), .ZN(n351) );
  INV_X1 U10 ( .A(n359), .ZN(n329) );
  INV_X1 U11 ( .A(n368), .ZN(n327) );
  NAND2_X1 U12 ( .A1(n320), .A2(n319), .ZN(n352) );
  NAND2_X1 U13 ( .A1(n345), .A2(n318), .ZN(n347) );
  AOI21_X1 U14 ( .B1(n378), .B2(A[8]), .A(n377), .ZN(n383) );
  NOR2_X1 U15 ( .A1(n378), .A2(A[8]), .ZN(n377) );
  OAI221_X1 U16 ( .B1(n386), .B2(n354), .C1(n334), .C2(n351), .A(n350), .ZN(
        vp[14]) );
  AOI22_X1 U17 ( .A1(A[13]), .A2(n382), .B1(A[14]), .B2(n379), .ZN(n350) );
  OAI221_X1 U18 ( .B1(n386), .B2(n367), .C1(n334), .C2(n330), .A(n364), .ZN(
        vp[3]) );
  AOI22_X1 U19 ( .A1(A[2]), .A2(n382), .B1(A[3]), .B2(n379), .ZN(n364) );
  OAI221_X1 U20 ( .B1(n386), .B2(n372), .C1(n334), .C2(n367), .A(n366), .ZN(
        vp[4]) );
  AOI22_X1 U21 ( .A1(A[3]), .A2(n382), .B1(A[4]), .B2(n379), .ZN(n366) );
  OAI221_X1 U22 ( .B1(n386), .B2(n328), .C1(n334), .C2(n372), .A(n371), .ZN(
        vp[5]) );
  AOI22_X1 U23 ( .A1(A[4]), .A2(n382), .B1(A[5]), .B2(n379), .ZN(n371) );
  OAI221_X1 U24 ( .B1(n386), .B2(n376), .C1(n334), .C2(n328), .A(n373), .ZN(
        vp[6]) );
  AOI22_X1 U25 ( .A1(A[5]), .A2(n382), .B1(A[6]), .B2(n379), .ZN(n373) );
  OAI221_X1 U26 ( .B1(n386), .B2(n381), .C1(n334), .C2(n376), .A(n375), .ZN(
        vp[7]) );
  AOI22_X1 U27 ( .A1(A[6]), .A2(n382), .B1(A[7]), .B2(n379), .ZN(n375) );
  OAI221_X1 U28 ( .B1(n386), .B2(n343), .C1(n333), .C2(n323), .A(n324), .ZN(
        vp[10]) );
  INV_X1 U29 ( .A(n340), .ZN(n324) );
  OAI22_X1 U30 ( .A1(n317), .A2(n335), .B1(n387), .B2(n334), .ZN(n340) );
  OAI221_X1 U31 ( .B1(n386), .B2(n321), .C1(n335), .C2(n323), .A(n344), .ZN(
        vp[11]) );
  AOI22_X1 U32 ( .A1(n322), .A2(n384), .B1(A[11]), .B2(n379), .ZN(n344) );
  INV_X1 U33 ( .A(n343), .ZN(n322) );
  OAI221_X1 U34 ( .B1(n386), .B2(n349), .C1(n334), .C2(n321), .A(n346), .ZN(
        vp[12]) );
  AOI22_X1 U35 ( .A1(A[11]), .A2(n382), .B1(A[12]), .B2(n379), .ZN(n346) );
  OAI221_X1 U36 ( .B1(n386), .B2(n351), .C1(n334), .C2(n349), .A(n348), .ZN(
        vp[13]) );
  AOI22_X1 U37 ( .A1(A[12]), .A2(n382), .B1(A[13]), .B2(n379), .ZN(n348) );
  OAI221_X1 U38 ( .B1(n386), .B2(n356), .C1(n334), .C2(n354), .A(n353), .ZN(
        vp[15]) );
  AOI22_X1 U39 ( .A1(A[14]), .A2(n382), .B1(A[15]), .B2(n379), .ZN(n353) );
  OAI221_X1 U40 ( .B1(n387), .B2(n386), .C1(n317), .C2(n333), .A(n385), .ZN(
        vp[9]) );
  AOI22_X1 U41 ( .A1(n384), .A2(n383), .B1(n382), .B2(A[8]), .ZN(n385) );
  OAI221_X1 U42 ( .B1(n326), .B2(n386), .C1(n334), .C2(n381), .A(n380), .ZN(
        vp[8]) );
  INV_X1 U43 ( .A(n383), .ZN(n326) );
  AOI22_X1 U44 ( .A1(A[7]), .A2(n382), .B1(n379), .B2(A[8]), .ZN(n380) );
  NOR2_X1 U45 ( .A1(n357), .A2(n336), .ZN(n384) );
  INV_X1 U46 ( .A(n339), .ZN(n336) );
  NOR2_X1 U47 ( .A1(n341), .A2(A[11]), .ZN(n345) );
  XNOR2_X1 U48 ( .A(n352), .B(A[14]), .ZN(n354) );
  XNOR2_X1 U49 ( .A(n329), .B(A[3]), .ZN(n367) );
  XNOR2_X1 U50 ( .A(n327), .B(A[6]), .ZN(n376) );
  NOR2_X1 U51 ( .A1(n360), .A2(A[2]), .ZN(n359) );
  NOR2_X1 U52 ( .A1(n369), .A2(A[5]), .ZN(n368) );
  XOR2_X1 U53 ( .A(n316), .B(A[15]), .Z(n356) );
  NOR2_X1 U54 ( .A1(n352), .A2(A[14]), .ZN(n316) );
  AOI21_X1 U55 ( .B1(n333), .B2(n386), .A(n332), .ZN(vp[0]) );
  OAI21_X1 U56 ( .B1(n331), .B2(n332), .A(n360), .ZN(n363) );
  OAI21_X1 U57 ( .B1(n357), .B2(n356), .A(n355), .ZN(vp[16]) );
  OAI21_X1 U58 ( .B1(n382), .B2(n379), .A(A[15]), .ZN(n355) );
  INV_X1 U59 ( .A(n379), .ZN(n333) );
  NAND2_X1 U60 ( .A1(n331), .A2(n332), .ZN(n360) );
  INV_X1 U61 ( .A(n382), .ZN(n335) );
  NAND2_X1 U62 ( .A1(n369), .A2(n365), .ZN(n372) );
  OAI21_X1 U63 ( .B1(A[3]), .B2(n329), .A(A[4]), .ZN(n365) );
  NAND2_X1 U64 ( .A1(n378), .A2(n374), .ZN(n381) );
  OAI21_X1 U65 ( .B1(A[6]), .B2(n327), .A(A[7]), .ZN(n374) );
  OR3_X1 U66 ( .A1(A[3]), .A2(A[4]), .A3(n329), .ZN(n369) );
  OR3_X1 U67 ( .A1(A[6]), .A2(A[7]), .A3(n327), .ZN(n378) );
  INV_X1 U68 ( .A(n361), .ZN(n330) );
  AOI21_X1 U69 ( .B1(n360), .B2(A[2]), .A(n359), .ZN(n361) );
  INV_X1 U70 ( .A(n370), .ZN(n328) );
  AOI21_X1 U71 ( .B1(n369), .B2(A[5]), .A(n368), .ZN(n370) );
  INV_X1 U72 ( .A(n342), .ZN(n321) );
  AOI21_X1 U73 ( .B1(n341), .B2(A[11]), .A(n345), .ZN(n342) );
  OAI21_X1 U74 ( .B1(b[1]), .B2(b[0]), .A(n338), .ZN(n339) );
  OAI221_X1 U75 ( .B1(n386), .B2(n363), .C1(n333), .C2(n331), .A(n358), .ZN(
        vp[1]) );
  OAI21_X1 U76 ( .B1(n382), .B2(n384), .A(\notA[0] ), .ZN(n358) );
  OAI221_X1 U77 ( .B1(n386), .B2(n330), .C1(n334), .C2(n363), .A(n362), .ZN(
        vp[2]) );
  AOI22_X1 U78 ( .A1(A[1]), .A2(n382), .B1(A[2]), .B2(n379), .ZN(n362) );
  INV_X1 U79 ( .A(\notA[0] ), .ZN(n332) );
  INV_X1 U80 ( .A(A[1]), .ZN(n331) );
  INV_X1 U81 ( .A(A[10]), .ZN(n323) );
  NAND2_X1 U82 ( .A1(b[1]), .A2(b[0]), .ZN(n338) );
  NAND2_X1 U83 ( .A1(b[2]), .A2(n338), .ZN(n357) );
  NAND2_X1 U84 ( .A1(n341), .A2(n337), .ZN(n343) );
  OAI21_X1 U85 ( .B1(A[9]), .B2(n325), .A(A[10]), .ZN(n337) );
  INV_X1 U86 ( .A(n377), .ZN(n325) );
  INV_X1 U87 ( .A(A[9]), .ZN(n317) );
  INV_X1 U88 ( .A(A[12]), .ZN(n318) );
  INV_X1 U89 ( .A(A[13]), .ZN(n319) );
endmodule


module BOOTH_ENCODER_WIDTH16_1 ( A, b, vp );
  input [15:0] A;
  input [2:0] b;
  output [16:0] vp;
  wire   \notA[0] , n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387;
  assign \notA[0]  = A[0];

  XOR2_X1 U90 ( .A(n377), .B(A[9]), .Z(n387) );
  NAND3_X1 U91 ( .A1(n323), .A2(n317), .A3(n377), .ZN(n341) );
  NOR2_X2 U3 ( .A1(n338), .A2(b[2]), .ZN(n382) );
  NOR2_X2 U4 ( .A1(n339), .A2(b[2]), .ZN(n379) );
  OR2_X1 U5 ( .A1(n339), .A2(n357), .ZN(n386) );
  INV_X1 U6 ( .A(n347), .ZN(n320) );
  INV_X1 U7 ( .A(n384), .ZN(n334) );
  OAI21_X1 U8 ( .B1(n345), .B2(n318), .A(n347), .ZN(n349) );
  OAI21_X1 U9 ( .B1(n320), .B2(n319), .A(n352), .ZN(n351) );
  INV_X1 U10 ( .A(n359), .ZN(n329) );
  INV_X1 U11 ( .A(n368), .ZN(n327) );
  NAND2_X1 U12 ( .A1(n320), .A2(n319), .ZN(n352) );
  NAND2_X1 U13 ( .A1(n345), .A2(n318), .ZN(n347) );
  AOI21_X1 U14 ( .B1(n378), .B2(A[8]), .A(n377), .ZN(n383) );
  NOR2_X1 U15 ( .A1(n378), .A2(A[8]), .ZN(n377) );
  OAI221_X1 U16 ( .B1(n386), .B2(n354), .C1(n334), .C2(n351), .A(n350), .ZN(
        vp[14]) );
  AOI22_X1 U17 ( .A1(A[13]), .A2(n382), .B1(A[14]), .B2(n379), .ZN(n350) );
  OAI221_X1 U18 ( .B1(n386), .B2(n367), .C1(n334), .C2(n330), .A(n364), .ZN(
        vp[3]) );
  AOI22_X1 U19 ( .A1(A[2]), .A2(n382), .B1(A[3]), .B2(n379), .ZN(n364) );
  OAI221_X1 U20 ( .B1(n386), .B2(n372), .C1(n334), .C2(n367), .A(n366), .ZN(
        vp[4]) );
  AOI22_X1 U21 ( .A1(A[3]), .A2(n382), .B1(A[4]), .B2(n379), .ZN(n366) );
  OAI221_X1 U22 ( .B1(n386), .B2(n328), .C1(n334), .C2(n372), .A(n371), .ZN(
        vp[5]) );
  AOI22_X1 U23 ( .A1(A[4]), .A2(n382), .B1(A[5]), .B2(n379), .ZN(n371) );
  OAI221_X1 U24 ( .B1(n386), .B2(n376), .C1(n334), .C2(n328), .A(n373), .ZN(
        vp[6]) );
  AOI22_X1 U25 ( .A1(A[5]), .A2(n382), .B1(A[6]), .B2(n379), .ZN(n373) );
  OAI221_X1 U26 ( .B1(n386), .B2(n381), .C1(n334), .C2(n376), .A(n375), .ZN(
        vp[7]) );
  AOI22_X1 U27 ( .A1(A[6]), .A2(n382), .B1(A[7]), .B2(n379), .ZN(n375) );
  OAI221_X1 U28 ( .B1(n386), .B2(n343), .C1(n333), .C2(n323), .A(n324), .ZN(
        vp[10]) );
  INV_X1 U29 ( .A(n340), .ZN(n324) );
  OAI22_X1 U30 ( .A1(n317), .A2(n335), .B1(n387), .B2(n334), .ZN(n340) );
  OAI221_X1 U31 ( .B1(n386), .B2(n321), .C1(n335), .C2(n323), .A(n344), .ZN(
        vp[11]) );
  AOI22_X1 U32 ( .A1(n322), .A2(n384), .B1(A[11]), .B2(n379), .ZN(n344) );
  INV_X1 U33 ( .A(n343), .ZN(n322) );
  OAI221_X1 U34 ( .B1(n386), .B2(n349), .C1(n334), .C2(n321), .A(n346), .ZN(
        vp[12]) );
  AOI22_X1 U35 ( .A1(A[11]), .A2(n382), .B1(A[12]), .B2(n379), .ZN(n346) );
  OAI221_X1 U36 ( .B1(n386), .B2(n351), .C1(n334), .C2(n349), .A(n348), .ZN(
        vp[13]) );
  AOI22_X1 U37 ( .A1(A[12]), .A2(n382), .B1(A[13]), .B2(n379), .ZN(n348) );
  OAI221_X1 U38 ( .B1(n386), .B2(n356), .C1(n334), .C2(n354), .A(n353), .ZN(
        vp[15]) );
  AOI22_X1 U39 ( .A1(A[14]), .A2(n382), .B1(A[15]), .B2(n379), .ZN(n353) );
  OAI221_X1 U40 ( .B1(n387), .B2(n386), .C1(n317), .C2(n333), .A(n385), .ZN(
        vp[9]) );
  AOI22_X1 U41 ( .A1(n384), .A2(n383), .B1(n382), .B2(A[8]), .ZN(n385) );
  OAI221_X1 U42 ( .B1(n326), .B2(n386), .C1(n334), .C2(n381), .A(n380), .ZN(
        vp[8]) );
  INV_X1 U43 ( .A(n383), .ZN(n326) );
  AOI22_X1 U44 ( .A1(A[7]), .A2(n382), .B1(n379), .B2(A[8]), .ZN(n380) );
  NOR2_X1 U45 ( .A1(n357), .A2(n336), .ZN(n384) );
  INV_X1 U46 ( .A(n339), .ZN(n336) );
  NOR2_X1 U47 ( .A1(n341), .A2(A[11]), .ZN(n345) );
  XNOR2_X1 U48 ( .A(n352), .B(A[14]), .ZN(n354) );
  XNOR2_X1 U49 ( .A(n329), .B(A[3]), .ZN(n367) );
  XNOR2_X1 U50 ( .A(n327), .B(A[6]), .ZN(n376) );
  NOR2_X1 U51 ( .A1(n360), .A2(A[2]), .ZN(n359) );
  NOR2_X1 U52 ( .A1(n369), .A2(A[5]), .ZN(n368) );
  XOR2_X1 U53 ( .A(n316), .B(A[15]), .Z(n356) );
  NOR2_X1 U54 ( .A1(n352), .A2(A[14]), .ZN(n316) );
  AOI21_X1 U55 ( .B1(n333), .B2(n386), .A(n332), .ZN(vp[0]) );
  OAI21_X1 U56 ( .B1(n331), .B2(n332), .A(n360), .ZN(n363) );
  OAI21_X1 U57 ( .B1(n357), .B2(n356), .A(n355), .ZN(vp[16]) );
  OAI21_X1 U58 ( .B1(n382), .B2(n379), .A(A[15]), .ZN(n355) );
  INV_X1 U59 ( .A(n379), .ZN(n333) );
  NAND2_X1 U60 ( .A1(n331), .A2(n332), .ZN(n360) );
  INV_X1 U61 ( .A(n382), .ZN(n335) );
  NAND2_X1 U62 ( .A1(n369), .A2(n365), .ZN(n372) );
  OAI21_X1 U63 ( .B1(A[3]), .B2(n329), .A(A[4]), .ZN(n365) );
  NAND2_X1 U64 ( .A1(n378), .A2(n374), .ZN(n381) );
  OAI21_X1 U65 ( .B1(A[6]), .B2(n327), .A(A[7]), .ZN(n374) );
  OR3_X1 U66 ( .A1(A[3]), .A2(A[4]), .A3(n329), .ZN(n369) );
  OR3_X1 U67 ( .A1(A[6]), .A2(A[7]), .A3(n327), .ZN(n378) );
  INV_X1 U68 ( .A(n361), .ZN(n330) );
  AOI21_X1 U69 ( .B1(n360), .B2(A[2]), .A(n359), .ZN(n361) );
  INV_X1 U70 ( .A(n370), .ZN(n328) );
  AOI21_X1 U71 ( .B1(n369), .B2(A[5]), .A(n368), .ZN(n370) );
  INV_X1 U72 ( .A(n342), .ZN(n321) );
  AOI21_X1 U73 ( .B1(n341), .B2(A[11]), .A(n345), .ZN(n342) );
  OAI21_X1 U74 ( .B1(b[1]), .B2(b[0]), .A(n338), .ZN(n339) );
  OAI221_X1 U75 ( .B1(n386), .B2(n363), .C1(n333), .C2(n331), .A(n358), .ZN(
        vp[1]) );
  OAI21_X1 U76 ( .B1(n382), .B2(n384), .A(\notA[0] ), .ZN(n358) );
  OAI221_X1 U77 ( .B1(n386), .B2(n330), .C1(n334), .C2(n363), .A(n362), .ZN(
        vp[2]) );
  AOI22_X1 U78 ( .A1(A[1]), .A2(n382), .B1(A[2]), .B2(n379), .ZN(n362) );
  INV_X1 U79 ( .A(\notA[0] ), .ZN(n332) );
  INV_X1 U80 ( .A(A[1]), .ZN(n331) );
  INV_X1 U81 ( .A(A[10]), .ZN(n323) );
  NAND2_X1 U82 ( .A1(b[1]), .A2(b[0]), .ZN(n338) );
  NAND2_X1 U83 ( .A1(b[2]), .A2(n338), .ZN(n357) );
  NAND2_X1 U84 ( .A1(n341), .A2(n337), .ZN(n343) );
  OAI21_X1 U85 ( .B1(A[9]), .B2(n325), .A(A[10]), .ZN(n337) );
  INV_X1 U86 ( .A(n377), .ZN(n325) );
  INV_X1 U87 ( .A(A[9]), .ZN(n317) );
  INV_X1 U88 ( .A(A[12]), .ZN(n318) );
  INV_X1 U89 ( .A(A[13]), .ZN(n319) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n2) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_MUL_WIDTH16_0 ( A, B, Ci, S, Partial, Co );
  input [16:0] A;
  input [16:0] B;
  output [16:0] S;
  output [1:0] Partial;
  input Ci;
  output Co;

  wire   [16:2] res;
  wire   [16:1] carry;
  assign S[14] = res[16];
  assign S[15] = res[16];
  assign S[16] = res[16];
  assign S[13] = res[15];
  assign S[12] = res[14];
  assign S[11] = res[13];
  assign S[10] = res[12];
  assign S[9] = res[11];
  assign S[8] = res[10];
  assign S[7] = res[9];
  assign S[6] = res[8];
  assign S[5] = res[7];
  assign S[4] = res[6];
  assign S[3] = res[5];
  assign S[2] = res[4];
  assign S[1] = res[3];
  assign S[0] = res[2];

  FA_0 sum0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(Partial[0]), .Co(carry[1]) );
  FA_199 sumI_1 ( .A(A[1]), .B(B[1]), .Ci(carry[1]), .S(Partial[1]), .Co(
        carry[2]) );
  FA_198 sumI_2 ( .A(A[2]), .B(B[2]), .Ci(carry[2]), .S(res[2]), .Co(carry[3])
         );
  FA_197 sumI_3 ( .A(A[3]), .B(B[3]), .Ci(carry[3]), .S(res[3]), .Co(carry[4])
         );
  FA_196 sumI_4 ( .A(A[4]), .B(B[4]), .Ci(carry[4]), .S(res[4]), .Co(carry[5])
         );
  FA_195 sumI_5 ( .A(A[5]), .B(B[5]), .Ci(carry[5]), .S(res[5]), .Co(carry[6])
         );
  FA_194 sumI_6 ( .A(A[6]), .B(B[6]), .Ci(carry[6]), .S(res[6]), .Co(carry[7])
         );
  FA_193 sumI_7 ( .A(A[7]), .B(B[7]), .Ci(carry[7]), .S(res[7]), .Co(carry[8])
         );
  FA_192 sumI_8 ( .A(A[8]), .B(B[8]), .Ci(carry[8]), .S(res[8]), .Co(carry[9])
         );
  FA_191 sumI_9 ( .A(A[9]), .B(B[9]), .Ci(carry[9]), .S(res[9]), .Co(carry[10]) );
  FA_190 sumI_10 ( .A(A[10]), .B(B[10]), .Ci(carry[10]), .S(res[10]), .Co(
        carry[11]) );
  FA_189 sumI_11 ( .A(A[11]), .B(B[11]), .Ci(carry[11]), .S(res[11]), .Co(
        carry[12]) );
  FA_188 sumI_12 ( .A(A[12]), .B(B[12]), .Ci(carry[12]), .S(res[12]), .Co(
        carry[13]) );
  FA_187 sumI_13 ( .A(A[13]), .B(B[13]), .Ci(carry[13]), .S(res[13]), .Co(
        carry[14]) );
  FA_186 sumI_14 ( .A(A[14]), .B(B[14]), .Ci(carry[14]), .S(res[14]), .Co(
        carry[15]) );
  FA_185 sumI_15 ( .A(A[15]), .B(B[15]), .Ci(carry[15]), .S(res[15]), .Co(
        carry[16]) );
  FA_184 sumTH ( .A(A[16]), .B(B[16]), .Ci(carry[16]), .S(res[16]), .Co(Co) );
endmodule


module FA_183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_MUL_WIDTH16_7 ( A, B, Ci, S, Partial, Co );
  input [16:0] A;
  input [16:0] B;
  output [16:0] S;
  output [1:0] Partial;
  input Ci;
  output Co;

  wire   [16:2] res;
  wire   [16:1] carry;
  assign S[14] = res[16];
  assign S[15] = res[16];
  assign S[16] = res[16];
  assign S[13] = res[15];
  assign S[12] = res[14];
  assign S[11] = res[13];
  assign S[10] = res[12];
  assign S[9] = res[11];
  assign S[8] = res[10];
  assign S[7] = res[9];
  assign S[6] = res[8];
  assign S[5] = res[7];
  assign S[4] = res[6];
  assign S[3] = res[5];
  assign S[2] = res[4];
  assign S[1] = res[3];
  assign S[0] = res[2];

  FA_183 sum0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(Partial[0]), .Co(carry[1]) );
  FA_182 sumI_1 ( .A(A[1]), .B(B[1]), .Ci(carry[1]), .S(Partial[1]), .Co(
        carry[2]) );
  FA_181 sumI_2 ( .A(A[2]), .B(B[2]), .Ci(carry[2]), .S(res[2]), .Co(carry[3])
         );
  FA_180 sumI_3 ( .A(A[3]), .B(B[3]), .Ci(carry[3]), .S(res[3]), .Co(carry[4])
         );
  FA_179 sumI_4 ( .A(A[4]), .B(B[4]), .Ci(carry[4]), .S(res[4]), .Co(carry[5])
         );
  FA_178 sumI_5 ( .A(A[5]), .B(B[5]), .Ci(carry[5]), .S(res[5]), .Co(carry[6])
         );
  FA_177 sumI_6 ( .A(A[6]), .B(B[6]), .Ci(carry[6]), .S(res[6]), .Co(carry[7])
         );
  FA_176 sumI_7 ( .A(A[7]), .B(B[7]), .Ci(carry[7]), .S(res[7]), .Co(carry[8])
         );
  FA_175 sumI_8 ( .A(A[8]), .B(B[8]), .Ci(carry[8]), .S(res[8]), .Co(carry[9])
         );
  FA_174 sumI_9 ( .A(A[9]), .B(B[9]), .Ci(carry[9]), .S(res[9]), .Co(carry[10]) );
  FA_173 sumI_10 ( .A(A[10]), .B(B[10]), .Ci(carry[10]), .S(res[10]), .Co(
        carry[11]) );
  FA_172 sumI_11 ( .A(A[11]), .B(B[11]), .Ci(carry[11]), .S(res[11]), .Co(
        carry[12]) );
  FA_171 sumI_12 ( .A(A[12]), .B(B[12]), .Ci(carry[12]), .S(res[12]), .Co(
        carry[13]) );
  FA_170 sumI_13 ( .A(A[13]), .B(B[13]), .Ci(carry[13]), .S(res[13]), .Co(
        carry[14]) );
  FA_169 sumI_14 ( .A(A[14]), .B(B[14]), .Ci(carry[14]), .S(res[14]), .Co(
        carry[15]) );
  FA_168 sumI_15 ( .A(A[15]), .B(B[15]), .Ci(carry[15]), .S(res[15]), .Co(
        carry[16]) );
  FA_167 sumTH ( .A(A[16]), .B(B[16]), .Ci(carry[16]), .S(res[16]), .Co(Co) );
endmodule


module FA_166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_MUL_WIDTH16_6 ( A, B, Ci, S, Partial, Co );
  input [16:0] A;
  input [16:0] B;
  output [16:0] S;
  output [1:0] Partial;
  input Ci;
  output Co;

  wire   [16:2] res;
  wire   [16:1] carry;
  assign S[14] = res[16];
  assign S[15] = res[16];
  assign S[16] = res[16];
  assign S[13] = res[15];
  assign S[12] = res[14];
  assign S[11] = res[13];
  assign S[10] = res[12];
  assign S[9] = res[11];
  assign S[8] = res[10];
  assign S[7] = res[9];
  assign S[6] = res[8];
  assign S[5] = res[7];
  assign S[4] = res[6];
  assign S[3] = res[5];
  assign S[2] = res[4];
  assign S[1] = res[3];
  assign S[0] = res[2];

  FA_166 sum0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(Partial[0]), .Co(carry[1]) );
  FA_165 sumI_1 ( .A(A[1]), .B(B[1]), .Ci(carry[1]), .S(Partial[1]), .Co(
        carry[2]) );
  FA_164 sumI_2 ( .A(A[2]), .B(B[2]), .Ci(carry[2]), .S(res[2]), .Co(carry[3])
         );
  FA_163 sumI_3 ( .A(A[3]), .B(B[3]), .Ci(carry[3]), .S(res[3]), .Co(carry[4])
         );
  FA_162 sumI_4 ( .A(A[4]), .B(B[4]), .Ci(carry[4]), .S(res[4]), .Co(carry[5])
         );
  FA_161 sumI_5 ( .A(A[5]), .B(B[5]), .Ci(carry[5]), .S(res[5]), .Co(carry[6])
         );
  FA_160 sumI_6 ( .A(A[6]), .B(B[6]), .Ci(carry[6]), .S(res[6]), .Co(carry[7])
         );
  FA_159 sumI_7 ( .A(A[7]), .B(B[7]), .Ci(carry[7]), .S(res[7]), .Co(carry[8])
         );
  FA_158 sumI_8 ( .A(A[8]), .B(B[8]), .Ci(carry[8]), .S(res[8]), .Co(carry[9])
         );
  FA_157 sumI_9 ( .A(A[9]), .B(B[9]), .Ci(carry[9]), .S(res[9]), .Co(carry[10]) );
  FA_156 sumI_10 ( .A(A[10]), .B(B[10]), .Ci(carry[10]), .S(res[10]), .Co(
        carry[11]) );
  FA_155 sumI_11 ( .A(A[11]), .B(B[11]), .Ci(carry[11]), .S(res[11]), .Co(
        carry[12]) );
  FA_154 sumI_12 ( .A(A[12]), .B(B[12]), .Ci(carry[12]), .S(res[12]), .Co(
        carry[13]) );
  FA_153 sumI_13 ( .A(A[13]), .B(B[13]), .Ci(carry[13]), .S(res[13]), .Co(
        carry[14]) );
  FA_152 sumI_14 ( .A(A[14]), .B(B[14]), .Ci(carry[14]), .S(res[14]), .Co(
        carry[15]) );
  FA_151 sumI_15 ( .A(A[15]), .B(B[15]), .Ci(carry[15]), .S(res[15]), .Co(
        carry[16]) );
  FA_150 sumTH ( .A(A[16]), .B(B[16]), .Ci(carry[16]), .S(res[16]), .Co(Co) );
endmodule


module FA_149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_MUL_WIDTH16_5 ( A, B, Ci, S, Partial, Co );
  input [16:0] A;
  input [16:0] B;
  output [16:0] S;
  output [1:0] Partial;
  input Ci;
  output Co;

  wire   [16:2] res;
  wire   [16:1] carry;
  assign S[14] = res[16];
  assign S[15] = res[16];
  assign S[16] = res[16];
  assign S[13] = res[15];
  assign S[12] = res[14];
  assign S[11] = res[13];
  assign S[10] = res[12];
  assign S[9] = res[11];
  assign S[8] = res[10];
  assign S[7] = res[9];
  assign S[6] = res[8];
  assign S[5] = res[7];
  assign S[4] = res[6];
  assign S[3] = res[5];
  assign S[2] = res[4];
  assign S[1] = res[3];
  assign S[0] = res[2];

  FA_149 sum0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(Partial[0]), .Co(carry[1]) );
  FA_148 sumI_1 ( .A(A[1]), .B(B[1]), .Ci(carry[1]), .S(Partial[1]), .Co(
        carry[2]) );
  FA_147 sumI_2 ( .A(A[2]), .B(B[2]), .Ci(carry[2]), .S(res[2]), .Co(carry[3])
         );
  FA_146 sumI_3 ( .A(A[3]), .B(B[3]), .Ci(carry[3]), .S(res[3]), .Co(carry[4])
         );
  FA_145 sumI_4 ( .A(A[4]), .B(B[4]), .Ci(carry[4]), .S(res[4]), .Co(carry[5])
         );
  FA_144 sumI_5 ( .A(A[5]), .B(B[5]), .Ci(carry[5]), .S(res[5]), .Co(carry[6])
         );
  FA_143 sumI_6 ( .A(A[6]), .B(B[6]), .Ci(carry[6]), .S(res[6]), .Co(carry[7])
         );
  FA_142 sumI_7 ( .A(A[7]), .B(B[7]), .Ci(carry[7]), .S(res[7]), .Co(carry[8])
         );
  FA_141 sumI_8 ( .A(A[8]), .B(B[8]), .Ci(carry[8]), .S(res[8]), .Co(carry[9])
         );
  FA_140 sumI_9 ( .A(A[9]), .B(B[9]), .Ci(carry[9]), .S(res[9]), .Co(carry[10]) );
  FA_139 sumI_10 ( .A(A[10]), .B(B[10]), .Ci(carry[10]), .S(res[10]), .Co(
        carry[11]) );
  FA_138 sumI_11 ( .A(A[11]), .B(B[11]), .Ci(carry[11]), .S(res[11]), .Co(
        carry[12]) );
  FA_137 sumI_12 ( .A(A[12]), .B(B[12]), .Ci(carry[12]), .S(res[12]), .Co(
        carry[13]) );
  FA_136 sumI_13 ( .A(A[13]), .B(B[13]), .Ci(carry[13]), .S(res[13]), .Co(
        carry[14]) );
  FA_135 sumI_14 ( .A(A[14]), .B(B[14]), .Ci(carry[14]), .S(res[14]), .Co(
        carry[15]) );
  FA_134 sumI_15 ( .A(A[15]), .B(B[15]), .Ci(carry[15]), .S(res[15]), .Co(
        carry[16]) );
  FA_133 sumTH ( .A(A[16]), .B(B[16]), .Ci(carry[16]), .S(res[16]), .Co(Co) );
endmodule


module FA_132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_MUL_WIDTH16_4 ( A, B, Ci, S, Partial, Co );
  input [16:0] A;
  input [16:0] B;
  output [16:0] S;
  output [1:0] Partial;
  input Ci;
  output Co;

  wire   [16:2] res;
  wire   [16:1] carry;
  assign S[14] = res[16];
  assign S[15] = res[16];
  assign S[16] = res[16];
  assign S[13] = res[15];
  assign S[12] = res[14];
  assign S[11] = res[13];
  assign S[10] = res[12];
  assign S[9] = res[11];
  assign S[8] = res[10];
  assign S[7] = res[9];
  assign S[6] = res[8];
  assign S[5] = res[7];
  assign S[4] = res[6];
  assign S[3] = res[5];
  assign S[2] = res[4];
  assign S[1] = res[3];
  assign S[0] = res[2];

  FA_132 sum0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(Partial[0]), .Co(carry[1]) );
  FA_131 sumI_1 ( .A(A[1]), .B(B[1]), .Ci(carry[1]), .S(Partial[1]), .Co(
        carry[2]) );
  FA_130 sumI_2 ( .A(A[2]), .B(B[2]), .Ci(carry[2]), .S(res[2]), .Co(carry[3])
         );
  FA_129 sumI_3 ( .A(A[3]), .B(B[3]), .Ci(carry[3]), .S(res[3]), .Co(carry[4])
         );
  FA_128 sumI_4 ( .A(A[4]), .B(B[4]), .Ci(carry[4]), .S(res[4]), .Co(carry[5])
         );
  FA_127 sumI_5 ( .A(A[5]), .B(B[5]), .Ci(carry[5]), .S(res[5]), .Co(carry[6])
         );
  FA_126 sumI_6 ( .A(A[6]), .B(B[6]), .Ci(carry[6]), .S(res[6]), .Co(carry[7])
         );
  FA_125 sumI_7 ( .A(A[7]), .B(B[7]), .Ci(carry[7]), .S(res[7]), .Co(carry[8])
         );
  FA_124 sumI_8 ( .A(A[8]), .B(B[8]), .Ci(carry[8]), .S(res[8]), .Co(carry[9])
         );
  FA_123 sumI_9 ( .A(A[9]), .B(B[9]), .Ci(carry[9]), .S(res[9]), .Co(carry[10]) );
  FA_122 sumI_10 ( .A(A[10]), .B(B[10]), .Ci(carry[10]), .S(res[10]), .Co(
        carry[11]) );
  FA_121 sumI_11 ( .A(A[11]), .B(B[11]), .Ci(carry[11]), .S(res[11]), .Co(
        carry[12]) );
  FA_120 sumI_12 ( .A(A[12]), .B(B[12]), .Ci(carry[12]), .S(res[12]), .Co(
        carry[13]) );
  FA_119 sumI_13 ( .A(A[13]), .B(B[13]), .Ci(carry[13]), .S(res[13]), .Co(
        carry[14]) );
  FA_118 sumI_14 ( .A(A[14]), .B(B[14]), .Ci(carry[14]), .S(res[14]), .Co(
        carry[15]) );
  FA_117 sumI_15 ( .A(A[15]), .B(B[15]), .Ci(carry[15]), .S(res[15]), .Co(
        carry[16]) );
  FA_116 sumTH ( .A(A[16]), .B(B[16]), .Ci(carry[16]), .S(res[16]), .Co(Co) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_MUL_WIDTH16_3 ( A, B, Ci, S, Partial, Co );
  input [16:0] A;
  input [16:0] B;
  output [16:0] S;
  output [1:0] Partial;
  input Ci;
  output Co;

  wire   [16:2] res;
  wire   [16:1] carry;
  assign S[14] = res[16];
  assign S[15] = res[16];
  assign S[16] = res[16];
  assign S[13] = res[15];
  assign S[12] = res[14];
  assign S[11] = res[13];
  assign S[10] = res[12];
  assign S[9] = res[11];
  assign S[8] = res[10];
  assign S[7] = res[9];
  assign S[6] = res[8];
  assign S[5] = res[7];
  assign S[4] = res[6];
  assign S[3] = res[5];
  assign S[2] = res[4];
  assign S[1] = res[3];
  assign S[0] = res[2];

  FA_115 sum0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(Partial[0]), .Co(carry[1]) );
  FA_114 sumI_1 ( .A(A[1]), .B(B[1]), .Ci(carry[1]), .S(Partial[1]), .Co(
        carry[2]) );
  FA_113 sumI_2 ( .A(A[2]), .B(B[2]), .Ci(carry[2]), .S(res[2]), .Co(carry[3])
         );
  FA_112 sumI_3 ( .A(A[3]), .B(B[3]), .Ci(carry[3]), .S(res[3]), .Co(carry[4])
         );
  FA_111 sumI_4 ( .A(A[4]), .B(B[4]), .Ci(carry[4]), .S(res[4]), .Co(carry[5])
         );
  FA_110 sumI_5 ( .A(A[5]), .B(B[5]), .Ci(carry[5]), .S(res[5]), .Co(carry[6])
         );
  FA_109 sumI_6 ( .A(A[6]), .B(B[6]), .Ci(carry[6]), .S(res[6]), .Co(carry[7])
         );
  FA_108 sumI_7 ( .A(A[7]), .B(B[7]), .Ci(carry[7]), .S(res[7]), .Co(carry[8])
         );
  FA_107 sumI_8 ( .A(A[8]), .B(B[8]), .Ci(carry[8]), .S(res[8]), .Co(carry[9])
         );
  FA_106 sumI_9 ( .A(A[9]), .B(B[9]), .Ci(carry[9]), .S(res[9]), .Co(carry[10]) );
  FA_105 sumI_10 ( .A(A[10]), .B(B[10]), .Ci(carry[10]), .S(res[10]), .Co(
        carry[11]) );
  FA_104 sumI_11 ( .A(A[11]), .B(B[11]), .Ci(carry[11]), .S(res[11]), .Co(
        carry[12]) );
  FA_103 sumI_12 ( .A(A[12]), .B(B[12]), .Ci(carry[12]), .S(res[12]), .Co(
        carry[13]) );
  FA_102 sumI_13 ( .A(A[13]), .B(B[13]), .Ci(carry[13]), .S(res[13]), .Co(
        carry[14]) );
  FA_101 sumI_14 ( .A(A[14]), .B(B[14]), .Ci(carry[14]), .S(res[14]), .Co(
        carry[15]) );
  FA_100 sumI_15 ( .A(A[15]), .B(B[15]), .Ci(carry[15]), .S(res[15]), .Co(
        carry[16]) );
  FA_99 sumTH ( .A(A[16]), .B(B[16]), .Ci(carry[16]), .S(res[16]), .Co(Co) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_MUL_WIDTH16_2 ( A, B, Ci, S, Partial, Co );
  input [16:0] A;
  input [16:0] B;
  output [16:0] S;
  output [1:0] Partial;
  input Ci;
  output Co;

  wire   [16:2] res;
  wire   [16:1] carry;
  assign S[14] = res[16];
  assign S[15] = res[16];
  assign S[16] = res[16];
  assign S[13] = res[15];
  assign S[12] = res[14];
  assign S[11] = res[13];
  assign S[10] = res[12];
  assign S[9] = res[11];
  assign S[8] = res[10];
  assign S[7] = res[9];
  assign S[6] = res[8];
  assign S[5] = res[7];
  assign S[4] = res[6];
  assign S[3] = res[5];
  assign S[2] = res[4];
  assign S[1] = res[3];
  assign S[0] = res[2];

  FA_98 sum0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(Partial[0]), .Co(carry[1]) );
  FA_97 sumI_1 ( .A(A[1]), .B(B[1]), .Ci(carry[1]), .S(Partial[1]), .Co(
        carry[2]) );
  FA_96 sumI_2 ( .A(A[2]), .B(B[2]), .Ci(carry[2]), .S(res[2]), .Co(carry[3])
         );
  FA_95 sumI_3 ( .A(A[3]), .B(B[3]), .Ci(carry[3]), .S(res[3]), .Co(carry[4])
         );
  FA_94 sumI_4 ( .A(A[4]), .B(B[4]), .Ci(carry[4]), .S(res[4]), .Co(carry[5])
         );
  FA_93 sumI_5 ( .A(A[5]), .B(B[5]), .Ci(carry[5]), .S(res[5]), .Co(carry[6])
         );
  FA_92 sumI_6 ( .A(A[6]), .B(B[6]), .Ci(carry[6]), .S(res[6]), .Co(carry[7])
         );
  FA_91 sumI_7 ( .A(A[7]), .B(B[7]), .Ci(carry[7]), .S(res[7]), .Co(carry[8])
         );
  FA_90 sumI_8 ( .A(A[8]), .B(B[8]), .Ci(carry[8]), .S(res[8]), .Co(carry[9])
         );
  FA_89 sumI_9 ( .A(A[9]), .B(B[9]), .Ci(carry[9]), .S(res[9]), .Co(carry[10])
         );
  FA_88 sumI_10 ( .A(A[10]), .B(B[10]), .Ci(carry[10]), .S(res[10]), .Co(
        carry[11]) );
  FA_87 sumI_11 ( .A(A[11]), .B(B[11]), .Ci(carry[11]), .S(res[11]), .Co(
        carry[12]) );
  FA_86 sumI_12 ( .A(A[12]), .B(B[12]), .Ci(carry[12]), .S(res[12]), .Co(
        carry[13]) );
  FA_85 sumI_13 ( .A(A[13]), .B(B[13]), .Ci(carry[13]), .S(res[13]), .Co(
        carry[14]) );
  FA_84 sumI_14 ( .A(A[14]), .B(B[14]), .Ci(carry[14]), .S(res[14]), .Co(
        carry[15]) );
  FA_83 sumI_15 ( .A(A[15]), .B(B[15]), .Ci(carry[15]), .S(res[15]), .Co(
        carry[16]) );
  FA_82 sumTH ( .A(A[16]), .B(B[16]), .Ci(carry[16]), .S(res[16]), .Co(Co) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n17), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n17) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n17), .B2(Ci), .ZN(n18) );
endmodule


module RCA_MUL_WIDTH16_1 ( A, B, Ci, S, Partial, Co );
  input [16:0] A;
  input [16:0] B;
  output [16:0] S;
  output [1:0] Partial;
  input Ci;
  output Co;

  wire   [16:2] res;
  wire   [16:1] carry;
  assign S[14] = res[16];
  assign S[15] = res[16];
  assign S[16] = res[16];
  assign S[13] = res[15];
  assign S[12] = res[14];
  assign S[11] = res[13];
  assign S[10] = res[12];
  assign S[9] = res[11];
  assign S[8] = res[10];
  assign S[7] = res[9];
  assign S[6] = res[8];
  assign S[5] = res[7];
  assign S[4] = res[6];
  assign S[3] = res[5];
  assign S[2] = res[4];
  assign S[1] = res[3];
  assign S[0] = res[2];

  FA_81 sum0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(Partial[0]), .Co(carry[1]) );
  FA_80 sumI_1 ( .A(A[1]), .B(B[1]), .Ci(carry[1]), .S(Partial[1]), .Co(
        carry[2]) );
  FA_79 sumI_2 ( .A(A[2]), .B(B[2]), .Ci(carry[2]), .S(res[2]), .Co(carry[3])
         );
  FA_78 sumI_3 ( .A(A[3]), .B(B[3]), .Ci(carry[3]), .S(res[3]), .Co(carry[4])
         );
  FA_77 sumI_4 ( .A(A[4]), .B(B[4]), .Ci(carry[4]), .S(res[4]), .Co(carry[5])
         );
  FA_76 sumI_5 ( .A(A[5]), .B(B[5]), .Ci(carry[5]), .S(res[5]), .Co(carry[6])
         );
  FA_75 sumI_6 ( .A(A[6]), .B(B[6]), .Ci(carry[6]), .S(res[6]), .Co(carry[7])
         );
  FA_74 sumI_7 ( .A(A[7]), .B(B[7]), .Ci(carry[7]), .S(res[7]), .Co(carry[8])
         );
  FA_73 sumI_8 ( .A(A[8]), .B(B[8]), .Ci(carry[8]), .S(res[8]), .Co(carry[9])
         );
  FA_72 sumI_9 ( .A(A[9]), .B(B[9]), .Ci(carry[9]), .S(res[9]), .Co(carry[10])
         );
  FA_71 sumI_10 ( .A(A[10]), .B(B[10]), .Ci(carry[10]), .S(res[10]), .Co(
        carry[11]) );
  FA_70 sumI_11 ( .A(A[11]), .B(B[11]), .Ci(carry[11]), .S(res[11]), .Co(
        carry[12]) );
  FA_69 sumI_12 ( .A(A[12]), .B(B[12]), .Ci(carry[12]), .S(res[12]), .Co(
        carry[13]) );
  FA_68 sumI_13 ( .A(A[13]), .B(B[13]), .Ci(carry[13]), .S(res[13]), .Co(
        carry[14]) );
  FA_67 sumI_14 ( .A(A[14]), .B(B[14]), .Ci(carry[14]), .S(res[14]), .Co(
        carry[15]) );
  FA_66 sumI_15 ( .A(A[15]), .B(B[15]), .Ci(carry[15]), .S(res[15]), .Co(
        carry[16]) );
  FA_65 sumTH ( .A(A[16]), .B(B[16]), .Ci(carry[16]), .S(res[16]), .Co(Co) );
endmodule


module MULTIPLIER_WIDTH16 ( A, B, P );
  input [15:0] A;
  input [15:0] B;
  output [31:0] P;
  wire   \outEnc[7][16] , \outEnc[7][15] , \outEnc[7][14] , \outEnc[7][13] ,
         \outEnc[7][12] , \outEnc[7][11] , \outEnc[7][10] , \outEnc[7][9] ,
         \outEnc[7][8] , \outEnc[7][7] , \outEnc[7][6] , \outEnc[7][5] ,
         \outEnc[7][4] , \outEnc[7][3] , \outEnc[7][2] , \outEnc[7][1] ,
         \outEnc[7][0] , \outEnc[6][16] , \outEnc[6][15] , \outEnc[6][14] ,
         \outEnc[6][13] , \outEnc[6][12] , \outEnc[6][11] , \outEnc[6][10] ,
         \outEnc[6][9] , \outEnc[6][8] , \outEnc[6][7] , \outEnc[6][6] ,
         \outEnc[6][5] , \outEnc[6][4] , \outEnc[6][3] , \outEnc[6][2] ,
         \outEnc[6][1] , \outEnc[6][0] , \outEnc[5][16] , \outEnc[5][15] ,
         \outEnc[5][14] , \outEnc[5][13] , \outEnc[5][12] , \outEnc[5][11] ,
         \outEnc[5][10] , \outEnc[5][9] , \outEnc[5][8] , \outEnc[5][7] ,
         \outEnc[5][6] , \outEnc[5][5] , \outEnc[5][4] , \outEnc[5][3] ,
         \outEnc[5][2] , \outEnc[5][1] , \outEnc[5][0] , \outEnc[4][16] ,
         \outEnc[4][15] , \outEnc[4][14] , \outEnc[4][13] , \outEnc[4][12] ,
         \outEnc[4][11] , \outEnc[4][10] , \outEnc[4][9] , \outEnc[4][8] ,
         \outEnc[4][7] , \outEnc[4][6] , \outEnc[4][5] , \outEnc[4][4] ,
         \outEnc[4][3] , \outEnc[4][2] , \outEnc[4][1] , \outEnc[4][0] ,
         \outEnc[3][16] , \outEnc[3][15] , \outEnc[3][14] , \outEnc[3][13] ,
         \outEnc[3][12] , \outEnc[3][11] , \outEnc[3][10] , \outEnc[3][9] ,
         \outEnc[3][8] , \outEnc[3][7] , \outEnc[3][6] , \outEnc[3][5] ,
         \outEnc[3][4] , \outEnc[3][3] , \outEnc[3][2] , \outEnc[3][1] ,
         \outEnc[3][0] , \outEnc[2][16] , \outEnc[2][15] , \outEnc[2][14] ,
         \outEnc[2][13] , \outEnc[2][12] , \outEnc[2][11] , \outEnc[2][10] ,
         \outEnc[2][9] , \outEnc[2][8] , \outEnc[2][7] , \outEnc[2][6] ,
         \outEnc[2][5] , \outEnc[2][4] , \outEnc[2][3] , \outEnc[2][2] ,
         \outEnc[2][1] , \outEnc[2][0] , \outEnc[1][16] , \outEnc[1][15] ,
         \outEnc[1][14] , \outEnc[1][13] , \outEnc[1][12] , \outEnc[1][11] ,
         \outEnc[1][10] , \outEnc[1][9] , \outEnc[1][8] , \outEnc[1][7] ,
         \outEnc[1][6] , \outEnc[1][5] , \outEnc[1][4] , \outEnc[1][3] ,
         \outEnc[1][2] , \outEnc[1][1] , \outEnc[1][0] , \outEnc[0][16] ,
         \outEnc[0][15] , \outEnc[0][14] , \outEnc[0][13] , \outEnc[0][12] ,
         \outEnc[0][11] , \outEnc[0][10] , \outEnc[0][9] , \outEnc[0][8] ,
         \outEnc[0][7] , \outEnc[0][6] , \outEnc[0][5] , \outEnc[0][4] ,
         \outEnc[0][3] , \outEnc[0][2] , \outEnc[0][1] , \outEnc[0][0] ,
         \outSum[6][16] , \outSum[6][15] , \outSum[6][14] , \outSum[6][13] ,
         \outSum[6][12] , \outSum[6][11] , \outSum[6][10] , \outSum[6][9] ,
         \outSum[6][8] , \outSum[6][7] , \outSum[6][6] , \outSum[6][5] ,
         \outSum[6][4] , \outSum[6][3] , \outSum[6][2] , \outSum[6][1] ,
         \outSum[6][0] , \outSum[5][16] , \outSum[5][15] , \outSum[5][14] ,
         \outSum[5][13] , \outSum[5][12] , \outSum[5][11] , \outSum[5][10] ,
         \outSum[5][9] , \outSum[5][8] , \outSum[5][7] , \outSum[5][6] ,
         \outSum[5][5] , \outSum[5][4] , \outSum[5][3] , \outSum[5][2] ,
         \outSum[5][1] , \outSum[5][0] , \outSum[4][16] , \outSum[4][15] ,
         \outSum[4][14] , \outSum[4][13] , \outSum[4][12] , \outSum[4][11] ,
         \outSum[4][10] , \outSum[4][9] , \outSum[4][8] , \outSum[4][7] ,
         \outSum[4][6] , \outSum[4][5] , \outSum[4][4] , \outSum[4][3] ,
         \outSum[4][2] , \outSum[4][1] , \outSum[4][0] , \outSum[3][16] ,
         \outSum[3][15] , \outSum[3][14] , \outSum[3][13] , \outSum[3][12] ,
         \outSum[3][11] , \outSum[3][10] , \outSum[3][9] , \outSum[3][8] ,
         \outSum[3][7] , \outSum[3][6] , \outSum[3][5] , \outSum[3][4] ,
         \outSum[3][3] , \outSum[3][2] , \outSum[3][1] , \outSum[3][0] ,
         \outSum[2][16] , \outSum[2][15] , \outSum[2][14] , \outSum[2][13] ,
         \outSum[2][12] , \outSum[2][11] , \outSum[2][10] , \outSum[2][9] ,
         \outSum[2][8] , \outSum[2][7] , \outSum[2][6] , \outSum[2][5] ,
         \outSum[2][4] , \outSum[2][3] , \outSum[2][2] , \outSum[2][1] ,
         \outSum[2][0] , \outSum[1][16] , \outSum[1][15] , \outSum[1][14] ,
         \outSum[1][13] , \outSum[1][12] , \outSum[1][11] , \outSum[1][10] ,
         \outSum[1][9] , \outSum[1][8] , \outSum[1][7] , \outSum[1][6] ,
         \outSum[1][5] , \outSum[1][4] , \outSum[1][3] , \outSum[1][2] ,
         \outSum[1][1] , \outSum[1][0] , \outSum[0][16] , \outSum[0][15] ,
         \outSum[0][14] , \outSum[0][13] , \outSum[0][12] , \outSum[0][11] ,
         \outSum[0][10] , \outSum[0][9] , \outSum[0][8] , \outSum[0][7] ,
         \outSum[0][6] , \outSum[0][5] , \outSum[0][4] , \outSum[0][3] ,
         \outSum[0][2] , \outSum[0][1] , \outSum[0][0] , n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133;
  wire   SYNOPSYS_UNCONNECTED__0;

  BOOTH_ENCODER_WIDTH16_0 enc0 ( .A({n133, n132, n129, n128, n127, A[10], n124, 
        n123, n120, n117, n115, n112, n109, n107, A[1:0]}), .b({B[1:0], 1'b0}), 
        .vp({\outEnc[0][16] , \outEnc[0][15] , \outEnc[0][14] , 
        \outEnc[0][13] , \outEnc[0][12] , \outEnc[0][11] , \outEnc[0][10] , 
        \outEnc[0][9] , \outEnc[0][8] , \outEnc[0][7] , \outEnc[0][6] , 
        \outEnc[0][5] , \outEnc[0][4] , \outEnc[0][3] , \outEnc[0][2] , 
        \outEnc[0][1] , \outEnc[0][0] }) );
  BOOTH_ENCODER_WIDTH16_7 ENCi_0 ( .A({n133, n132, n129, n128, n127, A[10], 
        n124, n123, n120, n117, n115, n112, n109, n107, A[1:0]}), .b(B[3:1]), 
        .vp({\outEnc[1][16] , \outEnc[1][15] , \outEnc[1][14] , 
        \outEnc[1][13] , \outEnc[1][12] , \outEnc[1][11] , \outEnc[1][10] , 
        \outEnc[1][9] , \outEnc[1][8] , \outEnc[1][7] , \outEnc[1][6] , 
        \outEnc[1][5] , \outEnc[1][4] , \outEnc[1][3] , \outEnc[1][2] , 
        \outEnc[1][1] , \outEnc[1][0] }) );
  BOOTH_ENCODER_WIDTH16_6 ENCi_1 ( .A({n133, n131, n129, n128, n126, A[10], 
        n124, n122, n119, n117, n114, n111, n109, n106, A[1:0]}), .b(B[5:3]), 
        .vp({\outEnc[2][16] , \outEnc[2][15] , \outEnc[2][14] , 
        \outEnc[2][13] , \outEnc[2][12] , \outEnc[2][11] , \outEnc[2][10] , 
        \outEnc[2][9] , \outEnc[2][8] , \outEnc[2][7] , \outEnc[2][6] , 
        \outEnc[2][5] , \outEnc[2][4] , \outEnc[2][3] , \outEnc[2][2] , 
        \outEnc[2][1] , \outEnc[2][0] }) );
  BOOTH_ENCODER_WIDTH16_5 ENCi_2 ( .A({n133, n131, n129, n128, n126, A[10], 
        n124, n122, n119, n117, n114, n111, n109, n106, A[1:0]}), .b(B[7:5]), 
        .vp({\outEnc[3][16] , \outEnc[3][15] , \outEnc[3][14] , 
        \outEnc[3][13] , \outEnc[3][12] , \outEnc[3][11] , \outEnc[3][10] , 
        \outEnc[3][9] , \outEnc[3][8] , \outEnc[3][7] , \outEnc[3][6] , 
        \outEnc[3][5] , \outEnc[3][4] , \outEnc[3][3] , \outEnc[3][2] , 
        \outEnc[3][1] , \outEnc[3][0] }) );
  BOOTH_ENCODER_WIDTH16_4 ENCi_3 ( .A({n133, n130, n129, n128, n125, A[10], 
        n124, n121, n118, n116, n113, n110, n108, n105, A[1:0]}), .b(B[9:7]), 
        .vp({\outEnc[4][16] , \outEnc[4][15] , \outEnc[4][14] , 
        \outEnc[4][13] , \outEnc[4][12] , \outEnc[4][11] , \outEnc[4][10] , 
        \outEnc[4][9] , \outEnc[4][8] , \outEnc[4][7] , \outEnc[4][6] , 
        \outEnc[4][5] , \outEnc[4][4] , \outEnc[4][3] , \outEnc[4][2] , 
        \outEnc[4][1] , \outEnc[4][0] }) );
  BOOTH_ENCODER_WIDTH16_3 ENCi_4 ( .A({n133, n130, n129, n128, n125, A[10], 
        n124, n121, n118, n116, n113, n110, n108, n105, A[1:0]}), .b(B[11:9]), 
        .vp({\outEnc[5][16] , \outEnc[5][15] , \outEnc[5][14] , 
        \outEnc[5][13] , \outEnc[5][12] , \outEnc[5][11] , \outEnc[5][10] , 
        \outEnc[5][9] , \outEnc[5][8] , \outEnc[5][7] , \outEnc[5][6] , 
        \outEnc[5][5] , \outEnc[5][4] , \outEnc[5][3] , \outEnc[5][2] , 
        \outEnc[5][1] , \outEnc[5][0] }) );
  BOOTH_ENCODER_WIDTH16_2 ENCi_5 ( .A({n133, n130, n129, n128, n125, A[10], 
        n124, n121, n118, n116, n113, n110, n108, n105, A[1:0]}), .b(B[13:11]), 
        .vp({\outEnc[6][16] , \outEnc[6][15] , \outEnc[6][14] , 
        \outEnc[6][13] , \outEnc[6][12] , \outEnc[6][11] , \outEnc[6][10] , 
        \outEnc[6][9] , \outEnc[6][8] , \outEnc[6][7] , \outEnc[6][6] , 
        \outEnc[6][5] , \outEnc[6][4] , \outEnc[6][3] , \outEnc[6][2] , 
        \outEnc[6][1] , \outEnc[6][0] }) );
  BOOTH_ENCODER_WIDTH16_1 ENCi_6 ( .A({n133, n131, n129, n128, n126, A[10], 
        n124, n122, n119, n116, n114, n111, n108, n106, A[1:0]}), .b(B[15:13]), 
        .vp({\outEnc[7][16] , \outEnc[7][15] , \outEnc[7][14] , 
        \outEnc[7][13] , \outEnc[7][12] , \outEnc[7][11] , \outEnc[7][10] , 
        \outEnc[7][9] , \outEnc[7][8] , \outEnc[7][7] , \outEnc[7][6] , 
        \outEnc[7][5] , \outEnc[7][4] , \outEnc[7][3] , \outEnc[7][2] , 
        \outEnc[7][1] , \outEnc[7][0] }) );
  RCA_MUL_WIDTH16_0 rca0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \outEnc[0][16] , \outEnc[0][15] , \outEnc[0][14] , \outEnc[0][13] , 
        \outEnc[0][12] , \outEnc[0][11] , \outEnc[0][10] , \outEnc[0][9] , 
        \outEnc[0][8] , \outEnc[0][7] , \outEnc[0][6] , \outEnc[0][5] , 
        \outEnc[0][4] , \outEnc[0][3] , \outEnc[0][2] , \outEnc[0][1] , 
        \outEnc[0][0] }), .Ci(1'b0), .S({\outSum[0][16] , \outSum[0][15] , 
        \outSum[0][14] , \outSum[0][13] , \outSum[0][12] , \outSum[0][11] , 
        \outSum[0][10] , \outSum[0][9] , \outSum[0][8] , \outSum[0][7] , 
        \outSum[0][6] , \outSum[0][5] , \outSum[0][4] , \outSum[0][3] , 
        \outSum[0][2] , \outSum[0][1] , \outSum[0][0] }), .Partial(P[1:0]) );
  RCA_MUL_WIDTH16_7 rcai_0 ( .A({\outSum[0][16] , \outSum[0][15] , 
        \outSum[0][14] , \outSum[0][13] , \outSum[0][12] , \outSum[0][11] , 
        \outSum[0][10] , \outSum[0][9] , \outSum[0][8] , \outSum[0][7] , 
        \outSum[0][6] , \outSum[0][5] , \outSum[0][4] , \outSum[0][3] , 
        \outSum[0][2] , \outSum[0][1] , \outSum[0][0] }), .B({\outEnc[1][16] , 
        \outEnc[1][15] , \outEnc[1][14] , \outEnc[1][13] , \outEnc[1][12] , 
        \outEnc[1][11] , \outEnc[1][10] , \outEnc[1][9] , \outEnc[1][8] , 
        \outEnc[1][7] , \outEnc[1][6] , \outEnc[1][5] , \outEnc[1][4] , 
        \outEnc[1][3] , \outEnc[1][2] , \outEnc[1][1] , \outEnc[1][0] }), .Ci(
        1'b0), .S({\outSum[1][16] , \outSum[1][15] , \outSum[1][14] , 
        \outSum[1][13] , \outSum[1][12] , \outSum[1][11] , \outSum[1][10] , 
        \outSum[1][9] , \outSum[1][8] , \outSum[1][7] , \outSum[1][6] , 
        \outSum[1][5] , \outSum[1][4] , \outSum[1][3] , \outSum[1][2] , 
        \outSum[1][1] , \outSum[1][0] }), .Partial(P[3:2]) );
  RCA_MUL_WIDTH16_6 rcai_1 ( .A({\outSum[1][16] , \outSum[1][15] , 
        \outSum[1][14] , \outSum[1][13] , \outSum[1][12] , \outSum[1][11] , 
        \outSum[1][10] , \outSum[1][9] , \outSum[1][8] , \outSum[1][7] , 
        \outSum[1][6] , \outSum[1][5] , \outSum[1][4] , \outSum[1][3] , 
        \outSum[1][2] , \outSum[1][1] , \outSum[1][0] }), .B({\outEnc[2][16] , 
        \outEnc[2][15] , \outEnc[2][14] , \outEnc[2][13] , \outEnc[2][12] , 
        \outEnc[2][11] , \outEnc[2][10] , \outEnc[2][9] , \outEnc[2][8] , 
        \outEnc[2][7] , \outEnc[2][6] , \outEnc[2][5] , \outEnc[2][4] , 
        \outEnc[2][3] , \outEnc[2][2] , \outEnc[2][1] , \outEnc[2][0] }), .Ci(
        1'b0), .S({\outSum[2][16] , \outSum[2][15] , \outSum[2][14] , 
        \outSum[2][13] , \outSum[2][12] , \outSum[2][11] , \outSum[2][10] , 
        \outSum[2][9] , \outSum[2][8] , \outSum[2][7] , \outSum[2][6] , 
        \outSum[2][5] , \outSum[2][4] , \outSum[2][3] , \outSum[2][2] , 
        \outSum[2][1] , \outSum[2][0] }), .Partial(P[5:4]) );
  RCA_MUL_WIDTH16_5 rcai_2 ( .A({\outSum[2][16] , \outSum[2][15] , 
        \outSum[2][14] , \outSum[2][13] , \outSum[2][12] , \outSum[2][11] , 
        \outSum[2][10] , \outSum[2][9] , \outSum[2][8] , \outSum[2][7] , 
        \outSum[2][6] , \outSum[2][5] , \outSum[2][4] , \outSum[2][3] , 
        \outSum[2][2] , \outSum[2][1] , \outSum[2][0] }), .B({\outEnc[3][16] , 
        \outEnc[3][15] , \outEnc[3][14] , \outEnc[3][13] , \outEnc[3][12] , 
        \outEnc[3][11] , \outEnc[3][10] , \outEnc[3][9] , \outEnc[3][8] , 
        \outEnc[3][7] , \outEnc[3][6] , \outEnc[3][5] , \outEnc[3][4] , 
        \outEnc[3][3] , \outEnc[3][2] , \outEnc[3][1] , \outEnc[3][0] }), .Ci(
        1'b0), .S({\outSum[3][16] , \outSum[3][15] , \outSum[3][14] , 
        \outSum[3][13] , \outSum[3][12] , \outSum[3][11] , \outSum[3][10] , 
        \outSum[3][9] , \outSum[3][8] , \outSum[3][7] , \outSum[3][6] , 
        \outSum[3][5] , \outSum[3][4] , \outSum[3][3] , \outSum[3][2] , 
        \outSum[3][1] , \outSum[3][0] }), .Partial(P[7:6]) );
  RCA_MUL_WIDTH16_4 rcai_3 ( .A({\outSum[3][16] , \outSum[3][15] , 
        \outSum[3][14] , \outSum[3][13] , \outSum[3][12] , \outSum[3][11] , 
        \outSum[3][10] , \outSum[3][9] , \outSum[3][8] , \outSum[3][7] , 
        \outSum[3][6] , \outSum[3][5] , \outSum[3][4] , \outSum[3][3] , 
        \outSum[3][2] , \outSum[3][1] , \outSum[3][0] }), .B({\outEnc[4][16] , 
        \outEnc[4][15] , \outEnc[4][14] , \outEnc[4][13] , \outEnc[4][12] , 
        \outEnc[4][11] , \outEnc[4][10] , \outEnc[4][9] , \outEnc[4][8] , 
        \outEnc[4][7] , \outEnc[4][6] , \outEnc[4][5] , \outEnc[4][4] , 
        \outEnc[4][3] , \outEnc[4][2] , \outEnc[4][1] , \outEnc[4][0] }), .Ci(
        1'b0), .S({\outSum[4][16] , \outSum[4][15] , \outSum[4][14] , 
        \outSum[4][13] , \outSum[4][12] , \outSum[4][11] , \outSum[4][10] , 
        \outSum[4][9] , \outSum[4][8] , \outSum[4][7] , \outSum[4][6] , 
        \outSum[4][5] , \outSum[4][4] , \outSum[4][3] , \outSum[4][2] , 
        \outSum[4][1] , \outSum[4][0] }), .Partial(P[9:8]) );
  RCA_MUL_WIDTH16_3 rcai_4 ( .A({\outSum[4][16] , \outSum[4][15] , 
        \outSum[4][14] , \outSum[4][13] , \outSum[4][12] , \outSum[4][11] , 
        \outSum[4][10] , \outSum[4][9] , \outSum[4][8] , \outSum[4][7] , 
        \outSum[4][6] , \outSum[4][5] , \outSum[4][4] , \outSum[4][3] , 
        \outSum[4][2] , \outSum[4][1] , \outSum[4][0] }), .B({\outEnc[5][16] , 
        \outEnc[5][15] , \outEnc[5][14] , \outEnc[5][13] , \outEnc[5][12] , 
        \outEnc[5][11] , \outEnc[5][10] , \outEnc[5][9] , \outEnc[5][8] , 
        \outEnc[5][7] , \outEnc[5][6] , \outEnc[5][5] , \outEnc[5][4] , 
        \outEnc[5][3] , \outEnc[5][2] , \outEnc[5][1] , \outEnc[5][0] }), .Ci(
        1'b0), .S({\outSum[5][16] , \outSum[5][15] , \outSum[5][14] , 
        \outSum[5][13] , \outSum[5][12] , \outSum[5][11] , \outSum[5][10] , 
        \outSum[5][9] , \outSum[5][8] , \outSum[5][7] , \outSum[5][6] , 
        \outSum[5][5] , \outSum[5][4] , \outSum[5][3] , \outSum[5][2] , 
        \outSum[5][1] , \outSum[5][0] }), .Partial(P[11:10]) );
  RCA_MUL_WIDTH16_2 rcai_5 ( .A({\outSum[5][16] , \outSum[5][15] , 
        \outSum[5][14] , \outSum[5][13] , \outSum[5][12] , \outSum[5][11] , 
        \outSum[5][10] , \outSum[5][9] , \outSum[5][8] , \outSum[5][7] , 
        \outSum[5][6] , \outSum[5][5] , \outSum[5][4] , \outSum[5][3] , 
        \outSum[5][2] , \outSum[5][1] , \outSum[5][0] }), .B({\outEnc[6][16] , 
        \outEnc[6][15] , \outEnc[6][14] , \outEnc[6][13] , \outEnc[6][12] , 
        \outEnc[6][11] , \outEnc[6][10] , \outEnc[6][9] , \outEnc[6][8] , 
        \outEnc[6][7] , \outEnc[6][6] , \outEnc[6][5] , \outEnc[6][4] , 
        \outEnc[6][3] , \outEnc[6][2] , \outEnc[6][1] , \outEnc[6][0] }), .Ci(
        1'b0), .S({\outSum[6][16] , \outSum[6][15] , \outSum[6][14] , 
        \outSum[6][13] , \outSum[6][12] , \outSum[6][11] , \outSum[6][10] , 
        \outSum[6][9] , \outSum[6][8] , \outSum[6][7] , \outSum[6][6] , 
        \outSum[6][5] , \outSum[6][4] , \outSum[6][3] , \outSum[6][2] , 
        \outSum[6][1] , \outSum[6][0] }), .Partial(P[13:12]) );
  RCA_MUL_WIDTH16_1 rcai_6 ( .A({\outSum[6][16] , \outSum[6][15] , 
        \outSum[6][14] , \outSum[6][13] , \outSum[6][12] , \outSum[6][11] , 
        \outSum[6][10] , \outSum[6][9] , \outSum[6][8] , \outSum[6][7] , 
        \outSum[6][6] , \outSum[6][5] , \outSum[6][4] , \outSum[6][3] , 
        \outSum[6][2] , \outSum[6][1] , \outSum[6][0] }), .B({\outEnc[7][16] , 
        \outEnc[7][15] , \outEnc[7][14] , \outEnc[7][13] , \outEnc[7][12] , 
        \outEnc[7][11] , \outEnc[7][10] , \outEnc[7][9] , \outEnc[7][8] , 
        \outEnc[7][7] , \outEnc[7][6] , \outEnc[7][5] , \outEnc[7][4] , 
        \outEnc[7][3] , \outEnc[7][2] , \outEnc[7][1] , \outEnc[7][0] }), .Ci(
        1'b0), .S({SYNOPSYS_UNCONNECTED__0, P[31:16]}), .Partial(P[15:14]) );
  BUF_X1 U2 ( .A(A[6]), .Z(n117) );
  BUF_X1 U3 ( .A(A[3]), .Z(n109) );
  BUF_X1 U4 ( .A(A[3]), .Z(n108) );
  BUF_X1 U5 ( .A(A[6]), .Z(n116) );
  BUF_X1 U6 ( .A(A[12]), .Z(n128) );
  BUF_X1 U7 ( .A(A[13]), .Z(n129) );
  BUF_X2 U8 ( .A(A[15]), .Z(n133) );
  BUF_X2 U9 ( .A(A[9]), .Z(n124) );
  CLKBUF_X1 U10 ( .A(A[2]), .Z(n105) );
  CLKBUF_X1 U11 ( .A(A[2]), .Z(n106) );
  CLKBUF_X1 U12 ( .A(A[2]), .Z(n107) );
  CLKBUF_X1 U13 ( .A(A[4]), .Z(n110) );
  CLKBUF_X1 U14 ( .A(A[4]), .Z(n111) );
  CLKBUF_X1 U15 ( .A(A[4]), .Z(n112) );
  CLKBUF_X1 U16 ( .A(A[5]), .Z(n113) );
  CLKBUF_X1 U17 ( .A(A[5]), .Z(n114) );
  CLKBUF_X1 U18 ( .A(A[5]), .Z(n115) );
  CLKBUF_X1 U19 ( .A(A[7]), .Z(n118) );
  CLKBUF_X1 U20 ( .A(A[7]), .Z(n119) );
  CLKBUF_X1 U21 ( .A(A[7]), .Z(n120) );
  CLKBUF_X1 U22 ( .A(A[8]), .Z(n121) );
  CLKBUF_X1 U23 ( .A(A[8]), .Z(n122) );
  CLKBUF_X1 U24 ( .A(A[8]), .Z(n123) );
  CLKBUF_X1 U25 ( .A(A[11]), .Z(n125) );
  CLKBUF_X1 U26 ( .A(A[11]), .Z(n126) );
  CLKBUF_X1 U27 ( .A(A[11]), .Z(n127) );
  CLKBUF_X1 U28 ( .A(A[14]), .Z(n130) );
  CLKBUF_X1 U29 ( .A(A[14]), .Z(n131) );
  CLKBUF_X1 U30 ( .A(A[14]), .Z(n132) );
endmodule


module ALU_WIDTH32_RADIX4 ( A, B, .OP({\OP[4] , \OP[3] , \OP[2] , \OP[1] , 
        \OP[0] }), Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input \OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] ;
  wire   s_Co, s_SIGN, s_C, s_ADD_SUB, N20, N22, N24, N25, N27, s_LE, s_NE,
         s_Z, n114, n3, n110, n112, n115, n109, n206, n207, n103, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n104, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346;
  wire   [4:0] OP;
  wire   [31:0] s_A_ADDER;
  wire   [31:0] S_B_ADDER;
  wire   [31:0] s_A_LOGIC;
  wire   [31:0] S_B_LOGIC;
  wire   [3:0] s_LOGIC;
  wire   [31:0] s_A_SHIFT;
  wire   [31:0] S_B_SHIFT;
  wire   [1:0] s_SHIFT;
  wire   [15:0] s_A_MULT;
  wire   [15:0] S_B_MULT;
  wire   [15:0] S_B_LHI;
  wire   [31:0] s_OUT;
  wire   [31:0] s_LOG;
  wire   [31:0] s_SHI;
  wire   [31:0] s_MULT;
  wire   SYNOPSYS_UNCONNECTED__0;

  DLH_X1 s_SIGN_reg ( .G(n104), .D(N27), .Q(s_SIGN) );
  DLH_X1 \s_A_ADDER_reg[31]  ( .G(n325), .D(A[31]), .Q(s_A_ADDER[31]) );
  DLH_X1 \s_A_ADDER_reg[30]  ( .G(n327), .D(A[30]), .Q(s_A_ADDER[30]) );
  DLH_X1 \s_A_ADDER_reg[29]  ( .G(n327), .D(A[29]), .Q(s_A_ADDER[29]) );
  DLH_X1 \s_A_ADDER_reg[28]  ( .G(n327), .D(A[28]), .Q(s_A_ADDER[28]) );
  DLH_X1 \s_A_ADDER_reg[27]  ( .G(n325), .D(A[27]), .Q(s_A_ADDER[27]) );
  DLH_X1 \s_A_ADDER_reg[26]  ( .G(n328), .D(A[26]), .Q(s_A_ADDER[26]) );
  DLH_X1 \s_A_ADDER_reg[25]  ( .G(n328), .D(A[25]), .Q(s_A_ADDER[25]) );
  DLH_X1 \s_A_ADDER_reg[24]  ( .G(n327), .D(A[24]), .Q(s_A_ADDER[24]) );
  DLH_X1 \s_A_ADDER_reg[23]  ( .G(n331), .D(A[23]), .Q(s_A_ADDER[23]) );
  DLH_X1 \s_A_ADDER_reg[22]  ( .G(n325), .D(A[22]), .Q(s_A_ADDER[22]) );
  DLH_X1 \s_A_ADDER_reg[21]  ( .G(n327), .D(A[21]), .Q(s_A_ADDER[21]) );
  DLH_X1 \s_A_ADDER_reg[20]  ( .G(n328), .D(A[20]), .Q(s_A_ADDER[20]) );
  DLH_X1 \s_A_ADDER_reg[19]  ( .G(n325), .D(A[19]), .Q(s_A_ADDER[19]) );
  DLH_X1 \s_A_ADDER_reg[18]  ( .G(n325), .D(A[18]), .Q(s_A_ADDER[18]) );
  DLH_X1 \s_A_ADDER_reg[17]  ( .G(n327), .D(A[17]), .Q(s_A_ADDER[17]) );
  DLH_X1 \s_A_ADDER_reg[16]  ( .G(n326), .D(A[16]), .Q(s_A_ADDER[16]) );
  DLH_X1 \s_A_ADDER_reg[15]  ( .G(n331), .D(A[15]), .Q(s_A_ADDER[15]) );
  DLH_X1 \s_A_ADDER_reg[14]  ( .G(n326), .D(A[14]), .Q(s_A_ADDER[14]) );
  DLH_X1 \s_A_ADDER_reg[13]  ( .G(n326), .D(A[13]), .Q(s_A_ADDER[13]) );
  DLH_X1 \s_A_ADDER_reg[12]  ( .G(n326), .D(A[12]), .Q(s_A_ADDER[12]) );
  DLH_X1 \s_A_ADDER_reg[11]  ( .G(n330), .D(A[11]), .Q(s_A_ADDER[11]) );
  DLH_X1 \s_A_ADDER_reg[10]  ( .G(n331), .D(A[10]), .Q(s_A_ADDER[10]) );
  DLH_X1 \s_A_ADDER_reg[9]  ( .G(n325), .D(A[9]), .Q(s_A_ADDER[9]) );
  DLH_X1 \s_A_ADDER_reg[8]  ( .G(n325), .D(A[8]), .Q(s_A_ADDER[8]) );
  DLH_X1 \s_A_ADDER_reg[7]  ( .G(n330), .D(A[7]), .Q(s_A_ADDER[7]) );
  DLH_X1 \s_A_ADDER_reg[6]  ( .G(n326), .D(A[6]), .Q(s_A_ADDER[6]) );
  DLH_X1 \s_A_ADDER_reg[5]  ( .G(n328), .D(A[5]), .Q(s_A_ADDER[5]) );
  DLH_X1 \s_A_ADDER_reg[4]  ( .G(n325), .D(A[4]), .Q(s_A_ADDER[4]) );
  DLH_X1 \s_A_ADDER_reg[3]  ( .G(n331), .D(A[3]), .Q(s_A_ADDER[3]) );
  DLH_X1 \s_A_ADDER_reg[2]  ( .G(n326), .D(A[2]), .Q(s_A_ADDER[2]) );
  DLH_X1 \s_A_ADDER_reg[1]  ( .G(n326), .D(A[1]), .Q(s_A_ADDER[1]) );
  DLH_X1 \s_A_ADDER_reg[0]  ( .G(n325), .D(A[0]), .Q(s_A_ADDER[0]) );
  DLH_X1 \S_B_ADDER_reg[31]  ( .G(n326), .D(B[31]), .Q(S_B_ADDER[31]) );
  DLH_X1 \S_B_ADDER_reg[30]  ( .G(n328), .D(B[30]), .Q(S_B_ADDER[30]) );
  DLH_X1 \S_B_ADDER_reg[29]  ( .G(n328), .D(B[29]), .Q(S_B_ADDER[29]) );
  DLH_X1 \S_B_ADDER_reg[28]  ( .G(n327), .D(B[28]), .Q(S_B_ADDER[28]) );
  DLH_X1 \S_B_ADDER_reg[27]  ( .G(n329), .D(B[27]), .Q(S_B_ADDER[27]) );
  DLH_X1 \S_B_ADDER_reg[26]  ( .G(n329), .D(B[26]), .Q(S_B_ADDER[26]) );
  DLH_X1 \S_B_ADDER_reg[25]  ( .G(n329), .D(B[25]), .Q(S_B_ADDER[25]) );
  DLH_X1 \S_B_ADDER_reg[24]  ( .G(n329), .D(B[24]), .Q(S_B_ADDER[24]) );
  DLH_X1 \S_B_ADDER_reg[23]  ( .G(n329), .D(B[23]), .Q(S_B_ADDER[23]) );
  DLH_X1 \S_B_ADDER_reg[22]  ( .G(n330), .D(B[22]), .Q(S_B_ADDER[22]) );
  DLH_X1 \S_B_ADDER_reg[21]  ( .G(n330), .D(B[21]), .Q(S_B_ADDER[21]) );
  DLH_X1 \S_B_ADDER_reg[20]  ( .G(n329), .D(B[20]), .Q(S_B_ADDER[20]) );
  DLH_X1 \S_B_ADDER_reg[19]  ( .G(n330), .D(B[19]), .Q(S_B_ADDER[19]) );
  DLH_X1 \S_B_ADDER_reg[18]  ( .G(n330), .D(B[18]), .Q(S_B_ADDER[18]) );
  DLH_X1 \S_B_ADDER_reg[17]  ( .G(n330), .D(B[17]), .Q(S_B_ADDER[17]) );
  DLH_X1 \S_B_ADDER_reg[16]  ( .G(n329), .D(B[16]), .Q(S_B_ADDER[16]) );
  DLH_X1 \S_B_ADDER_reg[15]  ( .G(n331), .D(B[15]), .Q(S_B_ADDER[15]) );
  DLH_X1 \S_B_ADDER_reg[14]  ( .G(n330), .D(B[14]), .Q(S_B_ADDER[14]) );
  DLH_X1 \S_B_ADDER_reg[13]  ( .G(n330), .D(B[13]), .Q(S_B_ADDER[13]) );
  DLH_X1 \S_B_ADDER_reg[12]  ( .G(n329), .D(B[12]), .Q(S_B_ADDER[12]) );
  DLH_X1 \S_B_ADDER_reg[11]  ( .G(n329), .D(B[11]), .Q(S_B_ADDER[11]) );
  DLH_X1 \S_B_ADDER_reg[10]  ( .G(n329), .D(B[10]), .Q(S_B_ADDER[10]) );
  DLH_X1 \S_B_ADDER_reg[9]  ( .G(n326), .D(B[9]), .Q(S_B_ADDER[9]) );
  DLH_X1 \S_B_ADDER_reg[8]  ( .G(n326), .D(B[8]), .Q(S_B_ADDER[8]) );
  DLH_X1 \S_B_ADDER_reg[7]  ( .G(n327), .D(B[7]), .Q(S_B_ADDER[7]) );
  DLH_X1 \S_B_ADDER_reg[6]  ( .G(n327), .D(B[6]), .Q(S_B_ADDER[6]) );
  DLH_X1 \S_B_ADDER_reg[5]  ( .G(n327), .D(B[5]), .Q(S_B_ADDER[5]) );
  DLH_X1 \S_B_ADDER_reg[4]  ( .G(n328), .D(B[4]), .Q(S_B_ADDER[4]) );
  DLH_X1 \S_B_ADDER_reg[3]  ( .G(n328), .D(B[3]), .Q(S_B_ADDER[3]) );
  DLH_X1 \S_B_ADDER_reg[2]  ( .G(n328), .D(B[2]), .Q(S_B_ADDER[2]) );
  DLH_X1 \S_B_ADDER_reg[1]  ( .G(n328), .D(B[1]), .Q(S_B_ADDER[1]) );
  DLH_X1 \S_B_ADDER_reg[0]  ( .G(n330), .D(B[0]), .Q(S_B_ADDER[0]) );
  DLH_X1 \s_A_LOGIC_reg[31]  ( .G(n320), .D(A[31]), .Q(s_A_LOGIC[31]) );
  DLH_X1 \s_A_LOGIC_reg[30]  ( .G(n320), .D(A[30]), .Q(s_A_LOGIC[30]) );
  DLH_X1 \s_A_LOGIC_reg[29]  ( .G(n319), .D(A[29]), .Q(s_A_LOGIC[29]) );
  DLH_X1 \s_A_LOGIC_reg[28]  ( .G(n319), .D(A[28]), .Q(s_A_LOGIC[28]) );
  DLH_X1 \s_A_LOGIC_reg[27]  ( .G(n320), .D(A[27]), .Q(s_A_LOGIC[27]) );
  DLH_X1 \s_A_LOGIC_reg[26]  ( .G(n320), .D(A[26]), .Q(s_A_LOGIC[26]) );
  DLH_X1 \s_A_LOGIC_reg[25]  ( .G(n321), .D(A[25]), .Q(s_A_LOGIC[25]) );
  DLH_X1 \s_A_LOGIC_reg[24]  ( .G(n320), .D(A[24]), .Q(s_A_LOGIC[24]) );
  DLH_X1 \s_A_LOGIC_reg[23]  ( .G(n322), .D(A[23]), .Q(s_A_LOGIC[23]) );
  DLH_X1 \s_A_LOGIC_reg[22]  ( .G(n320), .D(A[22]), .Q(s_A_LOGIC[22]) );
  DLH_X1 \s_A_LOGIC_reg[21]  ( .G(n321), .D(A[21]), .Q(s_A_LOGIC[21]) );
  DLH_X1 \s_A_LOGIC_reg[20]  ( .G(n319), .D(A[20]), .Q(s_A_LOGIC[20]) );
  DLH_X1 \s_A_LOGIC_reg[19]  ( .G(n321), .D(A[19]), .Q(s_A_LOGIC[19]) );
  DLH_X1 \s_A_LOGIC_reg[18]  ( .G(n319), .D(A[18]), .Q(s_A_LOGIC[18]) );
  DLH_X1 \s_A_LOGIC_reg[17]  ( .G(n319), .D(A[17]), .Q(s_A_LOGIC[17]) );
  DLH_X1 \s_A_LOGIC_reg[16]  ( .G(n320), .D(A[16]), .Q(s_A_LOGIC[16]) );
  DLH_X1 \s_A_LOGIC_reg[15]  ( .G(n320), .D(A[15]), .Q(s_A_LOGIC[15]) );
  DLH_X1 \s_A_LOGIC_reg[14]  ( .G(n320), .D(A[14]), .Q(s_A_LOGIC[14]) );
  DLH_X1 \s_A_LOGIC_reg[13]  ( .G(n319), .D(A[13]), .Q(s_A_LOGIC[13]) );
  DLH_X1 \s_A_LOGIC_reg[12]  ( .G(n319), .D(A[12]), .Q(s_A_LOGIC[12]) );
  DLH_X1 \s_A_LOGIC_reg[11]  ( .G(n320), .D(A[11]), .Q(s_A_LOGIC[11]) );
  DLH_X1 \s_A_LOGIC_reg[10]  ( .G(n321), .D(A[10]), .Q(s_A_LOGIC[10]) );
  DLH_X1 \s_A_LOGIC_reg[9]  ( .G(n320), .D(A[9]), .Q(s_A_LOGIC[9]) );
  DLH_X1 \s_A_LOGIC_reg[8]  ( .G(n321), .D(A[8]), .Q(s_A_LOGIC[8]) );
  DLH_X1 \s_A_LOGIC_reg[7]  ( .G(n321), .D(A[7]), .Q(s_A_LOGIC[7]) );
  DLH_X1 \s_A_LOGIC_reg[6]  ( .G(n321), .D(A[6]), .Q(s_A_LOGIC[6]) );
  DLH_X1 \s_A_LOGIC_reg[5]  ( .G(n320), .D(A[5]), .Q(s_A_LOGIC[5]) );
  DLH_X1 \s_A_LOGIC_reg[4]  ( .G(n320), .D(A[4]), .Q(s_A_LOGIC[4]) );
  DLH_X1 \s_A_LOGIC_reg[3]  ( .G(n320), .D(A[3]), .Q(s_A_LOGIC[3]) );
  DLH_X1 \s_A_LOGIC_reg[2]  ( .G(n320), .D(A[2]), .Q(s_A_LOGIC[2]) );
  DLH_X1 \s_A_LOGIC_reg[1]  ( .G(n321), .D(A[1]), .Q(s_A_LOGIC[1]) );
  DLH_X1 \s_A_LOGIC_reg[0]  ( .G(n321), .D(A[0]), .Q(s_A_LOGIC[0]) );
  DLH_X1 \S_B_LOGIC_reg[31]  ( .G(n320), .D(B[31]), .Q(S_B_LOGIC[31]) );
  DLH_X1 \S_B_LOGIC_reg[30]  ( .G(n321), .D(B[30]), .Q(S_B_LOGIC[30]) );
  DLH_X1 \S_B_LOGIC_reg[29]  ( .G(n322), .D(B[29]), .Q(S_B_LOGIC[29]) );
  DLH_X1 \S_B_LOGIC_reg[28]  ( .G(n321), .D(B[28]), .Q(S_B_LOGIC[28]) );
  DLH_X1 \S_B_LOGIC_reg[27]  ( .G(n321), .D(B[27]), .Q(S_B_LOGIC[27]) );
  DLH_X1 \S_B_LOGIC_reg[26]  ( .G(n321), .D(B[26]), .Q(S_B_LOGIC[26]) );
  DLH_X1 \S_B_LOGIC_reg[25]  ( .G(n321), .D(B[25]), .Q(S_B_LOGIC[25]) );
  DLH_X1 \S_B_LOGIC_reg[24]  ( .G(n321), .D(B[24]), .Q(S_B_LOGIC[24]) );
  DLH_X1 \S_B_LOGIC_reg[23]  ( .G(n321), .D(B[23]), .Q(S_B_LOGIC[23]) );
  DLH_X1 \S_B_LOGIC_reg[22]  ( .G(n322), .D(B[22]), .Q(S_B_LOGIC[22]) );
  DLH_X1 \S_B_LOGIC_reg[21]  ( .G(n321), .D(B[21]), .Q(S_B_LOGIC[21]) );
  DLH_X1 \S_B_LOGIC_reg[20]  ( .G(n322), .D(B[20]), .Q(S_B_LOGIC[20]) );
  DLH_X1 \S_B_LOGIC_reg[19]  ( .G(n321), .D(B[19]), .Q(S_B_LOGIC[19]) );
  DLH_X1 \S_B_LOGIC_reg[18]  ( .G(n321), .D(B[18]), .Q(S_B_LOGIC[18]) );
  DLH_X1 \S_B_LOGIC_reg[17]  ( .G(n321), .D(B[17]), .Q(S_B_LOGIC[17]) );
  DLH_X1 \S_B_LOGIC_reg[16]  ( .G(n321), .D(B[16]), .Q(S_B_LOGIC[16]) );
  DLH_X1 \S_B_LOGIC_reg[15]  ( .G(n320), .D(B[15]), .Q(S_B_LOGIC[15]) );
  DLH_X1 \S_B_LOGIC_reg[14]  ( .G(n320), .D(B[14]), .Q(S_B_LOGIC[14]) );
  DLH_X1 \S_B_LOGIC_reg[13]  ( .G(n320), .D(B[13]), .Q(S_B_LOGIC[13]) );
  DLH_X1 \S_B_LOGIC_reg[12]  ( .G(n320), .D(B[12]), .Q(S_B_LOGIC[12]) );
  DLH_X1 \S_B_LOGIC_reg[11]  ( .G(n322), .D(B[11]), .Q(S_B_LOGIC[11]) );
  DLH_X1 \S_B_LOGIC_reg[10]  ( .G(n322), .D(B[10]), .Q(S_B_LOGIC[10]) );
  DLH_X1 \S_B_LOGIC_reg[9]  ( .G(n322), .D(B[9]), .Q(S_B_LOGIC[9]) );
  DLH_X1 \S_B_LOGIC_reg[8]  ( .G(n320), .D(B[8]), .Q(S_B_LOGIC[8]) );
  DLH_X1 \S_B_LOGIC_reg[7]  ( .G(n319), .D(B[7]), .Q(S_B_LOGIC[7]) );
  DLH_X1 \S_B_LOGIC_reg[6]  ( .G(n320), .D(B[6]), .Q(S_B_LOGIC[6]) );
  DLH_X1 \S_B_LOGIC_reg[5]  ( .G(n320), .D(B[5]), .Q(S_B_LOGIC[5]) );
  DLH_X1 \S_B_LOGIC_reg[4]  ( .G(n320), .D(B[4]), .Q(S_B_LOGIC[4]) );
  DLH_X1 \S_B_LOGIC_reg[3]  ( .G(n320), .D(B[3]), .Q(S_B_LOGIC[3]) );
  DLH_X1 \S_B_LOGIC_reg[2]  ( .G(n321), .D(B[2]), .Q(S_B_LOGIC[2]) );
  DLH_X1 \S_B_LOGIC_reg[1]  ( .G(n321), .D(B[1]), .Q(S_B_LOGIC[1]) );
  DLH_X1 \S_B_LOGIC_reg[0]  ( .G(n320), .D(B[0]), .Q(S_B_LOGIC[0]) );
  DLH_X1 \s_A_SHIFT_reg[31]  ( .G(n315), .D(A[31]), .Q(s_A_SHIFT[31]) );
  DLH_X1 \s_A_SHIFT_reg[30]  ( .G(n315), .D(A[30]), .Q(s_A_SHIFT[30]) );
  DLH_X1 \s_A_SHIFT_reg[29]  ( .G(n315), .D(A[29]), .Q(s_A_SHIFT[29]) );
  DLH_X1 \s_A_SHIFT_reg[28]  ( .G(n315), .D(A[28]), .Q(s_A_SHIFT[28]) );
  DLH_X1 \s_A_SHIFT_reg[27]  ( .G(n315), .D(A[27]), .Q(s_A_SHIFT[27]) );
  DLH_X1 \s_A_SHIFT_reg[26]  ( .G(n315), .D(A[26]), .Q(s_A_SHIFT[26]) );
  DLH_X1 \s_A_SHIFT_reg[25]  ( .G(n315), .D(A[25]), .Q(s_A_SHIFT[25]) );
  DLH_X1 \s_A_SHIFT_reg[24]  ( .G(n315), .D(A[24]), .Q(s_A_SHIFT[24]) );
  DLH_X1 \s_A_SHIFT_reg[23]  ( .G(n314), .D(A[23]), .Q(s_A_SHIFT[23]) );
  DLH_X1 \s_A_SHIFT_reg[22]  ( .G(n314), .D(A[22]), .Q(s_A_SHIFT[22]) );
  DLH_X1 \s_A_SHIFT_reg[21]  ( .G(n315), .D(A[21]), .Q(s_A_SHIFT[21]) );
  DLH_X1 \s_A_SHIFT_reg[20]  ( .G(n315), .D(A[20]), .Q(s_A_SHIFT[20]) );
  DLH_X1 \s_A_SHIFT_reg[19]  ( .G(n315), .D(A[19]), .Q(s_A_SHIFT[19]) );
  DLH_X1 \s_A_SHIFT_reg[18]  ( .G(n315), .D(A[18]), .Q(s_A_SHIFT[18]) );
  DLH_X1 \s_A_SHIFT_reg[17]  ( .G(n315), .D(A[17]), .Q(s_A_SHIFT[17]) );
  DLH_X1 \s_A_SHIFT_reg[16]  ( .G(n314), .D(A[16]), .Q(s_A_SHIFT[16]) );
  DLH_X1 \s_A_SHIFT_reg[15]  ( .G(n314), .D(A[15]), .Q(s_A_SHIFT[15]) );
  DLH_X1 \s_A_SHIFT_reg[14]  ( .G(n314), .D(A[14]), .Q(s_A_SHIFT[14]) );
  DLH_X1 \s_A_SHIFT_reg[13]  ( .G(n314), .D(A[13]), .Q(s_A_SHIFT[13]) );
  DLH_X1 \s_A_SHIFT_reg[12]  ( .G(n314), .D(A[12]), .Q(s_A_SHIFT[12]) );
  DLH_X1 \s_A_SHIFT_reg[11]  ( .G(n315), .D(A[11]), .Q(s_A_SHIFT[11]) );
  DLH_X1 \s_A_SHIFT_reg[10]  ( .G(n314), .D(A[10]), .Q(s_A_SHIFT[10]) );
  DLH_X1 \s_A_SHIFT_reg[9]  ( .G(n314), .D(A[9]), .Q(s_A_SHIFT[9]) );
  DLH_X1 \s_A_SHIFT_reg[8]  ( .G(n314), .D(A[8]), .Q(s_A_SHIFT[8]) );
  DLH_X1 \s_A_SHIFT_reg[7]  ( .G(n314), .D(A[7]), .Q(s_A_SHIFT[7]) );
  DLH_X1 \s_A_SHIFT_reg[6]  ( .G(n314), .D(A[6]), .Q(s_A_SHIFT[6]) );
  DLH_X1 \s_A_SHIFT_reg[5]  ( .G(n314), .D(A[5]), .Q(s_A_SHIFT[5]) );
  DLH_X1 \s_A_SHIFT_reg[4]  ( .G(n314), .D(A[4]), .Q(s_A_SHIFT[4]) );
  DLH_X1 \s_A_SHIFT_reg[3]  ( .G(n314), .D(A[3]), .Q(s_A_SHIFT[3]) );
  DLH_X1 \s_A_SHIFT_reg[2]  ( .G(n314), .D(A[2]), .Q(s_A_SHIFT[2]) );
  DLH_X1 \s_A_SHIFT_reg[1]  ( .G(n314), .D(A[1]), .Q(s_A_SHIFT[1]) );
  DLH_X1 \s_A_SHIFT_reg[0]  ( .G(n315), .D(A[0]), .Q(s_A_SHIFT[0]) );
  DLH_X1 \S_B_SHIFT_reg[31]  ( .G(n313), .D(B[31]), .Q(S_B_SHIFT[31]) );
  DLH_X1 \S_B_SHIFT_reg[30]  ( .G(n315), .D(B[30]), .Q(S_B_SHIFT[30]) );
  DLH_X1 \S_B_SHIFT_reg[29]  ( .G(n314), .D(B[29]), .Q(S_B_SHIFT[29]) );
  DLH_X1 \S_B_SHIFT_reg[28]  ( .G(n313), .D(B[28]), .Q(S_B_SHIFT[28]) );
  DLH_X1 \S_B_SHIFT_reg[27]  ( .G(n314), .D(B[27]), .Q(S_B_SHIFT[27]) );
  DLH_X1 \S_B_SHIFT_reg[26]  ( .G(n314), .D(B[26]), .Q(S_B_SHIFT[26]) );
  DLH_X1 \S_B_SHIFT_reg[25]  ( .G(n313), .D(B[25]), .Q(S_B_SHIFT[25]) );
  DLH_X1 \S_B_SHIFT_reg[24]  ( .G(n314), .D(B[24]), .Q(S_B_SHIFT[24]) );
  DLH_X1 \S_B_SHIFT_reg[23]  ( .G(n314), .D(B[23]), .Q(S_B_SHIFT[23]) );
  DLH_X1 \S_B_SHIFT_reg[22]  ( .G(n314), .D(B[22]), .Q(S_B_SHIFT[22]) );
  DLH_X1 \S_B_SHIFT_reg[21]  ( .G(n314), .D(B[21]), .Q(S_B_SHIFT[21]) );
  DLH_X1 \S_B_SHIFT_reg[20]  ( .G(n315), .D(B[20]), .Q(S_B_SHIFT[20]) );
  DLH_X1 \S_B_SHIFT_reg[19]  ( .G(n315), .D(B[19]), .Q(S_B_SHIFT[19]) );
  DLH_X1 \S_B_SHIFT_reg[18]  ( .G(n315), .D(B[18]), .Q(S_B_SHIFT[18]) );
  DLH_X1 \S_B_SHIFT_reg[17]  ( .G(n315), .D(B[17]), .Q(S_B_SHIFT[17]) );
  DLH_X1 \S_B_SHIFT_reg[16]  ( .G(n315), .D(B[16]), .Q(S_B_SHIFT[16]) );
  DLH_X1 \S_B_SHIFT_reg[15]  ( .G(n315), .D(B[15]), .Q(S_B_SHIFT[15]) );
  DLH_X1 \S_B_SHIFT_reg[14]  ( .G(n316), .D(B[14]), .Q(S_B_SHIFT[14]) );
  DLH_X1 \S_B_SHIFT_reg[13]  ( .G(n316), .D(B[13]), .Q(S_B_SHIFT[13]) );
  DLH_X1 \S_B_SHIFT_reg[12]  ( .G(n313), .D(B[12]), .Q(S_B_SHIFT[12]) );
  DLH_X1 \S_B_SHIFT_reg[11]  ( .G(n313), .D(B[11]), .Q(S_B_SHIFT[11]) );
  DLH_X1 \S_B_SHIFT_reg[10]  ( .G(n313), .D(B[10]), .Q(S_B_SHIFT[10]) );
  DLH_X1 \S_B_SHIFT_reg[9]  ( .G(n315), .D(B[9]), .Q(S_B_SHIFT[9]) );
  DLH_X1 \S_B_SHIFT_reg[8]  ( .G(n315), .D(B[8]), .Q(S_B_SHIFT[8]) );
  DLH_X1 \S_B_SHIFT_reg[7]  ( .G(n316), .D(B[7]), .Q(S_B_SHIFT[7]) );
  DLH_X1 \S_B_SHIFT_reg[6]  ( .G(n316), .D(B[6]), .Q(S_B_SHIFT[6]) );
  DLH_X1 \S_B_SHIFT_reg[5]  ( .G(n316), .D(B[5]), .Q(S_B_SHIFT[5]) );
  DLH_X1 \S_B_SHIFT_reg[4]  ( .G(n313), .D(B[4]), .Q(S_B_SHIFT[4]) );
  DLH_X1 \S_B_SHIFT_reg[3]  ( .G(n313), .D(B[3]), .Q(S_B_SHIFT[3]) );
  DLH_X1 \S_B_SHIFT_reg[2]  ( .G(n314), .D(B[2]), .Q(S_B_SHIFT[2]) );
  DLH_X1 \S_B_SHIFT_reg[1]  ( .G(n314), .D(B[1]), .Q(S_B_SHIFT[1]) );
  DLH_X1 \S_B_SHIFT_reg[0]  ( .G(n313), .D(B[0]), .Q(S_B_SHIFT[0]) );
  DLH_X1 \s_SHIFT_reg[1]  ( .G(n315), .D(n103), .Q(s_SHIFT[1]) );
  DLH_X1 \s_SHIFT_reg[0]  ( .G(n315), .D(n114), .Q(s_SHIFT[0]) );
  DLH_X1 \s_A_MULT_reg[15]  ( .G(n307), .D(A[15]), .Q(s_A_MULT[15]) );
  DLH_X1 \s_A_MULT_reg[14]  ( .G(n308), .D(A[14]), .Q(s_A_MULT[14]) );
  DLH_X1 \s_A_MULT_reg[13]  ( .G(n308), .D(A[13]), .Q(s_A_MULT[13]) );
  DLH_X1 \s_A_MULT_reg[12]  ( .G(n308), .D(A[12]), .Q(s_A_MULT[12]) );
  DLH_X1 \s_A_MULT_reg[11]  ( .G(n308), .D(A[11]), .Q(s_A_MULT[11]) );
  DLH_X1 \s_A_MULT_reg[10]  ( .G(n308), .D(A[10]), .Q(s_A_MULT[10]) );
  DLH_X1 \s_A_MULT_reg[9]  ( .G(n308), .D(A[9]), .Q(s_A_MULT[9]) );
  DLH_X1 \s_A_MULT_reg[8]  ( .G(n308), .D(A[8]), .Q(s_A_MULT[8]) );
  DLH_X1 \s_A_MULT_reg[7]  ( .G(n308), .D(A[7]), .Q(s_A_MULT[7]) );
  DLH_X1 \s_A_MULT_reg[6]  ( .G(n307), .D(A[6]), .Q(s_A_MULT[6]) );
  DLH_X1 \s_A_MULT_reg[5]  ( .G(n308), .D(A[5]), .Q(s_A_MULT[5]) );
  DLH_X1 \s_A_MULT_reg[4]  ( .G(n308), .D(A[4]), .Q(s_A_MULT[4]) );
  DLH_X1 \s_A_MULT_reg[3]  ( .G(n308), .D(A[3]), .Q(s_A_MULT[3]) );
  DLH_X1 \s_A_MULT_reg[2]  ( .G(n307), .D(A[2]), .Q(s_A_MULT[2]) );
  DLH_X1 \s_A_MULT_reg[1]  ( .G(n308), .D(A[1]), .Q(s_A_MULT[1]) );
  DLH_X1 \s_A_MULT_reg[0]  ( .G(n307), .D(A[0]), .Q(s_A_MULT[0]) );
  DLH_X1 \S_B_MULT_reg[15]  ( .G(n308), .D(B[15]), .Q(S_B_MULT[15]) );
  DLH_X1 \S_B_MULT_reg[14]  ( .G(n307), .D(B[14]), .Q(S_B_MULT[14]) );
  DLH_X1 \S_B_MULT_reg[13]  ( .G(n307), .D(B[13]), .Q(S_B_MULT[13]) );
  DLH_X1 \S_B_MULT_reg[12]  ( .G(n308), .D(B[12]), .Q(S_B_MULT[12]) );
  DLH_X1 \S_B_MULT_reg[11]  ( .G(n308), .D(B[11]), .Q(S_B_MULT[11]) );
  DLH_X1 \S_B_MULT_reg[10]  ( .G(n308), .D(B[10]), .Q(S_B_MULT[10]) );
  DLH_X1 \S_B_MULT_reg[9]  ( .G(n308), .D(B[9]), .Q(S_B_MULT[9]) );
  DLH_X1 \S_B_MULT_reg[8]  ( .G(n308), .D(B[8]), .Q(S_B_MULT[8]) );
  DLH_X1 \S_B_MULT_reg[7]  ( .G(n307), .D(B[7]), .Q(S_B_MULT[7]) );
  DLH_X1 \S_B_MULT_reg[6]  ( .G(n307), .D(B[6]), .Q(S_B_MULT[6]) );
  DLH_X1 \S_B_MULT_reg[5]  ( .G(n308), .D(B[5]), .Q(S_B_MULT[5]) );
  DLH_X1 \S_B_MULT_reg[4]  ( .G(n308), .D(B[4]), .Q(S_B_MULT[4]) );
  DLH_X1 \S_B_MULT_reg[3]  ( .G(n308), .D(B[3]), .Q(S_B_MULT[3]) );
  DLH_X1 \S_B_MULT_reg[2]  ( .G(n308), .D(B[2]), .Q(S_B_MULT[2]) );
  DLH_X1 \S_B_MULT_reg[1]  ( .G(n308), .D(B[1]), .Q(S_B_MULT[1]) );
  DLH_X1 \S_B_MULT_reg[0]  ( .G(n308), .D(B[0]), .Q(S_B_MULT[0]) );
  DLH_X1 \S_B_LHI_reg[15]  ( .G(n310), .D(B[15]), .Q(S_B_LHI[15]) );
  DLH_X1 \S_B_LHI_reg[14]  ( .G(n310), .D(B[14]), .Q(S_B_LHI[14]) );
  DLH_X1 \S_B_LHI_reg[13]  ( .G(n310), .D(B[13]), .Q(S_B_LHI[13]) );
  DLH_X1 \S_B_LHI_reg[12]  ( .G(n310), .D(B[12]), .Q(S_B_LHI[12]) );
  DLH_X1 \S_B_LHI_reg[11]  ( .G(n310), .D(B[11]), .Q(S_B_LHI[11]) );
  DLH_X1 \S_B_LHI_reg[10]  ( .G(n310), .D(B[10]), .Q(S_B_LHI[10]) );
  DLH_X1 \S_B_LHI_reg[9]  ( .G(n310), .D(B[9]), .Q(S_B_LHI[9]) );
  DLH_X1 \S_B_LHI_reg[8]  ( .G(n310), .D(B[8]), .Q(S_B_LHI[8]) );
  DLH_X1 \S_B_LHI_reg[7]  ( .G(n310), .D(B[7]), .Q(S_B_LHI[7]) );
  DLH_X1 \S_B_LHI_reg[6]  ( .G(n310), .D(B[6]), .Q(S_B_LHI[6]) );
  DLH_X1 \S_B_LHI_reg[5]  ( .G(n310), .D(B[5]), .Q(S_B_LHI[5]) );
  DLH_X1 \S_B_LHI_reg[4]  ( .G(n310), .D(B[4]), .Q(S_B_LHI[4]) );
  DLH_X1 \S_B_LHI_reg[3]  ( .G(n310), .D(B[3]), .Q(S_B_LHI[3]) );
  DLH_X1 \S_B_LHI_reg[2]  ( .G(n310), .D(B[2]), .Q(S_B_LHI[2]) );
  DLH_X1 \S_B_LHI_reg[1]  ( .G(n310), .D(B[1]), .Q(S_B_LHI[1]) );
  DLH_X1 \S_B_LHI_reg[0]  ( .G(n310), .D(B[0]), .Q(S_B_LHI[0]) );
  DLH_X1 s_ADD_SUB_reg ( .G(n325), .D(n110), .Q(s_ADD_SUB) );
  DLH_X1 \s_LOGIC_reg[3]  ( .G(n321), .D(N24), .Q(s_LOGIC[3]) );
  DLH_X1 \s_LOGIC_reg[2]  ( .G(n321), .D(n334), .Q(s_LOGIC[2]) );
  DLH_X1 \s_LOGIC_reg[1]  ( .G(n321), .D(n334), .Q(s_LOGIC[1]) );
  XOR2_X1 U142 ( .A(s_SIGN), .B(s_Co), .Z(s_C) );
  NAND3_X1 U143 ( .A1(n81), .A2(n82), .A3(n83), .ZN(Y[0]) );
  OAI33_X1 U144 ( .A1(n338), .A2(s_NE), .A3(n341), .B1(n344), .B2(s_LE), .B3(
        n86), .ZN(n85) );
  OAI33_X1 U145 ( .A1(n90), .A2(n3), .A3(OP[2]), .B1(n342), .B2(n207), .B3(n86), .ZN(n89) );
  NAND3_X1 U146 ( .A1(OP[2]), .A2(n345), .A3(n97), .ZN(n17) );
  NAND3_X1 U147 ( .A1(n345), .A2(n340), .A3(OP[4]), .ZN(n90) );
  ADDER_SUBTRACTOR_WIDTH32_RADIX4 ADD_SUB ( .A(s_A_ADDER), .B(S_B_ADDER), .Ci(
        s_ADD_SUB), .S(s_OUT), .Co(s_Co) );
  ZERO_DETECTOR_WIDTH32_1 BIG_XNOR ( .A(s_OUT), .Y(s_Z) );
  LOGIC_WIDTH32 LOGICALS ( .R1(s_A_LOGIC), .R2(S_B_LOGIC), .S0(1'b0), .S1(
        s_LOGIC[1]), .S2(s_LOGIC[2]), .S3(s_LOGIC[3]), .Y(s_LOG) );
  COMPARATOR COMP ( .Z(s_Z), .C(s_C), .LE(s_LE), .LT(n206), .GE(n115), .GT(
        n207), .EQ(n3), .NE(s_NE) );
  SHIFTER_WIDTH32 SHIFT ( .R1(s_A_SHIFT), .R2(S_B_SHIFT), .SEL(s_SHIFT), .Y(
        s_SHI) );
  MULTIPLIER_WIDTH16 MULT ( .A(s_A_MULT), .B(S_B_MULT), .P({s_MULT[31], 
        SYNOPSYS_UNCONNECTED__0, s_MULT[29:0]}) );
  BUF_X1 U3 ( .A(n303), .Z(n305) );
  BUF_X1 U4 ( .A(n303), .Z(n306) );
  BUF_X1 U5 ( .A(n304), .Z(n307) );
  BUF_X1 U6 ( .A(n304), .Z(n308) );
  BUF_X1 U7 ( .A(n112), .Z(n309) );
  BUF_X1 U8 ( .A(n112), .Z(n310) );
  BUF_X1 U9 ( .A(n109), .Z(n303) );
  BUF_X1 U10 ( .A(n109), .Z(n304) );
  BUF_X1 U11 ( .A(N25), .Z(n311) );
  BUF_X1 U12 ( .A(N22), .Z(n317) );
  BUF_X1 U13 ( .A(N22), .Z(n318) );
  BUF_X1 U14 ( .A(N25), .Z(n312) );
  BUF_X1 U15 ( .A(N25), .Z(n313) );
  BUF_X1 U16 ( .A(N22), .Z(n319) );
  BUF_X1 U17 ( .A(n333), .Z(n300) );
  BUF_X1 U18 ( .A(n333), .Z(n301) );
  BUF_X1 U19 ( .A(n333), .Z(n302) );
  NOR2_X1 U20 ( .A1(n343), .A2(n337), .ZN(n103) );
  NOR2_X1 U21 ( .A1(n343), .A2(n338), .ZN(n112) );
  NOR2_X1 U22 ( .A1(n344), .A2(n337), .ZN(n109) );
  INV_X1 U23 ( .A(n92), .ZN(n341) );
  INV_X1 U24 ( .A(n104), .ZN(n336) );
  BUF_X1 U25 ( .A(N20), .Z(n323) );
  BUF_X1 U26 ( .A(N20), .Z(n324) );
  AOI222_X1 U27 ( .A1(s_SHI[16]), .A2(n312), .B1(s_OUT[16]), .B2(n302), .C1(
        s_LOG[16]), .C2(n318), .ZN(n68) );
  AOI222_X1 U28 ( .A1(s_SHI[17]), .A2(n312), .B1(s_OUT[17]), .B2(n302), .C1(
        s_LOG[17]), .C2(n318), .ZN(n66) );
  AOI222_X1 U29 ( .A1(s_SHI[18]), .A2(n313), .B1(s_OUT[18]), .B2(n302), .C1(
        s_LOG[18]), .C2(n319), .ZN(n64) );
  AOI222_X1 U30 ( .A1(s_SHI[27]), .A2(n313), .B1(s_OUT[27]), .B2(n302), .C1(
        s_LOG[27]), .C2(n319), .ZN(n44) );
  AOI222_X1 U31 ( .A1(s_SHI[28]), .A2(n313), .B1(s_OUT[28]), .B2(n302), .C1(
        s_LOG[28]), .C2(n319), .ZN(n42) );
  AOI222_X1 U32 ( .A1(s_SHI[29]), .A2(n312), .B1(s_OUT[29]), .B2(n302), .C1(
        s_LOG[29]), .C2(n318), .ZN(n40) );
  AOI222_X1 U33 ( .A1(s_SHI[30]), .A2(n313), .B1(s_OUT[30]), .B2(n302), .C1(
        s_LOG[30]), .C2(n319), .ZN(n36) );
  AOI222_X1 U34 ( .A1(s_SHI[31]), .A2(n313), .B1(s_OUT[31]), .B2(n302), .C1(
        s_LOG[31]), .C2(n319), .ZN(n34) );
  AOI222_X1 U35 ( .A1(s_SHI[19]), .A2(n312), .B1(s_OUT[19]), .B2(n301), .C1(
        s_LOG[19]), .C2(n318), .ZN(n62) );
  AOI222_X1 U36 ( .A1(s_SHI[20]), .A2(n313), .B1(s_OUT[20]), .B2(n301), .C1(
        s_LOG[20]), .C2(n319), .ZN(n58) );
  AOI222_X1 U37 ( .A1(s_SHI[21]), .A2(n312), .B1(s_OUT[21]), .B2(n301), .C1(
        s_LOG[21]), .C2(n318), .ZN(n56) );
  AOI222_X1 U38 ( .A1(s_SHI[22]), .A2(n312), .B1(s_OUT[22]), .B2(n301), .C1(
        s_LOG[22]), .C2(n318), .ZN(n54) );
  AOI222_X1 U39 ( .A1(s_SHI[23]), .A2(n312), .B1(s_OUT[23]), .B2(n301), .C1(
        s_LOG[23]), .C2(n318), .ZN(n52) );
  AOI222_X1 U40 ( .A1(s_SHI[24]), .A2(n313), .B1(s_OUT[24]), .B2(n301), .C1(
        s_LOG[24]), .C2(n319), .ZN(n50) );
  AOI222_X1 U41 ( .A1(s_SHI[25]), .A2(n312), .B1(s_OUT[25]), .B2(n301), .C1(
        s_LOG[25]), .C2(n318), .ZN(n48) );
  AOI222_X1 U42 ( .A1(s_SHI[26]), .A2(n313), .B1(s_OUT[26]), .B2(n301), .C1(
        s_LOG[26]), .C2(n319), .ZN(n46) );
  NOR2_X1 U43 ( .A1(n346), .A2(n342), .ZN(n92) );
  AOI221_X1 U44 ( .B1(n206), .B2(n84), .C1(n332), .C2(n346), .A(n85), .ZN(n83)
         );
  OAI22_X1 U45 ( .A1(n337), .A2(n341), .B1(n346), .B2(n91), .ZN(n84) );
  OAI21_X1 U46 ( .B1(n344), .B2(n18), .A(n17), .ZN(N22) );
  AOI22_X1 U47 ( .A1(s_SHI[1]), .A2(n311), .B1(s_MULT[1]), .B2(n307), .ZN(n59)
         );
  AOI22_X1 U48 ( .A1(s_SHI[3]), .A2(n311), .B1(s_MULT[3]), .B2(n306), .ZN(n31)
         );
  AOI22_X1 U49 ( .A1(s_SHI[7]), .A2(n311), .B1(s_MULT[7]), .B2(n306), .ZN(n23)
         );
  AOI22_X1 U50 ( .A1(s_SHI[11]), .A2(n311), .B1(s_MULT[11]), .B2(n307), .ZN(
        n77) );
  AOI22_X1 U51 ( .A1(s_SHI[13]), .A2(n311), .B1(s_MULT[13]), .B2(n307), .ZN(
        n73) );
  AOI22_X1 U52 ( .A1(s_SHI[15]), .A2(n311), .B1(s_MULT[15]), .B2(n307), .ZN(
        n69) );
  AOI22_X1 U53 ( .A1(s_SHI[5]), .A2(n312), .B1(s_MULT[5]), .B2(n306), .ZN(n27)
         );
  AOI22_X1 U54 ( .A1(s_SHI[9]), .A2(n312), .B1(s_MULT[9]), .B2(n306), .ZN(n19)
         );
  INV_X1 U55 ( .A(n101), .ZN(n337) );
  INV_X1 U56 ( .A(n100), .ZN(n338) );
  INV_X1 U57 ( .A(n98), .ZN(n344) );
  INV_X1 U58 ( .A(n96), .ZN(n343) );
  INV_X1 U59 ( .A(n93), .ZN(n333) );
  AND2_X1 U60 ( .A1(n90), .A2(n338), .ZN(n86) );
  OAI21_X1 U61 ( .B1(n342), .B2(n18), .A(n335), .ZN(N25) );
  INV_X1 U62 ( .A(n103), .ZN(n335) );
  OAI211_X1 U63 ( .C1(n92), .C2(n90), .A(n94), .B(n99), .ZN(n104) );
  AOI21_X1 U64 ( .B1(n100), .B2(n92), .A(n339), .ZN(n99) );
  INV_X1 U65 ( .A(n91), .ZN(n339) );
  OAI21_X1 U66 ( .B1(n18), .B2(n343), .A(n336), .ZN(n110) );
  NAND2_X1 U67 ( .A1(n93), .A2(n336), .ZN(N20) );
  NOR2_X1 U68 ( .A1(n94), .A2(n95), .ZN(N27) );
  XNOR2_X1 U69 ( .A(B[31]), .B(A[31]), .ZN(n95) );
  NOR2_X1 U70 ( .A1(n341), .A2(n18), .ZN(n114) );
  INV_X1 U71 ( .A(n17), .ZN(n334) );
  NOR3_X1 U72 ( .A1(n340), .A2(OP[4]), .A3(n345), .ZN(n100) );
  OAI221_X1 U73 ( .B1(n96), .B2(n345), .C1(OP[1]), .C2(n98), .A(n97), .ZN(n93)
         );
  NOR3_X1 U74 ( .A1(OP[1]), .A2(OP[4]), .A3(n340), .ZN(n101) );
  NOR2_X1 U75 ( .A1(n346), .A2(OP[2]), .ZN(n98) );
  NAND4_X1 U76 ( .A1(OP[4]), .A2(OP[1]), .A3(n342), .A4(n340), .ZN(n91) );
  NOR2_X1 U77 ( .A1(OP[4]), .A2(OP[3]), .ZN(n97) );
  NAND2_X1 U78 ( .A1(n97), .A2(OP[1]), .ZN(n18) );
  INV_X1 U79 ( .A(OP[2]), .ZN(n342) );
  AOI22_X1 U80 ( .A1(s_OUT[0]), .A2(n300), .B1(s_LOG[0]), .B2(n317), .ZN(n82)
         );
  NAND2_X1 U81 ( .A1(n59), .A2(n60), .ZN(Y[1]) );
  AOI22_X1 U82 ( .A1(s_OUT[1]), .A2(n300), .B1(s_LOG[1]), .B2(n317), .ZN(n60)
         );
  NAND2_X1 U83 ( .A1(n37), .A2(n38), .ZN(Y[2]) );
  AOI22_X1 U84 ( .A1(s_OUT[2]), .A2(n300), .B1(s_LOG[2]), .B2(n317), .ZN(n38)
         );
  NAND2_X1 U85 ( .A1(n31), .A2(n32), .ZN(Y[3]) );
  AOI22_X1 U86 ( .A1(s_OUT[3]), .A2(n300), .B1(s_LOG[3]), .B2(n317), .ZN(n32)
         );
  NAND2_X1 U87 ( .A1(n29), .A2(n30), .ZN(Y[4]) );
  AOI22_X1 U88 ( .A1(s_OUT[4]), .A2(n300), .B1(s_LOG[4]), .B2(n317), .ZN(n30)
         );
  NAND2_X1 U89 ( .A1(n23), .A2(n24), .ZN(Y[7]) );
  AOI22_X1 U90 ( .A1(s_OUT[7]), .A2(n300), .B1(s_LOG[7]), .B2(n317), .ZN(n24)
         );
  AOI22_X1 U91 ( .A1(s_SHI[2]), .A2(n311), .B1(s_MULT[2]), .B2(n307), .ZN(n37)
         );
  AOI22_X1 U92 ( .A1(s_SHI[4]), .A2(n311), .B1(s_MULT[4]), .B2(n306), .ZN(n29)
         );
  AOI22_X1 U93 ( .A1(s_SHI[10]), .A2(n311), .B1(s_MULT[10]), .B2(n307), .ZN(
        n79) );
  AOI22_X1 U94 ( .A1(s_SHI[12]), .A2(n311), .B1(s_MULT[12]), .B2(n307), .ZN(
        n75) );
  AOI22_X1 U95 ( .A1(s_SHI[14]), .A2(n311), .B1(s_MULT[14]), .B2(n307), .ZN(
        n71) );
  AOI22_X1 U96 ( .A1(s_SHI[6]), .A2(n312), .B1(s_MULT[6]), .B2(n306), .ZN(n25)
         );
  AOI22_X1 U97 ( .A1(s_SHI[8]), .A2(n312), .B1(s_MULT[8]), .B2(n306), .ZN(n21)
         );
  NOR2_X1 U98 ( .A1(OP[0]), .A2(OP[2]), .ZN(n96) );
  NAND2_X1 U99 ( .A1(n79), .A2(n80), .ZN(Y[10]) );
  AOI22_X1 U100 ( .A1(s_OUT[10]), .A2(n300), .B1(s_LOG[10]), .B2(n317), .ZN(
        n80) );
  NAND2_X1 U101 ( .A1(n77), .A2(n78), .ZN(Y[11]) );
  AOI22_X1 U102 ( .A1(s_OUT[11]), .A2(n301), .B1(s_LOG[11]), .B2(n317), .ZN(
        n78) );
  NAND2_X1 U103 ( .A1(n75), .A2(n76), .ZN(Y[12]) );
  AOI22_X1 U104 ( .A1(s_OUT[12]), .A2(n301), .B1(s_LOG[12]), .B2(n317), .ZN(
        n76) );
  NAND2_X1 U105 ( .A1(n73), .A2(n74), .ZN(Y[13]) );
  AOI22_X1 U106 ( .A1(s_OUT[13]), .A2(n301), .B1(s_LOG[13]), .B2(n317), .ZN(
        n74) );
  NAND2_X1 U107 ( .A1(n71), .A2(n72), .ZN(Y[14]) );
  AOI22_X1 U108 ( .A1(s_OUT[14]), .A2(n300), .B1(s_LOG[14]), .B2(n317), .ZN(
        n72) );
  NAND2_X1 U109 ( .A1(n69), .A2(n70), .ZN(Y[15]) );
  AOI22_X1 U110 ( .A1(s_OUT[15]), .A2(n301), .B1(s_LOG[15]), .B2(n317), .ZN(
        n70) );
  NAND2_X1 U111 ( .A1(n67), .A2(n68), .ZN(Y[16]) );
  AOI22_X1 U112 ( .A1(s_MULT[16]), .A2(n305), .B1(S_B_LHI[0]), .B2(n309), .ZN(
        n67) );
  NAND2_X1 U113 ( .A1(n65), .A2(n66), .ZN(Y[17]) );
  AOI22_X1 U114 ( .A1(s_MULT[17]), .A2(n305), .B1(S_B_LHI[1]), .B2(n309), .ZN(
        n65) );
  NAND2_X1 U115 ( .A1(n61), .A2(n62), .ZN(Y[19]) );
  AOI22_X1 U116 ( .A1(s_MULT[19]), .A2(n305), .B1(S_B_LHI[3]), .B2(n309), .ZN(
        n61) );
  NAND2_X1 U117 ( .A1(n55), .A2(n56), .ZN(Y[21]) );
  AOI22_X1 U118 ( .A1(s_MULT[21]), .A2(n305), .B1(S_B_LHI[5]), .B2(n309), .ZN(
        n55) );
  NAND2_X1 U119 ( .A1(n53), .A2(n54), .ZN(Y[22]) );
  AOI22_X1 U120 ( .A1(s_MULT[22]), .A2(n305), .B1(S_B_LHI[6]), .B2(n309), .ZN(
        n53) );
  NAND2_X1 U121 ( .A1(n51), .A2(n52), .ZN(Y[23]) );
  AOI22_X1 U122 ( .A1(s_MULT[23]), .A2(n305), .B1(S_B_LHI[7]), .B2(n309), .ZN(
        n51) );
  NAND2_X1 U123 ( .A1(n47), .A2(n48), .ZN(Y[25]) );
  AOI22_X1 U124 ( .A1(s_MULT[25]), .A2(n306), .B1(S_B_LHI[9]), .B2(n309), .ZN(
        n47) );
  NAND2_X1 U125 ( .A1(n39), .A2(n40), .ZN(Y[29]) );
  AOI22_X1 U126 ( .A1(s_MULT[29]), .A2(n306), .B1(S_B_LHI[13]), .B2(n310), 
        .ZN(n39) );
  AOI22_X1 U127 ( .A1(s_SHI[0]), .A2(n311), .B1(s_MULT[0]), .B2(n306), .ZN(n81) );
  INV_X1 U128 ( .A(OP[0]), .ZN(n346) );
  INV_X1 U129 ( .A(OP[3]), .ZN(n340) );
  INV_X1 U130 ( .A(OP[1]), .ZN(n345) );
  INV_X1 U131 ( .A(n87), .ZN(n332) );
  AOI21_X1 U132 ( .B1(n115), .B2(n88), .A(n89), .ZN(n87) );
  OAI21_X1 U133 ( .B1(n342), .B2(n337), .A(n91), .ZN(n88) );
  NAND2_X1 U134 ( .A1(n63), .A2(n64), .ZN(Y[18]) );
  AOI22_X1 U135 ( .A1(s_MULT[18]), .A2(n305), .B1(S_B_LHI[2]), .B2(n309), .ZN(
        n63) );
  NAND2_X1 U136 ( .A1(n57), .A2(n58), .ZN(Y[20]) );
  AOI22_X1 U137 ( .A1(s_MULT[20]), .A2(n305), .B1(S_B_LHI[4]), .B2(n309), .ZN(
        n57) );
  NAND2_X1 U138 ( .A1(n49), .A2(n50), .ZN(Y[24]) );
  AOI22_X1 U139 ( .A1(s_MULT[24]), .A2(n305), .B1(S_B_LHI[8]), .B2(n309), .ZN(
        n49) );
  NAND2_X1 U140 ( .A1(n45), .A2(n46), .ZN(Y[26]) );
  AOI22_X1 U141 ( .A1(s_MULT[26]), .A2(n305), .B1(S_B_LHI[10]), .B2(n309), 
        .ZN(n45) );
  NAND2_X1 U148 ( .A1(n43), .A2(n44), .ZN(Y[27]) );
  AOI22_X1 U149 ( .A1(s_MULT[27]), .A2(n306), .B1(S_B_LHI[11]), .B2(n309), 
        .ZN(n43) );
  NAND2_X1 U150 ( .A1(n41), .A2(n42), .ZN(Y[28]) );
  AOI22_X1 U151 ( .A1(s_MULT[28]), .A2(n306), .B1(S_B_LHI[12]), .B2(n310), 
        .ZN(n41) );
  NAND2_X1 U152 ( .A1(n35), .A2(n36), .ZN(Y[30]) );
  AOI22_X1 U153 ( .A1(s_MULT[31]), .A2(n305), .B1(S_B_LHI[14]), .B2(n310), 
        .ZN(n35) );
  NAND2_X1 U154 ( .A1(n33), .A2(n34), .ZN(Y[31]) );
  AOI22_X1 U155 ( .A1(s_MULT[31]), .A2(n305), .B1(S_B_LHI[15]), .B2(n310), 
        .ZN(n33) );
  NAND2_X1 U156 ( .A1(n27), .A2(n28), .ZN(Y[5]) );
  AOI22_X1 U157 ( .A1(s_OUT[5]), .A2(n300), .B1(s_LOG[5]), .B2(n318), .ZN(n28)
         );
  NAND2_X1 U158 ( .A1(n25), .A2(n26), .ZN(Y[6]) );
  AOI22_X1 U159 ( .A1(s_OUT[6]), .A2(n300), .B1(s_LOG[6]), .B2(n318), .ZN(n26)
         );
  NAND2_X1 U160 ( .A1(n21), .A2(n22), .ZN(Y[8]) );
  AOI22_X1 U161 ( .A1(s_OUT[8]), .A2(n300), .B1(s_LOG[8]), .B2(n318), .ZN(n22)
         );
  NAND2_X1 U162 ( .A1(n19), .A2(n20), .ZN(Y[9]) );
  AOI22_X1 U163 ( .A1(s_OUT[9]), .A2(n300), .B1(s_LOG[9]), .B2(n318), .ZN(n20)
         );
  AOI221_X1 U164 ( .B1(n101), .B2(n92), .C1(n98), .C2(n100), .A(n102), .ZN(n94) );
  AOI211_X1 U165 ( .C1(n337), .C2(n338), .A(OP[0]), .B(n342), .ZN(n102) );
  OAI22_X1 U166 ( .A1(OP[0]), .A2(n17), .B1(n344), .B2(n18), .ZN(N24) );
  CLKBUF_X1 U167 ( .A(N25), .Z(n314) );
  CLKBUF_X1 U168 ( .A(N25), .Z(n315) );
  CLKBUF_X1 U169 ( .A(N25), .Z(n316) );
  CLKBUF_X1 U170 ( .A(N22), .Z(n320) );
  CLKBUF_X1 U171 ( .A(N22), .Z(n321) );
  CLKBUF_X1 U172 ( .A(N22), .Z(n322) );
  CLKBUF_X1 U173 ( .A(n323), .Z(n325) );
  CLKBUF_X1 U174 ( .A(n323), .Z(n326) );
  CLKBUF_X1 U175 ( .A(n323), .Z(n327) );
  CLKBUF_X1 U176 ( .A(n323), .Z(n328) );
  CLKBUF_X1 U177 ( .A(n324), .Z(n329) );
  CLKBUF_X1 U178 ( .A(n324), .Z(n330) );
  CLKBUF_X1 U179 ( .A(n324), .Z(n331) );
endmodule


module REGISTER_GENERIC_WIDTH32_6 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298;

  DFF_X1 \DOUT_reg[31]  ( .D(n68), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[30]  ( .D(n69), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[29]  ( .D(n70), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[28]  ( .D(n71), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[27]  ( .D(n72), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n73), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[25]  ( .D(n74), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[24]  ( .D(n75), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[22]  ( .D(n77), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[21]  ( .D(n78), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[20]  ( .D(n79), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n80), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n81), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n83), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n84), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n89), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n90), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n91), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n92), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n93), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n94), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n95), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n96), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n97), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n98), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n262) );
  BUF_X1 U4 ( .A(n35), .Z(n261) );
  BUF_X1 U5 ( .A(n35), .Z(n260) );
  BUF_X1 U6 ( .A(n34), .Z(n265) );
  NAND2_X1 U7 ( .A1(RST), .A2(n263), .ZN(n35) );
  BUF_X1 U8 ( .A(n34), .Z(n263) );
  BUF_X1 U9 ( .A(n34), .Z(n264) );
  OAI22_X1 U10 ( .A1(n36), .A2(n265), .B1(n262), .B2(n266), .ZN(n99) );
  INV_X1 U11 ( .A(DIN[0]), .ZN(n266) );
  OAI22_X1 U12 ( .A1(n37), .A2(n265), .B1(n262), .B2(n277), .ZN(n98) );
  INV_X1 U13 ( .A(DIN[1]), .ZN(n277) );
  OAI22_X1 U14 ( .A1(n38), .A2(n265), .B1(n262), .B2(n276), .ZN(n97) );
  INV_X1 U15 ( .A(DIN[2]), .ZN(n276) );
  OAI22_X1 U16 ( .A1(n39), .A2(n265), .B1(n262), .B2(n275), .ZN(n96) );
  INV_X1 U17 ( .A(DIN[3]), .ZN(n275) );
  OAI22_X1 U18 ( .A1(n40), .A2(n265), .B1(n262), .B2(n281), .ZN(n95) );
  INV_X1 U19 ( .A(DIN[4]), .ZN(n281) );
  OAI22_X1 U20 ( .A1(n43), .A2(n265), .B1(n262), .B2(n278), .ZN(n92) );
  INV_X1 U21 ( .A(DIN[7]), .ZN(n278) );
  OAI22_X1 U22 ( .A1(n46), .A2(n264), .B1(n261), .B2(n283), .ZN(n89) );
  INV_X1 U23 ( .A(DIN[10]), .ZN(n283) );
  OAI22_X1 U24 ( .A1(n47), .A2(n264), .B1(n261), .B2(n282), .ZN(n88) );
  INV_X1 U25 ( .A(DIN[11]), .ZN(n282) );
  OAI22_X1 U26 ( .A1(n48), .A2(n264), .B1(n261), .B2(n274), .ZN(n87) );
  INV_X1 U27 ( .A(DIN[12]), .ZN(n274) );
  OAI22_X1 U28 ( .A1(n49), .A2(n264), .B1(n261), .B2(n273), .ZN(n86) );
  INV_X1 U29 ( .A(DIN[13]), .ZN(n273) );
  OAI22_X1 U30 ( .A1(n50), .A2(n264), .B1(n261), .B2(n272), .ZN(n85) );
  INV_X1 U31 ( .A(DIN[14]), .ZN(n272) );
  OAI22_X1 U32 ( .A1(n51), .A2(n264), .B1(n261), .B2(n271), .ZN(n84) );
  INV_X1 U33 ( .A(DIN[15]), .ZN(n271) );
  OAI22_X1 U34 ( .A1(n52), .A2(n264), .B1(n261), .B2(n289), .ZN(n83) );
  INV_X1 U35 ( .A(DIN[16]), .ZN(n289) );
  OAI22_X1 U36 ( .A1(n53), .A2(n264), .B1(n261), .B2(n288), .ZN(n82) );
  INV_X1 U37 ( .A(DIN[17]), .ZN(n288) );
  OAI22_X1 U38 ( .A1(n55), .A2(n264), .B1(n261), .B2(n286), .ZN(n80) );
  INV_X1 U39 ( .A(DIN[19]), .ZN(n286) );
  OAI22_X1 U40 ( .A1(n57), .A2(n263), .B1(n260), .B2(n269), .ZN(n78) );
  INV_X1 U41 ( .A(DIN[21]), .ZN(n269) );
  OAI22_X1 U42 ( .A1(n58), .A2(n263), .B1(n260), .B2(n268), .ZN(n77) );
  INV_X1 U43 ( .A(DIN[22]), .ZN(n268) );
  OAI22_X1 U44 ( .A1(n59), .A2(n263), .B1(n260), .B2(n267), .ZN(n76) );
  INV_X1 U45 ( .A(DIN[23]), .ZN(n267) );
  OAI22_X1 U46 ( .A1(n61), .A2(n263), .B1(n260), .B2(n292), .ZN(n74) );
  INV_X1 U47 ( .A(DIN[25]), .ZN(n292) );
  OAI22_X1 U48 ( .A1(n65), .A2(n263), .B1(n260), .B2(n296), .ZN(n70) );
  INV_X1 U49 ( .A(DIN[29]), .ZN(n296) );
  NAND2_X1 U50 ( .A1(n298), .A2(RST), .ZN(n34) );
  INV_X1 U51 ( .A(EN), .ZN(n298) );
  OAI22_X1 U52 ( .A1(n54), .A2(n264), .B1(n261), .B2(n287), .ZN(n81) );
  INV_X1 U53 ( .A(DIN[18]), .ZN(n287) );
  OAI22_X1 U54 ( .A1(n56), .A2(n264), .B1(n261), .B2(n270), .ZN(n79) );
  INV_X1 U55 ( .A(DIN[20]), .ZN(n270) );
  OAI22_X1 U56 ( .A1(n60), .A2(n263), .B1(n260), .B2(n293), .ZN(n75) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n293) );
  OAI22_X1 U58 ( .A1(n62), .A2(n263), .B1(n260), .B2(n291), .ZN(n73) );
  INV_X1 U59 ( .A(DIN[26]), .ZN(n291) );
  OAI22_X1 U60 ( .A1(n63), .A2(n263), .B1(n260), .B2(n290), .ZN(n72) );
  INV_X1 U61 ( .A(DIN[27]), .ZN(n290) );
  OAI22_X1 U62 ( .A1(n64), .A2(n263), .B1(n260), .B2(n297), .ZN(n71) );
  INV_X1 U63 ( .A(DIN[28]), .ZN(n297) );
  OAI22_X1 U64 ( .A1(n66), .A2(n263), .B1(n260), .B2(n295), .ZN(n69) );
  INV_X1 U65 ( .A(DIN[30]), .ZN(n295) );
  OAI22_X1 U66 ( .A1(n67), .A2(n263), .B1(n260), .B2(n294), .ZN(n68) );
  INV_X1 U67 ( .A(DIN[31]), .ZN(n294) );
  OAI22_X1 U68 ( .A1(n41), .A2(n265), .B1(n262), .B2(n280), .ZN(n94) );
  INV_X1 U69 ( .A(DIN[5]), .ZN(n280) );
  OAI22_X1 U70 ( .A1(n42), .A2(n265), .B1(n262), .B2(n279), .ZN(n93) );
  INV_X1 U71 ( .A(DIN[6]), .ZN(n279) );
  OAI22_X1 U72 ( .A1(n44), .A2(n265), .B1(n262), .B2(n285), .ZN(n91) );
  INV_X1 U73 ( .A(DIN[8]), .ZN(n285) );
  OAI22_X1 U74 ( .A1(n45), .A2(n264), .B1(n262), .B2(n284), .ZN(n90) );
  INV_X1 U75 ( .A(DIN[9]), .ZN(n284) );
endmodule


module MUX31_GENERIC_NBIT32_3 ( S2, S1, S0, SEL, Y );
  input [31:0] S2;
  input [31:0] S1;
  input [31:0] S0;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n310, n311;

  BUF_X1 U2 ( .A(n37), .Z(n273) );
  BUF_X1 U3 ( .A(n37), .Z(n272) );
  BUF_X1 U4 ( .A(n36), .Z(n276) );
  BUF_X1 U5 ( .A(n36), .Z(n275) );
  BUF_X1 U6 ( .A(n36), .Z(n277) );
  BUF_X1 U7 ( .A(n38), .Z(n270) );
  BUF_X1 U8 ( .A(n38), .Z(n269) );
  BUF_X1 U9 ( .A(n37), .Z(n274) );
  BUF_X1 U10 ( .A(n38), .Z(n271) );
  INV_X1 U11 ( .A(SEL[0]), .ZN(n311) );
  NOR3_X1 U12 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n311), .ZN(n36) );
  NOR3_X1 U13 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n310), .ZN(n37) );
  AND3_X1 U14 ( .A1(n311), .A2(n310), .A3(SEL[2]), .ZN(n38) );
  INV_X1 U15 ( .A(SEL[1]), .ZN(n310) );
  INV_X1 U16 ( .A(n46), .ZN(Y[23]) );
  INV_X1 U17 ( .A(n47), .ZN(Y[22]) );
  INV_X1 U18 ( .A(n48), .ZN(Y[21]) );
  INV_X1 U19 ( .A(n60), .ZN(Y[9]) );
  INV_X1 U20 ( .A(n61), .ZN(Y[8]) );
  INV_X1 U21 ( .A(n62), .ZN(Y[7]) );
  INV_X1 U22 ( .A(n64), .ZN(Y[5]) );
  INV_X1 U23 ( .A(n65), .ZN(Y[4]) );
  INV_X1 U24 ( .A(n66), .ZN(Y[3]) );
  INV_X1 U25 ( .A(n39), .ZN(Y[30]) );
  INV_X1 U26 ( .A(n67), .ZN(Y[2]) );
  INV_X1 U27 ( .A(n40), .ZN(Y[29]) );
  INV_X1 U28 ( .A(n42), .ZN(Y[27]) );
  INV_X1 U29 ( .A(n43), .ZN(Y[26]) );
  INV_X1 U30 ( .A(n44), .ZN(Y[25]) );
  AOI222_X1 U31 ( .A1(S0[21]), .A2(n276), .B1(S1[21]), .B2(n273), .C1(S2[21]), 
        .C2(n270), .ZN(n48) );
  AOI222_X1 U32 ( .A1(S0[22]), .A2(n277), .B1(S1[22]), .B2(n273), .C1(S2[22]), 
        .C2(n270), .ZN(n47) );
  AOI222_X1 U33 ( .A1(S0[23]), .A2(n277), .B1(S1[23]), .B2(n273), .C1(S2[23]), 
        .C2(n270), .ZN(n46) );
  AOI222_X1 U34 ( .A1(S0[3]), .A2(n275), .B1(S1[3]), .B2(n272), .C1(S2[3]), 
        .C2(n269), .ZN(n66) );
  AOI222_X1 U35 ( .A1(S0[4]), .A2(n275), .B1(S1[4]), .B2(n272), .C1(S2[4]), 
        .C2(n269), .ZN(n65) );
  AOI222_X1 U36 ( .A1(S0[5]), .A2(n275), .B1(S1[5]), .B2(n272), .C1(S2[5]), 
        .C2(n269), .ZN(n64) );
  AOI222_X1 U37 ( .A1(S0[7]), .A2(n275), .B1(S1[7]), .B2(n272), .C1(S2[7]), 
        .C2(n269), .ZN(n62) );
  AOI222_X1 U38 ( .A1(S0[8]), .A2(n275), .B1(S1[8]), .B2(n272), .C1(S2[8]), 
        .C2(n269), .ZN(n61) );
  AOI222_X1 U39 ( .A1(S0[9]), .A2(n275), .B1(S1[9]), .B2(n272), .C1(S2[9]), 
        .C2(n269), .ZN(n60) );
  AOI222_X1 U40 ( .A1(S0[2]), .A2(n275), .B1(S1[2]), .B2(n272), .C1(S2[2]), 
        .C2(n269), .ZN(n67) );
  AOI222_X1 U41 ( .A1(S0[29]), .A2(n277), .B1(S1[29]), .B2(n274), .C1(S2[29]), 
        .C2(n271), .ZN(n40) );
  AOI222_X1 U42 ( .A1(S0[30]), .A2(n277), .B1(S1[30]), .B2(n274), .C1(S2[30]), 
        .C2(n271), .ZN(n39) );
  AOI222_X1 U43 ( .A1(S0[25]), .A2(n277), .B1(S1[25]), .B2(n274), .C1(S2[25]), 
        .C2(n271), .ZN(n44) );
  AOI222_X1 U44 ( .A1(S0[26]), .A2(n277), .B1(S1[26]), .B2(n274), .C1(S2[26]), 
        .C2(n271), .ZN(n43) );
  AOI222_X1 U45 ( .A1(S0[27]), .A2(n277), .B1(S1[27]), .B2(n274), .C1(S2[27]), 
        .C2(n271), .ZN(n42) );
  INV_X1 U46 ( .A(n49), .ZN(Y[20]) );
  AOI222_X1 U47 ( .A1(S0[20]), .A2(n276), .B1(S1[20]), .B2(n273), .C1(S2[20]), 
        .C2(n270), .ZN(n49) );
  INV_X1 U48 ( .A(n52), .ZN(Y[17]) );
  AOI222_X1 U49 ( .A1(S0[17]), .A2(n276), .B1(S1[17]), .B2(n273), .C1(S2[17]), 
        .C2(n270), .ZN(n52) );
  INV_X1 U50 ( .A(n56), .ZN(Y[13]) );
  AOI222_X1 U51 ( .A1(S0[13]), .A2(n276), .B1(S1[13]), .B2(n273), .C1(S2[13]), 
        .C2(n270), .ZN(n56) );
  INV_X1 U52 ( .A(n69), .ZN(Y[0]) );
  AOI222_X1 U53 ( .A1(S0[0]), .A2(n275), .B1(S1[0]), .B2(n272), .C1(S2[0]), 
        .C2(n269), .ZN(n69) );
  INV_X1 U54 ( .A(n63), .ZN(Y[6]) );
  AOI222_X1 U55 ( .A1(S0[6]), .A2(n275), .B1(S1[6]), .B2(n272), .C1(S2[6]), 
        .C2(n269), .ZN(n63) );
  INV_X1 U56 ( .A(n35), .ZN(Y[31]) );
  AOI222_X1 U57 ( .A1(S0[31]), .A2(n277), .B1(S1[31]), .B2(n274), .C1(S2[31]), 
        .C2(n271), .ZN(n35) );
  INV_X1 U58 ( .A(n41), .ZN(Y[28]) );
  AOI222_X1 U59 ( .A1(S0[28]), .A2(n277), .B1(S1[28]), .B2(n274), .C1(S2[28]), 
        .C2(n271), .ZN(n41) );
  INV_X1 U60 ( .A(n45), .ZN(Y[24]) );
  AOI222_X1 U61 ( .A1(S0[24]), .A2(n277), .B1(S1[24]), .B2(n274), .C1(S2[24]), 
        .C2(n271), .ZN(n45) );
  INV_X1 U62 ( .A(n51), .ZN(Y[18]) );
  AOI222_X1 U63 ( .A1(S0[18]), .A2(n276), .B1(S1[18]), .B2(n273), .C1(S2[18]), 
        .C2(n270), .ZN(n51) );
  INV_X1 U64 ( .A(n55), .ZN(Y[14]) );
  AOI222_X1 U65 ( .A1(S0[14]), .A2(n276), .B1(S1[14]), .B2(n273), .C1(S2[14]), 
        .C2(n270), .ZN(n55) );
  INV_X1 U66 ( .A(n59), .ZN(Y[10]) );
  AOI222_X1 U67 ( .A1(S0[10]), .A2(n275), .B1(S1[10]), .B2(n272), .C1(S2[10]), 
        .C2(n269), .ZN(n59) );
  INV_X1 U68 ( .A(n50), .ZN(Y[19]) );
  AOI222_X1 U69 ( .A1(S0[19]), .A2(n276), .B1(S1[19]), .B2(n273), .C1(S2[19]), 
        .C2(n270), .ZN(n50) );
  INV_X1 U70 ( .A(n54), .ZN(Y[15]) );
  AOI222_X1 U71 ( .A1(S0[15]), .A2(n276), .B1(S1[15]), .B2(n273), .C1(S2[15]), 
        .C2(n270), .ZN(n54) );
  INV_X1 U72 ( .A(n58), .ZN(Y[11]) );
  AOI222_X1 U73 ( .A1(S0[11]), .A2(n276), .B1(S1[11]), .B2(n272), .C1(S2[11]), 
        .C2(n269), .ZN(n58) );
  INV_X1 U74 ( .A(n68), .ZN(Y[1]) );
  AOI222_X1 U75 ( .A1(S0[1]), .A2(n275), .B1(S1[1]), .B2(n272), .C1(S2[1]), 
        .C2(n269), .ZN(n68) );
  INV_X1 U76 ( .A(n53), .ZN(Y[16]) );
  AOI222_X1 U77 ( .A1(S0[16]), .A2(n276), .B1(S1[16]), .B2(n273), .C1(S2[16]), 
        .C2(n270), .ZN(n53) );
  INV_X1 U78 ( .A(n57), .ZN(Y[12]) );
  AOI222_X1 U79 ( .A1(S0[12]), .A2(n276), .B1(S1[12]), .B2(n273), .C1(S2[12]), 
        .C2(n270), .ZN(n57) );
endmodule


module ZERO_DETECTOR_WIDTH32_0 ( A, Y );
  input [31:0] A;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NOR4_X1 U1 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n6) );
  NOR4_X1 U2 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n10) );
  NOR4_X1 U3 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n9) );
  NOR4_X1 U4 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n8) );
  NOR4_X1 U5 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n7) );
  NAND4_X1 U6 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NOR4_X1 U7 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n3) );
  NOR4_X1 U8 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n4) );
  NOR4_X1 U9 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n5) );
  NOR2_X1 U10 ( .A1(n1), .A2(n2), .ZN(Y) );
  NAND4_X1 U11 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
endmodule


module BRANCH_UNIT_WIDTH32 ( Z, EQ_COND, JUMP_EN, BRANCH );
  input Z, EQ_COND, JUMP_EN;
  output BRANCH;
  wire   n1;

  AND2_X1 U1 ( .A1(n1), .A2(JUMP_EN), .ZN(BRANCH) );
  XNOR2_X1 U2 ( .A(Z), .B(EQ_COND), .ZN(n1) );
endmodule


module REGISTER_GENERIC_WIDTH32_5 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296;

  DFF_X1 \DOUT_reg[31]  ( .D(n68), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[30]  ( .D(n69), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[29]  ( .D(n70), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[28]  ( .D(n71), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[27]  ( .D(n72), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n73), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[25]  ( .D(n74), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[24]  ( .D(n75), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[22]  ( .D(n77), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[21]  ( .D(n78), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[20]  ( .D(n79), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n80), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n81), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n83), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n84), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n89), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n90), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n91), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n92), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n93), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n94), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n95), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n96), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n97), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n98), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n260) );
  BUF_X1 U4 ( .A(n35), .Z(n259) );
  BUF_X1 U5 ( .A(n35), .Z(n258) );
  BUF_X1 U6 ( .A(n34), .Z(n263) );
  NAND2_X1 U7 ( .A1(RST), .A2(n261), .ZN(n35) );
  BUF_X1 U8 ( .A(n34), .Z(n261) );
  BUF_X1 U9 ( .A(n34), .Z(n262) );
  OAI22_X1 U10 ( .A1(n36), .A2(n263), .B1(n260), .B2(n295), .ZN(n99) );
  INV_X1 U11 ( .A(DIN[0]), .ZN(n295) );
  OAI22_X1 U12 ( .A1(n37), .A2(n263), .B1(n260), .B2(n294), .ZN(n98) );
  INV_X1 U13 ( .A(DIN[1]), .ZN(n294) );
  OAI22_X1 U14 ( .A1(n38), .A2(n263), .B1(n260), .B2(n293), .ZN(n97) );
  INV_X1 U15 ( .A(DIN[2]), .ZN(n293) );
  OAI22_X1 U16 ( .A1(n39), .A2(n263), .B1(n260), .B2(n292), .ZN(n96) );
  INV_X1 U17 ( .A(DIN[3]), .ZN(n292) );
  OAI22_X1 U18 ( .A1(n40), .A2(n263), .B1(n260), .B2(n291), .ZN(n95) );
  INV_X1 U19 ( .A(DIN[4]), .ZN(n291) );
  OAI22_X1 U20 ( .A1(n41), .A2(n263), .B1(n260), .B2(n290), .ZN(n94) );
  INV_X1 U21 ( .A(DIN[5]), .ZN(n290) );
  OAI22_X1 U22 ( .A1(n42), .A2(n263), .B1(n260), .B2(n289), .ZN(n93) );
  INV_X1 U23 ( .A(DIN[6]), .ZN(n289) );
  OAI22_X1 U24 ( .A1(n43), .A2(n263), .B1(n260), .B2(n288), .ZN(n92) );
  INV_X1 U25 ( .A(DIN[7]), .ZN(n288) );
  OAI22_X1 U26 ( .A1(n44), .A2(n263), .B1(n260), .B2(n287), .ZN(n91) );
  INV_X1 U27 ( .A(DIN[8]), .ZN(n287) );
  OAI22_X1 U28 ( .A1(n45), .A2(n262), .B1(n260), .B2(n286), .ZN(n90) );
  INV_X1 U29 ( .A(DIN[9]), .ZN(n286) );
  OAI22_X1 U30 ( .A1(n46), .A2(n262), .B1(n259), .B2(n285), .ZN(n89) );
  INV_X1 U31 ( .A(DIN[10]), .ZN(n285) );
  OAI22_X1 U32 ( .A1(n47), .A2(n262), .B1(n259), .B2(n284), .ZN(n88) );
  INV_X1 U33 ( .A(DIN[11]), .ZN(n284) );
  OAI22_X1 U34 ( .A1(n48), .A2(n262), .B1(n259), .B2(n283), .ZN(n87) );
  INV_X1 U35 ( .A(DIN[12]), .ZN(n283) );
  OAI22_X1 U36 ( .A1(n49), .A2(n262), .B1(n259), .B2(n282), .ZN(n86) );
  INV_X1 U37 ( .A(DIN[13]), .ZN(n282) );
  OAI22_X1 U38 ( .A1(n50), .A2(n262), .B1(n259), .B2(n281), .ZN(n85) );
  INV_X1 U39 ( .A(DIN[14]), .ZN(n281) );
  OAI22_X1 U40 ( .A1(n51), .A2(n262), .B1(n259), .B2(n280), .ZN(n84) );
  INV_X1 U41 ( .A(DIN[15]), .ZN(n280) );
  OAI22_X1 U42 ( .A1(n52), .A2(n262), .B1(n259), .B2(n279), .ZN(n83) );
  INV_X1 U43 ( .A(DIN[16]), .ZN(n279) );
  OAI22_X1 U44 ( .A1(n53), .A2(n262), .B1(n259), .B2(n278), .ZN(n82) );
  INV_X1 U45 ( .A(DIN[17]), .ZN(n278) );
  OAI22_X1 U46 ( .A1(n54), .A2(n262), .B1(n259), .B2(n277), .ZN(n81) );
  INV_X1 U47 ( .A(DIN[18]), .ZN(n277) );
  OAI22_X1 U48 ( .A1(n55), .A2(n262), .B1(n259), .B2(n276), .ZN(n80) );
  INV_X1 U49 ( .A(DIN[19]), .ZN(n276) );
  OAI22_X1 U50 ( .A1(n56), .A2(n262), .B1(n259), .B2(n275), .ZN(n79) );
  INV_X1 U51 ( .A(DIN[20]), .ZN(n275) );
  OAI22_X1 U52 ( .A1(n57), .A2(n261), .B1(n258), .B2(n274), .ZN(n78) );
  INV_X1 U53 ( .A(DIN[21]), .ZN(n274) );
  OAI22_X1 U54 ( .A1(n58), .A2(n261), .B1(n258), .B2(n273), .ZN(n77) );
  INV_X1 U55 ( .A(DIN[22]), .ZN(n273) );
  OAI22_X1 U56 ( .A1(n59), .A2(n261), .B1(n258), .B2(n272), .ZN(n76) );
  INV_X1 U57 ( .A(DIN[23]), .ZN(n272) );
  OAI22_X1 U58 ( .A1(n60), .A2(n261), .B1(n258), .B2(n271), .ZN(n75) );
  INV_X1 U59 ( .A(DIN[24]), .ZN(n271) );
  OAI22_X1 U60 ( .A1(n61), .A2(n261), .B1(n258), .B2(n270), .ZN(n74) );
  INV_X1 U61 ( .A(DIN[25]), .ZN(n270) );
  OAI22_X1 U62 ( .A1(n62), .A2(n261), .B1(n258), .B2(n269), .ZN(n73) );
  INV_X1 U63 ( .A(DIN[26]), .ZN(n269) );
  OAI22_X1 U64 ( .A1(n63), .A2(n261), .B1(n258), .B2(n268), .ZN(n72) );
  INV_X1 U65 ( .A(DIN[27]), .ZN(n268) );
  OAI22_X1 U66 ( .A1(n64), .A2(n261), .B1(n258), .B2(n267), .ZN(n71) );
  INV_X1 U67 ( .A(DIN[28]), .ZN(n267) );
  OAI22_X1 U68 ( .A1(n65), .A2(n261), .B1(n258), .B2(n266), .ZN(n70) );
  INV_X1 U69 ( .A(DIN[29]), .ZN(n266) );
  OAI22_X1 U70 ( .A1(n66), .A2(n261), .B1(n258), .B2(n265), .ZN(n69) );
  INV_X1 U71 ( .A(DIN[30]), .ZN(n265) );
  OAI22_X1 U72 ( .A1(n67), .A2(n261), .B1(n258), .B2(n264), .ZN(n68) );
  INV_X1 U73 ( .A(DIN[31]), .ZN(n264) );
  NAND2_X1 U74 ( .A1(n296), .A2(RST), .ZN(n34) );
  INV_X1 U75 ( .A(EN), .ZN(n296) );
endmodule


module REGISTER_GENERIC_WIDTH5_2 ( CLK, RST, EN, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST, EN;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n44, n45, n46, n47,
         n48, n49, n50, n51;

  DFF_X1 \DOUT_reg[4]  ( .D(n14), .CK(CLK), .Q(DOUT[4]), .QN(n13) );
  DFF_X1 \DOUT_reg[3]  ( .D(n15), .CK(CLK), .Q(DOUT[3]), .QN(n12) );
  DFF_X1 \DOUT_reg[2]  ( .D(n16), .CK(CLK), .Q(DOUT[2]), .QN(n11) );
  DFF_X1 \DOUT_reg[1]  ( .D(n17), .CK(CLK), .Q(DOUT[1]), .QN(n10) );
  DFF_X1 \DOUT_reg[0]  ( .D(n18), .CK(CLK), .Q(DOUT[0]), .QN(n9) );
  AND2_X1 U3 ( .A1(RST), .A2(n51), .ZN(n49) );
  NAND2_X1 U4 ( .A1(n44), .A2(RST), .ZN(n51) );
  INV_X1 U5 ( .A(EN), .ZN(n44) );
  OAI21_X1 U6 ( .B1(n9), .B2(n51), .A(n50), .ZN(n18) );
  NAND2_X1 U7 ( .A1(DIN[0]), .A2(n49), .ZN(n50) );
  OAI21_X1 U8 ( .B1(n10), .B2(n51), .A(n48), .ZN(n17) );
  NAND2_X1 U9 ( .A1(DIN[1]), .A2(n49), .ZN(n48) );
  OAI21_X1 U10 ( .B1(n11), .B2(n51), .A(n47), .ZN(n16) );
  NAND2_X1 U11 ( .A1(DIN[2]), .A2(n49), .ZN(n47) );
  OAI21_X1 U12 ( .B1(n12), .B2(n51), .A(n46), .ZN(n15) );
  NAND2_X1 U13 ( .A1(DIN[3]), .A2(n49), .ZN(n46) );
  OAI21_X1 U14 ( .B1(n13), .B2(n51), .A(n45), .ZN(n14) );
  NAND2_X1 U15 ( .A1(DIN[4]), .A2(n49), .ZN(n45) );
endmodule


module REGISTER_GENERIC_WIDTH32_4 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296;

  DFF_X1 \DOUT_reg[31]  ( .D(n68), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[30]  ( .D(n69), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[29]  ( .D(n70), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[28]  ( .D(n71), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[27]  ( .D(n72), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n73), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[25]  ( .D(n74), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[24]  ( .D(n75), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[22]  ( .D(n77), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[21]  ( .D(n78), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[20]  ( .D(n79), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n80), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n81), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n83), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n84), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n89), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n90), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n91), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n92), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n93), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n94), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n95), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n96), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n97), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n98), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n260) );
  BUF_X1 U4 ( .A(n35), .Z(n259) );
  BUF_X1 U5 ( .A(n35), .Z(n258) );
  BUF_X1 U6 ( .A(n34), .Z(n263) );
  NAND2_X1 U7 ( .A1(RST), .A2(n261), .ZN(n35) );
  BUF_X1 U8 ( .A(n34), .Z(n261) );
  BUF_X1 U9 ( .A(n34), .Z(n262) );
  OAI22_X1 U10 ( .A1(n36), .A2(n263), .B1(n260), .B2(n295), .ZN(n99) );
  INV_X1 U11 ( .A(DIN[0]), .ZN(n295) );
  OAI22_X1 U12 ( .A1(n37), .A2(n263), .B1(n260), .B2(n294), .ZN(n98) );
  INV_X1 U13 ( .A(DIN[1]), .ZN(n294) );
  OAI22_X1 U14 ( .A1(n38), .A2(n263), .B1(n260), .B2(n293), .ZN(n97) );
  INV_X1 U15 ( .A(DIN[2]), .ZN(n293) );
  OAI22_X1 U16 ( .A1(n39), .A2(n263), .B1(n260), .B2(n292), .ZN(n96) );
  INV_X1 U17 ( .A(DIN[3]), .ZN(n292) );
  OAI22_X1 U18 ( .A1(n40), .A2(n263), .B1(n260), .B2(n291), .ZN(n95) );
  INV_X1 U19 ( .A(DIN[4]), .ZN(n291) );
  OAI22_X1 U20 ( .A1(n41), .A2(n263), .B1(n260), .B2(n290), .ZN(n94) );
  INV_X1 U21 ( .A(DIN[5]), .ZN(n290) );
  OAI22_X1 U22 ( .A1(n42), .A2(n263), .B1(n260), .B2(n289), .ZN(n93) );
  INV_X1 U23 ( .A(DIN[6]), .ZN(n289) );
  OAI22_X1 U24 ( .A1(n43), .A2(n263), .B1(n260), .B2(n288), .ZN(n92) );
  INV_X1 U25 ( .A(DIN[7]), .ZN(n288) );
  OAI22_X1 U26 ( .A1(n44), .A2(n263), .B1(n260), .B2(n287), .ZN(n91) );
  INV_X1 U27 ( .A(DIN[8]), .ZN(n287) );
  OAI22_X1 U28 ( .A1(n45), .A2(n262), .B1(n260), .B2(n286), .ZN(n90) );
  INV_X1 U29 ( .A(DIN[9]), .ZN(n286) );
  OAI22_X1 U30 ( .A1(n46), .A2(n262), .B1(n259), .B2(n285), .ZN(n89) );
  INV_X1 U31 ( .A(DIN[10]), .ZN(n285) );
  OAI22_X1 U32 ( .A1(n47), .A2(n262), .B1(n259), .B2(n284), .ZN(n88) );
  INV_X1 U33 ( .A(DIN[11]), .ZN(n284) );
  OAI22_X1 U34 ( .A1(n48), .A2(n262), .B1(n259), .B2(n283), .ZN(n87) );
  INV_X1 U35 ( .A(DIN[12]), .ZN(n283) );
  OAI22_X1 U36 ( .A1(n49), .A2(n262), .B1(n259), .B2(n282), .ZN(n86) );
  INV_X1 U37 ( .A(DIN[13]), .ZN(n282) );
  OAI22_X1 U38 ( .A1(n50), .A2(n262), .B1(n259), .B2(n281), .ZN(n85) );
  INV_X1 U39 ( .A(DIN[14]), .ZN(n281) );
  OAI22_X1 U40 ( .A1(n51), .A2(n262), .B1(n259), .B2(n280), .ZN(n84) );
  INV_X1 U41 ( .A(DIN[15]), .ZN(n280) );
  OAI22_X1 U42 ( .A1(n52), .A2(n262), .B1(n259), .B2(n279), .ZN(n83) );
  INV_X1 U43 ( .A(DIN[16]), .ZN(n279) );
  OAI22_X1 U44 ( .A1(n53), .A2(n262), .B1(n259), .B2(n278), .ZN(n82) );
  INV_X1 U45 ( .A(DIN[17]), .ZN(n278) );
  OAI22_X1 U46 ( .A1(n54), .A2(n262), .B1(n259), .B2(n277), .ZN(n81) );
  INV_X1 U47 ( .A(DIN[18]), .ZN(n277) );
  OAI22_X1 U48 ( .A1(n55), .A2(n262), .B1(n259), .B2(n276), .ZN(n80) );
  INV_X1 U49 ( .A(DIN[19]), .ZN(n276) );
  OAI22_X1 U50 ( .A1(n56), .A2(n262), .B1(n259), .B2(n275), .ZN(n79) );
  INV_X1 U51 ( .A(DIN[20]), .ZN(n275) );
  OAI22_X1 U52 ( .A1(n57), .A2(n261), .B1(n258), .B2(n274), .ZN(n78) );
  INV_X1 U53 ( .A(DIN[21]), .ZN(n274) );
  OAI22_X1 U54 ( .A1(n58), .A2(n261), .B1(n258), .B2(n273), .ZN(n77) );
  INV_X1 U55 ( .A(DIN[22]), .ZN(n273) );
  OAI22_X1 U56 ( .A1(n59), .A2(n261), .B1(n258), .B2(n272), .ZN(n76) );
  INV_X1 U57 ( .A(DIN[23]), .ZN(n272) );
  OAI22_X1 U58 ( .A1(n60), .A2(n261), .B1(n258), .B2(n271), .ZN(n75) );
  INV_X1 U59 ( .A(DIN[24]), .ZN(n271) );
  OAI22_X1 U60 ( .A1(n61), .A2(n261), .B1(n258), .B2(n270), .ZN(n74) );
  INV_X1 U61 ( .A(DIN[25]), .ZN(n270) );
  OAI22_X1 U62 ( .A1(n62), .A2(n261), .B1(n258), .B2(n269), .ZN(n73) );
  INV_X1 U63 ( .A(DIN[26]), .ZN(n269) );
  OAI22_X1 U64 ( .A1(n63), .A2(n261), .B1(n258), .B2(n268), .ZN(n72) );
  INV_X1 U65 ( .A(DIN[27]), .ZN(n268) );
  OAI22_X1 U66 ( .A1(n64), .A2(n261), .B1(n258), .B2(n267), .ZN(n71) );
  INV_X1 U67 ( .A(DIN[28]), .ZN(n267) );
  OAI22_X1 U68 ( .A1(n65), .A2(n261), .B1(n258), .B2(n266), .ZN(n70) );
  INV_X1 U69 ( .A(DIN[29]), .ZN(n266) );
  OAI22_X1 U70 ( .A1(n66), .A2(n261), .B1(n258), .B2(n265), .ZN(n69) );
  INV_X1 U71 ( .A(DIN[30]), .ZN(n265) );
  OAI22_X1 U72 ( .A1(n67), .A2(n261), .B1(n258), .B2(n264), .ZN(n68) );
  INV_X1 U73 ( .A(DIN[31]), .ZN(n264) );
  NAND2_X1 U74 ( .A1(n296), .A2(RST), .ZN(n34) );
  INV_X1 U75 ( .A(EN), .ZN(n296) );
endmodule


module SIGN_EXTEND_WIDTH_IN8_WIDTH_OUT32_0 ( A, S, Y );
  input [7:0] A;
  output [31:0] Y;
  input S;
  wire   N0, \Y[31] , \Y[19] ;
  assign Y[7] = A[7];
  assign Y[6] = A[6];
  assign Y[5] = A[5];
  assign Y[4] = A[4];
  assign Y[3] = A[3];
  assign Y[2] = A[2];
  assign Y[1] = A[1];
  assign Y[0] = A[0];
  assign Y[20] = \Y[31] ;
  assign Y[21] = \Y[31] ;
  assign Y[22] = \Y[31] ;
  assign Y[23] = \Y[31] ;
  assign Y[24] = \Y[31] ;
  assign Y[25] = \Y[31] ;
  assign Y[26] = \Y[31] ;
  assign Y[27] = \Y[31] ;
  assign Y[28] = \Y[31] ;
  assign Y[29] = \Y[31] ;
  assign Y[30] = \Y[31] ;
  assign Y[31] = \Y[31] ;
  assign Y[8] = \Y[19] ;
  assign Y[9] = \Y[19] ;
  assign Y[10] = \Y[19] ;
  assign Y[11] = \Y[19] ;
  assign Y[12] = \Y[19] ;
  assign Y[13] = \Y[19] ;
  assign Y[14] = \Y[19] ;
  assign Y[15] = \Y[19] ;
  assign Y[16] = \Y[19] ;
  assign Y[17] = \Y[19] ;
  assign Y[18] = \Y[19] ;
  assign Y[19] = \Y[19] ;

  BUF_X1 U1 ( .A(N0), .Z(\Y[19] ) );
  BUF_X1 U2 ( .A(N0), .Z(\Y[31] ) );
  AND2_X1 U3 ( .A1(S), .A2(A[7]), .ZN(N0) );
endmodule


module SIGN_EXTEND_WIDTH_IN16_WIDTH_OUT32_2 ( A, S, Y );
  input [15:0] A;
  output [31:0] Y;
  input S;
  wire   N0;
  assign Y[15] = A[15];
  assign Y[14] = A[14];
  assign Y[13] = A[13];
  assign Y[12] = A[12];
  assign Y[11] = A[11];
  assign Y[10] = A[10];
  assign Y[9] = A[9];
  assign Y[8] = A[8];
  assign Y[7] = A[7];
  assign Y[6] = A[6];
  assign Y[5] = A[5];
  assign Y[4] = A[4];
  assign Y[3] = A[3];
  assign Y[2] = A[2];
  assign Y[1] = A[1];
  assign Y[0] = A[0];
  assign Y[16] = N0;
  assign Y[17] = N0;
  assign Y[18] = N0;
  assign Y[19] = N0;
  assign Y[20] = N0;
  assign Y[21] = N0;
  assign Y[22] = N0;
  assign Y[23] = N0;
  assign Y[24] = N0;
  assign Y[25] = N0;
  assign Y[26] = N0;
  assign Y[27] = N0;
  assign Y[28] = N0;
  assign Y[29] = N0;
  assign Y[30] = N0;
  assign Y[31] = N0;

  AND2_X1 U1 ( .A1(S), .A2(A[15]), .ZN(N0) );
endmodule


module MUX31_GENERIC_NBIT32_2 ( S2, S1, S0, SEL, Y );
  input [31:0] S2;
  input [31:0] S1;
  input [31:0] S0;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n285, n286;

  BUF_X1 U2 ( .A(n37), .Z(n247) );
  BUF_X1 U3 ( .A(n37), .Z(n248) );
  BUF_X1 U4 ( .A(n36), .Z(n250) );
  BUF_X1 U5 ( .A(n36), .Z(n251) );
  BUF_X1 U6 ( .A(n36), .Z(n252) );
  BUF_X1 U7 ( .A(n38), .Z(n244) );
  BUF_X1 U8 ( .A(n38), .Z(n245) );
  BUF_X1 U9 ( .A(n37), .Z(n249) );
  BUF_X1 U10 ( .A(n38), .Z(n246) );
  NOR3_X1 U11 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n285), .ZN(n37) );
  NOR3_X1 U12 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n286), .ZN(n36) );
  INV_X1 U13 ( .A(n69), .ZN(Y[0]) );
  AOI222_X1 U14 ( .A1(S0[0]), .A2(n250), .B1(S1[0]), .B2(n247), .C1(S2[0]), 
        .C2(n244), .ZN(n69) );
  INV_X1 U15 ( .A(n68), .ZN(Y[1]) );
  AOI222_X1 U16 ( .A1(S0[1]), .A2(n250), .B1(S1[1]), .B2(n247), .C1(S2[1]), 
        .C2(n244), .ZN(n68) );
  INV_X1 U17 ( .A(n67), .ZN(Y[2]) );
  AOI222_X1 U18 ( .A1(S0[2]), .A2(n250), .B1(S1[2]), .B2(n247), .C1(S2[2]), 
        .C2(n244), .ZN(n67) );
  INV_X1 U19 ( .A(n66), .ZN(Y[3]) );
  AOI222_X1 U20 ( .A1(S0[3]), .A2(n250), .B1(S1[3]), .B2(n247), .C1(S2[3]), 
        .C2(n244), .ZN(n66) );
  INV_X1 U21 ( .A(n65), .ZN(Y[4]) );
  AOI222_X1 U22 ( .A1(S0[4]), .A2(n250), .B1(S1[4]), .B2(n247), .C1(S2[4]), 
        .C2(n244), .ZN(n65) );
  INV_X1 U23 ( .A(n64), .ZN(Y[5]) );
  AOI222_X1 U24 ( .A1(S0[5]), .A2(n250), .B1(S1[5]), .B2(n247), .C1(S2[5]), 
        .C2(n244), .ZN(n64) );
  INV_X1 U25 ( .A(n63), .ZN(Y[6]) );
  AOI222_X1 U26 ( .A1(S0[6]), .A2(n250), .B1(S1[6]), .B2(n247), .C1(S2[6]), 
        .C2(n244), .ZN(n63) );
  INV_X1 U27 ( .A(n62), .ZN(Y[7]) );
  AOI222_X1 U28 ( .A1(S0[7]), .A2(n250), .B1(S1[7]), .B2(n247), .C1(S2[7]), 
        .C2(n244), .ZN(n62) );
  INV_X1 U29 ( .A(n61), .ZN(Y[8]) );
  AOI222_X1 U30 ( .A1(S0[8]), .A2(n250), .B1(S1[8]), .B2(n247), .C1(S2[8]), 
        .C2(n244), .ZN(n61) );
  INV_X1 U31 ( .A(n60), .ZN(Y[9]) );
  AOI222_X1 U32 ( .A1(S0[9]), .A2(n250), .B1(S1[9]), .B2(n247), .C1(S2[9]), 
        .C2(n244), .ZN(n60) );
  INV_X1 U33 ( .A(n59), .ZN(Y[10]) );
  AOI222_X1 U34 ( .A1(S0[10]), .A2(n250), .B1(S1[10]), .B2(n247), .C1(S2[10]), 
        .C2(n244), .ZN(n59) );
  INV_X1 U35 ( .A(n58), .ZN(Y[11]) );
  AOI222_X1 U36 ( .A1(S0[11]), .A2(n251), .B1(S1[11]), .B2(n247), .C1(S2[11]), 
        .C2(n244), .ZN(n58) );
  INV_X1 U37 ( .A(n57), .ZN(Y[12]) );
  AOI222_X1 U38 ( .A1(S0[12]), .A2(n251), .B1(S1[12]), .B2(n248), .C1(S2[12]), 
        .C2(n245), .ZN(n57) );
  INV_X1 U39 ( .A(n56), .ZN(Y[13]) );
  AOI222_X1 U40 ( .A1(S0[13]), .A2(n251), .B1(S1[13]), .B2(n248), .C1(S2[13]), 
        .C2(n245), .ZN(n56) );
  INV_X1 U41 ( .A(n55), .ZN(Y[14]) );
  AOI222_X1 U42 ( .A1(S0[14]), .A2(n251), .B1(S1[14]), .B2(n248), .C1(S2[14]), 
        .C2(n245), .ZN(n55) );
  INV_X1 U43 ( .A(n54), .ZN(Y[15]) );
  AOI222_X1 U44 ( .A1(S0[15]), .A2(n251), .B1(S1[15]), .B2(n248), .C1(S2[15]), 
        .C2(n245), .ZN(n54) );
  INV_X1 U45 ( .A(n53), .ZN(Y[16]) );
  AOI222_X1 U46 ( .A1(S0[16]), .A2(n251), .B1(S1[16]), .B2(n248), .C1(S2[16]), 
        .C2(n245), .ZN(n53) );
  INV_X1 U47 ( .A(n52), .ZN(Y[17]) );
  AOI222_X1 U48 ( .A1(S0[17]), .A2(n251), .B1(S1[17]), .B2(n248), .C1(S2[17]), 
        .C2(n245), .ZN(n52) );
  INV_X1 U49 ( .A(n51), .ZN(Y[18]) );
  AOI222_X1 U50 ( .A1(S0[18]), .A2(n251), .B1(S1[18]), .B2(n248), .C1(S2[18]), 
        .C2(n245), .ZN(n51) );
  INV_X1 U51 ( .A(n50), .ZN(Y[19]) );
  AOI222_X1 U52 ( .A1(S0[19]), .A2(n251), .B1(S1[19]), .B2(n248), .C1(S2[19]), 
        .C2(n245), .ZN(n50) );
  INV_X1 U53 ( .A(n49), .ZN(Y[20]) );
  AOI222_X1 U54 ( .A1(S0[20]), .A2(n251), .B1(S1[20]), .B2(n248), .C1(S2[20]), 
        .C2(n245), .ZN(n49) );
  INV_X1 U55 ( .A(n48), .ZN(Y[21]) );
  AOI222_X1 U56 ( .A1(S0[21]), .A2(n251), .B1(S1[21]), .B2(n248), .C1(S2[21]), 
        .C2(n245), .ZN(n48) );
  INV_X1 U57 ( .A(n47), .ZN(Y[22]) );
  AOI222_X1 U58 ( .A1(S0[22]), .A2(n252), .B1(S1[22]), .B2(n248), .C1(S2[22]), 
        .C2(n245), .ZN(n47) );
  INV_X1 U59 ( .A(n46), .ZN(Y[23]) );
  AOI222_X1 U60 ( .A1(S0[23]), .A2(n252), .B1(S1[23]), .B2(n248), .C1(S2[23]), 
        .C2(n245), .ZN(n46) );
  AND3_X1 U61 ( .A1(n286), .A2(n285), .A3(SEL[2]), .ZN(n38) );
  INV_X1 U62 ( .A(n35), .ZN(Y[31]) );
  AOI222_X1 U63 ( .A1(S0[31]), .A2(n252), .B1(S1[31]), .B2(n249), .C1(S2[31]), 
        .C2(n246), .ZN(n35) );
  INV_X1 U64 ( .A(n45), .ZN(Y[24]) );
  AOI222_X1 U65 ( .A1(S0[24]), .A2(n252), .B1(S1[24]), .B2(n249), .C1(S2[24]), 
        .C2(n246), .ZN(n45) );
  INV_X1 U66 ( .A(n44), .ZN(Y[25]) );
  AOI222_X1 U67 ( .A1(S0[25]), .A2(n252), .B1(S1[25]), .B2(n249), .C1(S2[25]), 
        .C2(n246), .ZN(n44) );
  INV_X1 U68 ( .A(n43), .ZN(Y[26]) );
  AOI222_X1 U69 ( .A1(S0[26]), .A2(n252), .B1(S1[26]), .B2(n249), .C1(S2[26]), 
        .C2(n246), .ZN(n43) );
  INV_X1 U70 ( .A(n42), .ZN(Y[27]) );
  AOI222_X1 U71 ( .A1(S0[27]), .A2(n252), .B1(S1[27]), .B2(n249), .C1(S2[27]), 
        .C2(n246), .ZN(n42) );
  INV_X1 U72 ( .A(n41), .ZN(Y[28]) );
  AOI222_X1 U73 ( .A1(S0[28]), .A2(n252), .B1(S1[28]), .B2(n249), .C1(S2[28]), 
        .C2(n246), .ZN(n41) );
  INV_X1 U74 ( .A(n40), .ZN(Y[29]) );
  AOI222_X1 U75 ( .A1(S0[29]), .A2(n252), .B1(S1[29]), .B2(n249), .C1(S2[29]), 
        .C2(n246), .ZN(n40) );
  INV_X1 U76 ( .A(n39), .ZN(Y[30]) );
  AOI222_X1 U77 ( .A1(S0[30]), .A2(n252), .B1(S1[30]), .B2(n249), .C1(S2[30]), 
        .C2(n246), .ZN(n39) );
  INV_X1 U78 ( .A(SEL[1]), .ZN(n285) );
  INV_X1 U79 ( .A(SEL[0]), .ZN(n286) );
endmodule


module MUX21_GENERIC_NBIT32_3 ( S1, S0, SEL, Y );
  input [31:0] S1;
  input [31:0] S0;
  output [31:0] Y;
  input SEL;
  wire   net77337, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266;
  assign net77337 = SEL;

  INV_X1 U1 ( .A(n266), .ZN(n257) );
  INV_X1 U2 ( .A(n266), .ZN(n256) );
  BUF_X1 U3 ( .A(n254), .Z(n261) );
  BUF_X1 U4 ( .A(n253), .Z(n258) );
  BUF_X1 U5 ( .A(n253), .Z(n260) );
  BUF_X1 U6 ( .A(n254), .Z(n262) );
  BUF_X1 U7 ( .A(n253), .Z(n259) );
  BUF_X1 U8 ( .A(n255), .Z(n264) );
  BUF_X1 U9 ( .A(n254), .Z(n263) );
  BUF_X1 U10 ( .A(n255), .Z(n266) );
  BUF_X1 U11 ( .A(n255), .Z(n265) );
  BUF_X1 U12 ( .A(net77337), .Z(n255) );
  BUF_X1 U13 ( .A(net77337), .Z(n253) );
  BUF_X1 U14 ( .A(net77337), .Z(n254) );
  INV_X1 U15 ( .A(n49), .ZN(Y[16]) );
  AOI22_X1 U16 ( .A1(S0[16]), .A2(n257), .B1(S1[16]), .B2(n261), .ZN(n49) );
  INV_X1 U17 ( .A(n51), .ZN(Y[14]) );
  AOI22_X1 U18 ( .A1(S0[14]), .A2(n257), .B1(S1[14]), .B2(n261), .ZN(n51) );
  INV_X1 U19 ( .A(n55), .ZN(Y[10]) );
  AOI22_X1 U20 ( .A1(S0[10]), .A2(n256), .B1(S1[10]), .B2(n263), .ZN(n55) );
  INV_X1 U21 ( .A(n46), .ZN(Y[19]) );
  AOI22_X1 U22 ( .A1(S0[19]), .A2(n257), .B1(S1[19]), .B2(n260), .ZN(n46) );
  INV_X1 U23 ( .A(n48), .ZN(Y[17]) );
  AOI22_X1 U24 ( .A1(S0[17]), .A2(n257), .B1(S1[17]), .B2(n261), .ZN(n48) );
  INV_X1 U25 ( .A(n53), .ZN(Y[12]) );
  AOI22_X1 U26 ( .A1(S0[12]), .A2(n257), .B1(S1[12]), .B2(n262), .ZN(n53) );
  INV_X1 U27 ( .A(n50), .ZN(Y[15]) );
  AOI22_X1 U28 ( .A1(S0[15]), .A2(n257), .B1(S1[15]), .B2(n261), .ZN(n50) );
  INV_X1 U29 ( .A(n47), .ZN(Y[18]) );
  AOI22_X1 U30 ( .A1(S0[18]), .A2(n257), .B1(S1[18]), .B2(n260), .ZN(n47) );
  INV_X1 U31 ( .A(n65), .ZN(Y[0]) );
  AOI22_X1 U32 ( .A1(S0[0]), .A2(n256), .B1(S1[0]), .B2(n265), .ZN(n65) );
  INV_X1 U33 ( .A(n54), .ZN(Y[11]) );
  AOI22_X1 U34 ( .A1(S0[11]), .A2(n256), .B1(S1[11]), .B2(n262), .ZN(n54) );
  INV_X1 U35 ( .A(n61), .ZN(Y[4]) );
  AOI22_X1 U36 ( .A1(S0[4]), .A2(n256), .B1(S1[4]), .B2(n264), .ZN(n61) );
  INV_X1 U37 ( .A(n44), .ZN(Y[21]) );
  AOI22_X1 U38 ( .A1(S0[21]), .A2(n257), .B1(S1[21]), .B2(n260), .ZN(n44) );
  INV_X1 U39 ( .A(n43), .ZN(Y[22]) );
  AOI22_X1 U40 ( .A1(S0[22]), .A2(n257), .B1(S1[22]), .B2(n259), .ZN(n43) );
  INV_X1 U41 ( .A(n56), .ZN(Y[9]) );
  AOI22_X1 U42 ( .A1(S0[9]), .A2(n256), .B1(S1[9]), .B2(n263), .ZN(n56) );
  INV_X1 U43 ( .A(n60), .ZN(Y[5]) );
  AOI22_X1 U44 ( .A1(S0[5]), .A2(n256), .B1(S1[5]), .B2(n264), .ZN(n60) );
  INV_X1 U45 ( .A(n64), .ZN(Y[1]) );
  AOI22_X1 U46 ( .A1(S0[1]), .A2(n256), .B1(S1[1]), .B2(n265), .ZN(n64) );
  INV_X1 U47 ( .A(n63), .ZN(Y[2]) );
  AOI22_X1 U48 ( .A1(S0[2]), .A2(n256), .B1(S1[2]), .B2(n265), .ZN(n63) );
  INV_X1 U49 ( .A(n52), .ZN(Y[13]) );
  AOI22_X1 U50 ( .A1(S0[13]), .A2(n257), .B1(S1[13]), .B2(n262), .ZN(n52) );
  INV_X1 U51 ( .A(n42), .ZN(Y[23]) );
  AOI22_X1 U52 ( .A1(S0[23]), .A2(n257), .B1(S1[23]), .B2(n262), .ZN(n42) );
  INV_X1 U53 ( .A(n45), .ZN(Y[20]) );
  AOI22_X1 U54 ( .A1(S0[20]), .A2(n257), .B1(S1[20]), .B2(n260), .ZN(n45) );
  INV_X1 U55 ( .A(n57), .ZN(Y[8]) );
  AOI22_X1 U56 ( .A1(S0[8]), .A2(n256), .B1(S1[8]), .B2(n263), .ZN(n57) );
  INV_X1 U57 ( .A(n62), .ZN(Y[3]) );
  AOI22_X1 U58 ( .A1(S0[3]), .A2(n256), .B1(S1[3]), .B2(n264), .ZN(n62) );
  INV_X1 U59 ( .A(n59), .ZN(Y[6]) );
  AOI22_X1 U60 ( .A1(S0[6]), .A2(n256), .B1(S1[6]), .B2(n264), .ZN(n59) );
  INV_X1 U61 ( .A(n58), .ZN(Y[7]) );
  AOI22_X1 U62 ( .A1(S0[7]), .A2(n256), .B1(S1[7]), .B2(n263), .ZN(n58) );
  INV_X1 U63 ( .A(n39), .ZN(Y[26]) );
  AOI22_X1 U64 ( .A1(S0[26]), .A2(n257), .B1(S1[26]), .B2(n259), .ZN(n39) );
  INV_X1 U65 ( .A(n37), .ZN(Y[28]) );
  AOI22_X1 U66 ( .A1(S0[28]), .A2(n256), .B1(S1[28]), .B2(n258), .ZN(n37) );
  INV_X1 U67 ( .A(n35), .ZN(Y[30]) );
  AOI22_X1 U68 ( .A1(S0[30]), .A2(n257), .B1(S1[30]), .B2(n258), .ZN(n35) );
  INV_X1 U69 ( .A(n41), .ZN(Y[24]) );
  AOI22_X1 U70 ( .A1(S0[24]), .A2(n257), .B1(S1[24]), .B2(n259), .ZN(n41) );
  INV_X1 U71 ( .A(n36), .ZN(Y[29]) );
  AOI22_X1 U72 ( .A1(S0[29]), .A2(n256), .B1(S1[29]), .B2(n258), .ZN(n36) );
  INV_X1 U73 ( .A(n38), .ZN(Y[27]) );
  AOI22_X1 U74 ( .A1(S0[27]), .A2(n257), .B1(S1[27]), .B2(n258), .ZN(n38) );
  INV_X1 U75 ( .A(n40), .ZN(Y[25]) );
  AOI22_X1 U76 ( .A1(S0[25]), .A2(n256), .B1(S1[25]), .B2(n259), .ZN(n40) );
  INV_X1 U77 ( .A(n34), .ZN(Y[31]) );
  AOI22_X1 U78 ( .A1(S0[31]), .A2(n256), .B1(n265), .B2(S1[31]), .ZN(n34) );
endmodule


module MUX21_GENERIC_NBIT32_2 ( S1, S0, SEL, Y );
  input [31:0] S1;
  input [31:0] S0;
  output [31:0] Y;
  input SEL;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294;

  INV_X1 U1 ( .A(n294), .ZN(n284) );
  INV_X1 U2 ( .A(n294), .ZN(n285) );
  BUF_X1 U3 ( .A(n283), .Z(n292) );
  BUF_X1 U4 ( .A(n282), .Z(n291) );
  BUF_X1 U5 ( .A(n282), .Z(n289) );
  BUF_X1 U6 ( .A(n281), .Z(n288) );
  BUF_X1 U7 ( .A(n282), .Z(n290) );
  BUF_X1 U8 ( .A(n281), .Z(n287) );
  BUF_X1 U9 ( .A(n281), .Z(n286) );
  BUF_X1 U10 ( .A(n283), .Z(n294) );
  BUF_X1 U11 ( .A(n283), .Z(n293) );
  BUF_X1 U12 ( .A(SEL), .Z(n283) );
  BUF_X1 U13 ( .A(SEL), .Z(n282) );
  BUF_X1 U14 ( .A(SEL), .Z(n281) );
  INV_X1 U15 ( .A(n34), .ZN(Y[31]) );
  AOI22_X1 U16 ( .A1(S0[31]), .A2(n284), .B1(n293), .B2(S1[31]), .ZN(n34) );
  INV_X1 U17 ( .A(n41), .ZN(Y[24]) );
  AOI22_X1 U18 ( .A1(S0[24]), .A2(n285), .B1(S1[24]), .B2(n287), .ZN(n41) );
  INV_X1 U19 ( .A(n40), .ZN(Y[25]) );
  AOI22_X1 U20 ( .A1(S0[25]), .A2(n284), .B1(S1[25]), .B2(n287), .ZN(n40) );
  INV_X1 U21 ( .A(n39), .ZN(Y[26]) );
  AOI22_X1 U22 ( .A1(S0[26]), .A2(n285), .B1(S1[26]), .B2(n287), .ZN(n39) );
  INV_X1 U23 ( .A(n38), .ZN(Y[27]) );
  AOI22_X1 U24 ( .A1(S0[27]), .A2(n284), .B1(S1[27]), .B2(n286), .ZN(n38) );
  INV_X1 U25 ( .A(n37), .ZN(Y[28]) );
  AOI22_X1 U26 ( .A1(S0[28]), .A2(n285), .B1(S1[28]), .B2(n286), .ZN(n37) );
  INV_X1 U27 ( .A(n36), .ZN(Y[29]) );
  AOI22_X1 U28 ( .A1(S0[29]), .A2(n284), .B1(S1[29]), .B2(n286), .ZN(n36) );
  INV_X1 U29 ( .A(n35), .ZN(Y[30]) );
  AOI22_X1 U30 ( .A1(S0[30]), .A2(n285), .B1(S1[30]), .B2(n286), .ZN(n35) );
  INV_X1 U31 ( .A(n49), .ZN(Y[16]) );
  AOI22_X1 U32 ( .A1(S0[16]), .A2(n285), .B1(S1[16]), .B2(n289), .ZN(n49) );
  INV_X1 U33 ( .A(n48), .ZN(Y[17]) );
  AOI22_X1 U34 ( .A1(S0[17]), .A2(n285), .B1(S1[17]), .B2(n289), .ZN(n48) );
  INV_X1 U35 ( .A(n47), .ZN(Y[18]) );
  AOI22_X1 U36 ( .A1(S0[18]), .A2(n285), .B1(S1[18]), .B2(n288), .ZN(n47) );
  INV_X1 U37 ( .A(n46), .ZN(Y[19]) );
  AOI22_X1 U38 ( .A1(S0[19]), .A2(n285), .B1(S1[19]), .B2(n288), .ZN(n46) );
  INV_X1 U39 ( .A(n45), .ZN(Y[20]) );
  AOI22_X1 U40 ( .A1(S0[20]), .A2(n285), .B1(S1[20]), .B2(n288), .ZN(n45) );
  INV_X1 U41 ( .A(n44), .ZN(Y[21]) );
  AOI22_X1 U42 ( .A1(S0[21]), .A2(n285), .B1(S1[21]), .B2(n288), .ZN(n44) );
  INV_X1 U43 ( .A(n43), .ZN(Y[22]) );
  AOI22_X1 U44 ( .A1(S0[22]), .A2(n285), .B1(S1[22]), .B2(n287), .ZN(n43) );
  INV_X1 U45 ( .A(n42), .ZN(Y[23]) );
  AOI22_X1 U46 ( .A1(S0[23]), .A2(n285), .B1(S1[23]), .B2(n290), .ZN(n42) );
  INV_X1 U47 ( .A(n65), .ZN(Y[0]) );
  AOI22_X1 U48 ( .A1(S0[0]), .A2(n284), .B1(S1[0]), .B2(n293), .ZN(n65) );
  INV_X1 U49 ( .A(n64), .ZN(Y[1]) );
  AOI22_X1 U50 ( .A1(S0[1]), .A2(n284), .B1(S1[1]), .B2(n293), .ZN(n64) );
  INV_X1 U51 ( .A(n63), .ZN(Y[2]) );
  AOI22_X1 U52 ( .A1(S0[2]), .A2(n284), .B1(S1[2]), .B2(n293), .ZN(n63) );
  INV_X1 U53 ( .A(n62), .ZN(Y[3]) );
  AOI22_X1 U54 ( .A1(S0[3]), .A2(n284), .B1(S1[3]), .B2(n292), .ZN(n62) );
  INV_X1 U55 ( .A(n61), .ZN(Y[4]) );
  AOI22_X1 U56 ( .A1(S0[4]), .A2(n284), .B1(S1[4]), .B2(n292), .ZN(n61) );
  INV_X1 U57 ( .A(n60), .ZN(Y[5]) );
  AOI22_X1 U58 ( .A1(S0[5]), .A2(n284), .B1(S1[5]), .B2(n292), .ZN(n60) );
  INV_X1 U59 ( .A(n59), .ZN(Y[6]) );
  AOI22_X1 U60 ( .A1(S0[6]), .A2(n284), .B1(S1[6]), .B2(n292), .ZN(n59) );
  INV_X1 U61 ( .A(n58), .ZN(Y[7]) );
  AOI22_X1 U62 ( .A1(S0[7]), .A2(n284), .B1(S1[7]), .B2(n291), .ZN(n58) );
  INV_X1 U63 ( .A(n57), .ZN(Y[8]) );
  AOI22_X1 U64 ( .A1(S0[8]), .A2(n284), .B1(S1[8]), .B2(n291), .ZN(n57) );
  INV_X1 U65 ( .A(n56), .ZN(Y[9]) );
  AOI22_X1 U66 ( .A1(S0[9]), .A2(n284), .B1(S1[9]), .B2(n291), .ZN(n56) );
  INV_X1 U67 ( .A(n55), .ZN(Y[10]) );
  AOI22_X1 U68 ( .A1(S0[10]), .A2(n284), .B1(S1[10]), .B2(n291), .ZN(n55) );
  INV_X1 U69 ( .A(n54), .ZN(Y[11]) );
  AOI22_X1 U70 ( .A1(S0[11]), .A2(n284), .B1(S1[11]), .B2(n290), .ZN(n54) );
  INV_X1 U71 ( .A(n53), .ZN(Y[12]) );
  AOI22_X1 U72 ( .A1(S0[12]), .A2(n285), .B1(S1[12]), .B2(n290), .ZN(n53) );
  INV_X1 U73 ( .A(n52), .ZN(Y[13]) );
  AOI22_X1 U74 ( .A1(S0[13]), .A2(n285), .B1(S1[13]), .B2(n290), .ZN(n52) );
  INV_X1 U75 ( .A(n51), .ZN(Y[14]) );
  AOI22_X1 U76 ( .A1(S0[14]), .A2(n285), .B1(S1[14]), .B2(n289), .ZN(n51) );
  INV_X1 U77 ( .A(n50), .ZN(Y[15]) );
  AOI22_X1 U78 ( .A1(S0[15]), .A2(n285), .B1(S1[15]), .B2(n289), .ZN(n50) );
endmodule


module SIGN_EXTEND_WIDTH_IN8_WIDTH_OUT32_1 ( A, S, Y );
  input [7:0] A;
  output [31:0] Y;
  input S;
  wire   N0, \Y[31] , \Y[19] ;
  assign Y[7] = A[7];
  assign Y[6] = A[6];
  assign Y[5] = A[5];
  assign Y[4] = A[4];
  assign Y[3] = A[3];
  assign Y[2] = A[2];
  assign Y[1] = A[1];
  assign Y[0] = A[0];
  assign Y[20] = \Y[31] ;
  assign Y[21] = \Y[31] ;
  assign Y[22] = \Y[31] ;
  assign Y[23] = \Y[31] ;
  assign Y[24] = \Y[31] ;
  assign Y[25] = \Y[31] ;
  assign Y[26] = \Y[31] ;
  assign Y[27] = \Y[31] ;
  assign Y[28] = \Y[31] ;
  assign Y[29] = \Y[31] ;
  assign Y[30] = \Y[31] ;
  assign Y[31] = \Y[31] ;
  assign Y[8] = \Y[19] ;
  assign Y[9] = \Y[19] ;
  assign Y[10] = \Y[19] ;
  assign Y[11] = \Y[19] ;
  assign Y[12] = \Y[19] ;
  assign Y[13] = \Y[19] ;
  assign Y[14] = \Y[19] ;
  assign Y[15] = \Y[19] ;
  assign Y[16] = \Y[19] ;
  assign Y[17] = \Y[19] ;
  assign Y[18] = \Y[19] ;
  assign Y[19] = \Y[19] ;

  BUF_X1 U1 ( .A(N0), .Z(\Y[19] ) );
  BUF_X1 U2 ( .A(N0), .Z(\Y[31] ) );
  AND2_X1 U3 ( .A1(S), .A2(A[7]), .ZN(N0) );
endmodule


module SIGN_EXTEND_WIDTH_IN16_WIDTH_OUT32_1 ( A, S, Y );
  input [15:0] A;
  output [31:0] Y;
  input S;
  wire   N0;
  assign Y[15] = A[15];
  assign Y[14] = A[14];
  assign Y[13] = A[13];
  assign Y[12] = A[12];
  assign Y[11] = A[11];
  assign Y[10] = A[10];
  assign Y[9] = A[9];
  assign Y[8] = A[8];
  assign Y[7] = A[7];
  assign Y[6] = A[6];
  assign Y[5] = A[5];
  assign Y[4] = A[4];
  assign Y[3] = A[3];
  assign Y[2] = A[2];
  assign Y[1] = A[1];
  assign Y[0] = A[0];
  assign Y[16] = N0;
  assign Y[17] = N0;
  assign Y[18] = N0;
  assign Y[19] = N0;
  assign Y[20] = N0;
  assign Y[21] = N0;
  assign Y[22] = N0;
  assign Y[23] = N0;
  assign Y[24] = N0;
  assign Y[25] = N0;
  assign Y[26] = N0;
  assign Y[27] = N0;
  assign Y[28] = N0;
  assign Y[29] = N0;
  assign Y[30] = N0;
  assign Y[31] = N0;

  AND2_X1 U1 ( .A1(S), .A2(A[15]), .ZN(N0) );
endmodule


module MUX31_GENERIC_NBIT32_1 ( S2, S1, S0, SEL, Y );
  input [31:0] S2;
  input [31:0] S1;
  input [31:0] S0;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n285, n286;

  BUF_X1 U2 ( .A(n37), .Z(n247) );
  BUF_X1 U3 ( .A(n37), .Z(n248) );
  BUF_X1 U4 ( .A(n36), .Z(n250) );
  BUF_X1 U5 ( .A(n36), .Z(n251) );
  BUF_X1 U6 ( .A(n36), .Z(n252) );
  BUF_X1 U7 ( .A(n38), .Z(n244) );
  BUF_X1 U8 ( .A(n38), .Z(n245) );
  BUF_X1 U9 ( .A(n37), .Z(n249) );
  BUF_X1 U10 ( .A(n38), .Z(n246) );
  INV_X1 U11 ( .A(n53), .ZN(Y[16]) );
  AOI222_X1 U12 ( .A1(S0[16]), .A2(n251), .B1(S1[16]), .B2(n248), .C1(S2[16]), 
        .C2(n245), .ZN(n53) );
  INV_X1 U13 ( .A(n52), .ZN(Y[17]) );
  AOI222_X1 U14 ( .A1(S0[17]), .A2(n251), .B1(S1[17]), .B2(n248), .C1(S2[17]), 
        .C2(n245), .ZN(n52) );
  INV_X1 U15 ( .A(n51), .ZN(Y[18]) );
  AOI222_X1 U16 ( .A1(S0[18]), .A2(n251), .B1(S1[18]), .B2(n248), .C1(S2[18]), 
        .C2(n245), .ZN(n51) );
  INV_X1 U17 ( .A(n50), .ZN(Y[19]) );
  AOI222_X1 U18 ( .A1(S0[19]), .A2(n251), .B1(S1[19]), .B2(n248), .C1(S2[19]), 
        .C2(n245), .ZN(n50) );
  INV_X1 U19 ( .A(n49), .ZN(Y[20]) );
  AOI222_X1 U20 ( .A1(S0[20]), .A2(n251), .B1(S1[20]), .B2(n248), .C1(S2[20]), 
        .C2(n245), .ZN(n49) );
  INV_X1 U21 ( .A(n48), .ZN(Y[21]) );
  AOI222_X1 U22 ( .A1(S0[21]), .A2(n251), .B1(S1[21]), .B2(n248), .C1(S2[21]), 
        .C2(n245), .ZN(n48) );
  INV_X1 U23 ( .A(n47), .ZN(Y[22]) );
  AOI222_X1 U24 ( .A1(S0[22]), .A2(n252), .B1(S1[22]), .B2(n248), .C1(S2[22]), 
        .C2(n245), .ZN(n47) );
  INV_X1 U25 ( .A(n46), .ZN(Y[23]) );
  AOI222_X1 U26 ( .A1(S0[23]), .A2(n252), .B1(S1[23]), .B2(n248), .C1(S2[23]), 
        .C2(n245), .ZN(n46) );
  INV_X1 U27 ( .A(n45), .ZN(Y[24]) );
  AOI222_X1 U28 ( .A1(S0[24]), .A2(n252), .B1(S1[24]), .B2(n249), .C1(S2[24]), 
        .C2(n246), .ZN(n45) );
  INV_X1 U29 ( .A(n44), .ZN(Y[25]) );
  AOI222_X1 U30 ( .A1(S0[25]), .A2(n252), .B1(S1[25]), .B2(n249), .C1(S2[25]), 
        .C2(n246), .ZN(n44) );
  INV_X1 U31 ( .A(n43), .ZN(Y[26]) );
  AOI222_X1 U32 ( .A1(S0[26]), .A2(n252), .B1(S1[26]), .B2(n249), .C1(S2[26]), 
        .C2(n246), .ZN(n43) );
  INV_X1 U33 ( .A(n42), .ZN(Y[27]) );
  AOI222_X1 U34 ( .A1(S0[27]), .A2(n252), .B1(S1[27]), .B2(n249), .C1(S2[27]), 
        .C2(n246), .ZN(n42) );
  INV_X1 U35 ( .A(n41), .ZN(Y[28]) );
  AOI222_X1 U36 ( .A1(S0[28]), .A2(n252), .B1(S1[28]), .B2(n249), .C1(S2[28]), 
        .C2(n246), .ZN(n41) );
  INV_X1 U37 ( .A(n40), .ZN(Y[29]) );
  AOI222_X1 U38 ( .A1(S0[29]), .A2(n252), .B1(S1[29]), .B2(n249), .C1(S2[29]), 
        .C2(n246), .ZN(n40) );
  INV_X1 U39 ( .A(n39), .ZN(Y[30]) );
  AOI222_X1 U40 ( .A1(S0[30]), .A2(n252), .B1(S1[30]), .B2(n249), .C1(S2[30]), 
        .C2(n246), .ZN(n39) );
  INV_X1 U41 ( .A(n35), .ZN(Y[31]) );
  AOI222_X1 U42 ( .A1(S0[31]), .A2(n252), .B1(S1[31]), .B2(n249), .C1(S2[31]), 
        .C2(n246), .ZN(n35) );
  NOR3_X1 U43 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n286), .ZN(n36) );
  NOR3_X1 U44 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n285), .ZN(n37) );
  AND3_X1 U45 ( .A1(n286), .A2(n285), .A3(SEL[2]), .ZN(n38) );
  INV_X1 U46 ( .A(SEL[1]), .ZN(n285) );
  INV_X1 U47 ( .A(SEL[0]), .ZN(n286) );
  INV_X1 U48 ( .A(n69), .ZN(Y[0]) );
  AOI222_X1 U49 ( .A1(S0[0]), .A2(n250), .B1(S1[0]), .B2(n247), .C1(S2[0]), 
        .C2(n244), .ZN(n69) );
  INV_X1 U50 ( .A(n68), .ZN(Y[1]) );
  AOI222_X1 U51 ( .A1(S0[1]), .A2(n250), .B1(S1[1]), .B2(n247), .C1(S2[1]), 
        .C2(n244), .ZN(n68) );
  INV_X1 U52 ( .A(n67), .ZN(Y[2]) );
  AOI222_X1 U53 ( .A1(S0[2]), .A2(n250), .B1(S1[2]), .B2(n247), .C1(S2[2]), 
        .C2(n244), .ZN(n67) );
  INV_X1 U54 ( .A(n66), .ZN(Y[3]) );
  AOI222_X1 U55 ( .A1(S0[3]), .A2(n250), .B1(S1[3]), .B2(n247), .C1(S2[3]), 
        .C2(n244), .ZN(n66) );
  INV_X1 U56 ( .A(n65), .ZN(Y[4]) );
  AOI222_X1 U57 ( .A1(S0[4]), .A2(n250), .B1(S1[4]), .B2(n247), .C1(S2[4]), 
        .C2(n244), .ZN(n65) );
  INV_X1 U58 ( .A(n64), .ZN(Y[5]) );
  AOI222_X1 U59 ( .A1(S0[5]), .A2(n250), .B1(S1[5]), .B2(n247), .C1(S2[5]), 
        .C2(n244), .ZN(n64) );
  INV_X1 U60 ( .A(n63), .ZN(Y[6]) );
  AOI222_X1 U61 ( .A1(S0[6]), .A2(n250), .B1(S1[6]), .B2(n247), .C1(S2[6]), 
        .C2(n244), .ZN(n63) );
  INV_X1 U62 ( .A(n62), .ZN(Y[7]) );
  AOI222_X1 U63 ( .A1(S0[7]), .A2(n250), .B1(S1[7]), .B2(n247), .C1(S2[7]), 
        .C2(n244), .ZN(n62) );
  INV_X1 U64 ( .A(n61), .ZN(Y[8]) );
  AOI222_X1 U65 ( .A1(S0[8]), .A2(n250), .B1(S1[8]), .B2(n247), .C1(S2[8]), 
        .C2(n244), .ZN(n61) );
  INV_X1 U66 ( .A(n60), .ZN(Y[9]) );
  AOI222_X1 U67 ( .A1(S0[9]), .A2(n250), .B1(S1[9]), .B2(n247), .C1(S2[9]), 
        .C2(n244), .ZN(n60) );
  INV_X1 U68 ( .A(n59), .ZN(Y[10]) );
  AOI222_X1 U69 ( .A1(S0[10]), .A2(n250), .B1(S1[10]), .B2(n247), .C1(S2[10]), 
        .C2(n244), .ZN(n59) );
  INV_X1 U70 ( .A(n58), .ZN(Y[11]) );
  AOI222_X1 U71 ( .A1(S0[11]), .A2(n251), .B1(S1[11]), .B2(n247), .C1(S2[11]), 
        .C2(n244), .ZN(n58) );
  INV_X1 U72 ( .A(n57), .ZN(Y[12]) );
  AOI222_X1 U73 ( .A1(S0[12]), .A2(n251), .B1(S1[12]), .B2(n248), .C1(S2[12]), 
        .C2(n245), .ZN(n57) );
  INV_X1 U74 ( .A(n56), .ZN(Y[13]) );
  AOI222_X1 U75 ( .A1(S0[13]), .A2(n251), .B1(S1[13]), .B2(n248), .C1(S2[13]), 
        .C2(n245), .ZN(n56) );
  INV_X1 U76 ( .A(n55), .ZN(Y[14]) );
  AOI222_X1 U77 ( .A1(S0[14]), .A2(n251), .B1(S1[14]), .B2(n248), .C1(S2[14]), 
        .C2(n245), .ZN(n55) );
  INV_X1 U78 ( .A(n54), .ZN(Y[15]) );
  AOI222_X1 U79 ( .A1(S0[15]), .A2(n251), .B1(S1[15]), .B2(n248), .C1(S2[15]), 
        .C2(n245), .ZN(n54) );
endmodule


module REGISTER_GENERIC_WIDTH32_3 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296;

  DFF_X1 \DOUT_reg[31]  ( .D(n68), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[30]  ( .D(n69), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[29]  ( .D(n70), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[28]  ( .D(n71), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[27]  ( .D(n72), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n73), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[25]  ( .D(n74), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[24]  ( .D(n75), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[22]  ( .D(n77), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[21]  ( .D(n78), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[20]  ( .D(n79), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n80), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n81), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n83), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n84), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n89), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n90), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n91), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n92), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n93), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n94), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n95), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n96), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n97), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n98), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n260) );
  BUF_X1 U4 ( .A(n35), .Z(n259) );
  BUF_X1 U5 ( .A(n35), .Z(n258) );
  BUF_X1 U6 ( .A(n34), .Z(n263) );
  NAND2_X1 U7 ( .A1(RST), .A2(n261), .ZN(n35) );
  BUF_X1 U8 ( .A(n34), .Z(n261) );
  BUF_X1 U9 ( .A(n34), .Z(n262) );
  NAND2_X1 U10 ( .A1(n264), .A2(RST), .ZN(n34) );
  INV_X1 U11 ( .A(EN), .ZN(n264) );
  OAI22_X1 U12 ( .A1(n36), .A2(n263), .B1(n260), .B2(n296), .ZN(n99) );
  INV_X1 U13 ( .A(DIN[0]), .ZN(n296) );
  OAI22_X1 U14 ( .A1(n37), .A2(n263), .B1(n260), .B2(n295), .ZN(n98) );
  INV_X1 U15 ( .A(DIN[1]), .ZN(n295) );
  OAI22_X1 U16 ( .A1(n38), .A2(n263), .B1(n260), .B2(n294), .ZN(n97) );
  INV_X1 U17 ( .A(DIN[2]), .ZN(n294) );
  OAI22_X1 U18 ( .A1(n39), .A2(n263), .B1(n260), .B2(n293), .ZN(n96) );
  INV_X1 U19 ( .A(DIN[3]), .ZN(n293) );
  OAI22_X1 U20 ( .A1(n40), .A2(n263), .B1(n260), .B2(n292), .ZN(n95) );
  INV_X1 U21 ( .A(DIN[4]), .ZN(n292) );
  OAI22_X1 U22 ( .A1(n41), .A2(n263), .B1(n260), .B2(n291), .ZN(n94) );
  INV_X1 U23 ( .A(DIN[5]), .ZN(n291) );
  OAI22_X1 U24 ( .A1(n42), .A2(n263), .B1(n260), .B2(n290), .ZN(n93) );
  INV_X1 U25 ( .A(DIN[6]), .ZN(n290) );
  OAI22_X1 U26 ( .A1(n43), .A2(n263), .B1(n260), .B2(n289), .ZN(n92) );
  INV_X1 U27 ( .A(DIN[7]), .ZN(n289) );
  OAI22_X1 U28 ( .A1(n44), .A2(n263), .B1(n260), .B2(n288), .ZN(n91) );
  INV_X1 U29 ( .A(DIN[8]), .ZN(n288) );
  OAI22_X1 U30 ( .A1(n45), .A2(n262), .B1(n260), .B2(n287), .ZN(n90) );
  INV_X1 U31 ( .A(DIN[9]), .ZN(n287) );
  OAI22_X1 U32 ( .A1(n46), .A2(n262), .B1(n259), .B2(n286), .ZN(n89) );
  INV_X1 U33 ( .A(DIN[10]), .ZN(n286) );
  OAI22_X1 U34 ( .A1(n47), .A2(n262), .B1(n259), .B2(n285), .ZN(n88) );
  INV_X1 U35 ( .A(DIN[11]), .ZN(n285) );
  OAI22_X1 U36 ( .A1(n48), .A2(n262), .B1(n259), .B2(n284), .ZN(n87) );
  INV_X1 U37 ( .A(DIN[12]), .ZN(n284) );
  OAI22_X1 U38 ( .A1(n49), .A2(n262), .B1(n259), .B2(n283), .ZN(n86) );
  INV_X1 U39 ( .A(DIN[13]), .ZN(n283) );
  OAI22_X1 U40 ( .A1(n50), .A2(n262), .B1(n259), .B2(n282), .ZN(n85) );
  INV_X1 U41 ( .A(DIN[14]), .ZN(n282) );
  OAI22_X1 U42 ( .A1(n51), .A2(n262), .B1(n259), .B2(n281), .ZN(n84) );
  INV_X1 U43 ( .A(DIN[15]), .ZN(n281) );
  OAI22_X1 U44 ( .A1(n52), .A2(n262), .B1(n259), .B2(n280), .ZN(n83) );
  INV_X1 U45 ( .A(DIN[16]), .ZN(n280) );
  OAI22_X1 U46 ( .A1(n53), .A2(n262), .B1(n259), .B2(n279), .ZN(n82) );
  INV_X1 U47 ( .A(DIN[17]), .ZN(n279) );
  OAI22_X1 U48 ( .A1(n54), .A2(n262), .B1(n259), .B2(n278), .ZN(n81) );
  INV_X1 U49 ( .A(DIN[18]), .ZN(n278) );
  OAI22_X1 U50 ( .A1(n55), .A2(n262), .B1(n259), .B2(n277), .ZN(n80) );
  INV_X1 U51 ( .A(DIN[19]), .ZN(n277) );
  OAI22_X1 U52 ( .A1(n56), .A2(n262), .B1(n259), .B2(n276), .ZN(n79) );
  INV_X1 U53 ( .A(DIN[20]), .ZN(n276) );
  OAI22_X1 U54 ( .A1(n57), .A2(n261), .B1(n258), .B2(n275), .ZN(n78) );
  INV_X1 U55 ( .A(DIN[21]), .ZN(n275) );
  OAI22_X1 U56 ( .A1(n58), .A2(n261), .B1(n258), .B2(n274), .ZN(n77) );
  INV_X1 U57 ( .A(DIN[22]), .ZN(n274) );
  OAI22_X1 U58 ( .A1(n59), .A2(n261), .B1(n258), .B2(n273), .ZN(n76) );
  INV_X1 U59 ( .A(DIN[23]), .ZN(n273) );
  OAI22_X1 U60 ( .A1(n60), .A2(n261), .B1(n258), .B2(n272), .ZN(n75) );
  INV_X1 U61 ( .A(DIN[24]), .ZN(n272) );
  OAI22_X1 U62 ( .A1(n61), .A2(n261), .B1(n258), .B2(n271), .ZN(n74) );
  INV_X1 U63 ( .A(DIN[25]), .ZN(n271) );
  OAI22_X1 U64 ( .A1(n62), .A2(n261), .B1(n258), .B2(n270), .ZN(n73) );
  INV_X1 U65 ( .A(DIN[26]), .ZN(n270) );
  OAI22_X1 U66 ( .A1(n63), .A2(n261), .B1(n258), .B2(n269), .ZN(n72) );
  INV_X1 U67 ( .A(DIN[27]), .ZN(n269) );
  OAI22_X1 U68 ( .A1(n64), .A2(n261), .B1(n258), .B2(n268), .ZN(n71) );
  INV_X1 U69 ( .A(DIN[28]), .ZN(n268) );
  OAI22_X1 U70 ( .A1(n65), .A2(n261), .B1(n258), .B2(n267), .ZN(n70) );
  INV_X1 U71 ( .A(DIN[29]), .ZN(n267) );
  OAI22_X1 U72 ( .A1(n66), .A2(n261), .B1(n258), .B2(n266), .ZN(n69) );
  INV_X1 U73 ( .A(DIN[30]), .ZN(n266) );
  OAI22_X1 U74 ( .A1(n67), .A2(n261), .B1(n258), .B2(n265), .ZN(n68) );
  INV_X1 U75 ( .A(DIN[31]), .ZN(n265) );
endmodule


module REGISTER_GENERIC_WIDTH5_1 ( CLK, RST, EN, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST, EN;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n2, n3, n4, n5, n6,
         n7, n8, n30;

  DFF_X1 \DOUT_reg[3]  ( .D(n15), .CK(CLK), .Q(DOUT[3]), .QN(n12) );
  DFF_X1 \DOUT_reg[1]  ( .D(n17), .CK(CLK), .Q(DOUT[1]), .QN(n10) );
  DFF_X1 \DOUT_reg[0]  ( .D(n18), .CK(CLK), .Q(DOUT[0]), .QN(n9) );
  DFF_X1 \DOUT_reg[2]  ( .D(n16), .CK(CLK), .Q(DOUT[2]), .QN(n11) );
  DFF_X1 \DOUT_reg[4]  ( .D(n14), .CK(CLK), .Q(DOUT[4]), .QN(n13) );
  AND2_X1 U3 ( .A1(RST), .A2(n2), .ZN(n4) );
  OAI21_X1 U4 ( .B1(n13), .B2(n2), .A(n8), .ZN(n14) );
  NAND2_X1 U5 ( .A1(DIN[4]), .A2(n4), .ZN(n8) );
  OAI21_X1 U6 ( .B1(n11), .B2(n2), .A(n6), .ZN(n16) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(n4), .ZN(n6) );
  OAI21_X1 U8 ( .B1(n9), .B2(n2), .A(n3), .ZN(n18) );
  NAND2_X1 U9 ( .A1(DIN[0]), .A2(n4), .ZN(n3) );
  OAI21_X1 U10 ( .B1(n10), .B2(n2), .A(n5), .ZN(n17) );
  NAND2_X1 U11 ( .A1(DIN[1]), .A2(n4), .ZN(n5) );
  OAI21_X1 U12 ( .B1(n12), .B2(n2), .A(n7), .ZN(n15) );
  NAND2_X1 U13 ( .A1(DIN[3]), .A2(n4), .ZN(n7) );
  NAND2_X1 U14 ( .A1(n30), .A2(RST), .ZN(n2) );
  INV_X1 U15 ( .A(EN), .ZN(n30) );
endmodule


module REGISTER_GENERIC_WIDTH32_2 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300;

  DFF_X1 \DOUT_reg[31]  ( .D(n68), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[30]  ( .D(n69), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[29]  ( .D(n70), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[28]  ( .D(n71), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[27]  ( .D(n72), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n73), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[25]  ( .D(n74), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[24]  ( .D(n75), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[22]  ( .D(n77), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[21]  ( .D(n78), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[20]  ( .D(n79), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n80), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n81), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n83), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n84), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n89), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n90), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n91), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n92), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n93), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n94), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n95), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n96), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n97), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n98), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n264) );
  BUF_X1 U4 ( .A(n35), .Z(n263) );
  BUF_X1 U5 ( .A(n35), .Z(n262) );
  NAND2_X1 U6 ( .A1(RST), .A2(n265), .ZN(n35) );
  BUF_X1 U7 ( .A(n34), .Z(n267) );
  BUF_X1 U8 ( .A(n34), .Z(n265) );
  BUF_X1 U9 ( .A(n34), .Z(n266) );
  NAND2_X1 U10 ( .A1(n300), .A2(RST), .ZN(n34) );
  INV_X1 U11 ( .A(EN), .ZN(n300) );
  OAI22_X1 U12 ( .A1(n36), .A2(n267), .B1(n264), .B2(n299), .ZN(n99) );
  INV_X1 U13 ( .A(DIN[0]), .ZN(n299) );
  OAI22_X1 U14 ( .A1(n37), .A2(n267), .B1(n264), .B2(n298), .ZN(n98) );
  INV_X1 U15 ( .A(DIN[1]), .ZN(n298) );
  OAI22_X1 U16 ( .A1(n38), .A2(n267), .B1(n264), .B2(n297), .ZN(n97) );
  INV_X1 U17 ( .A(DIN[2]), .ZN(n297) );
  OAI22_X1 U18 ( .A1(n39), .A2(n267), .B1(n264), .B2(n296), .ZN(n96) );
  INV_X1 U19 ( .A(DIN[3]), .ZN(n296) );
  OAI22_X1 U20 ( .A1(n40), .A2(n267), .B1(n264), .B2(n295), .ZN(n95) );
  INV_X1 U21 ( .A(DIN[4]), .ZN(n295) );
  OAI22_X1 U22 ( .A1(n41), .A2(n267), .B1(n264), .B2(n294), .ZN(n94) );
  INV_X1 U23 ( .A(DIN[5]), .ZN(n294) );
  OAI22_X1 U24 ( .A1(n42), .A2(n267), .B1(n264), .B2(n293), .ZN(n93) );
  INV_X1 U25 ( .A(DIN[6]), .ZN(n293) );
  OAI22_X1 U26 ( .A1(n43), .A2(n267), .B1(n264), .B2(n292), .ZN(n92) );
  INV_X1 U27 ( .A(DIN[7]), .ZN(n292) );
  OAI22_X1 U28 ( .A1(n44), .A2(n267), .B1(n264), .B2(n291), .ZN(n91) );
  INV_X1 U29 ( .A(DIN[8]), .ZN(n291) );
  OAI22_X1 U30 ( .A1(n45), .A2(n266), .B1(n264), .B2(n290), .ZN(n90) );
  INV_X1 U31 ( .A(DIN[9]), .ZN(n290) );
  OAI22_X1 U32 ( .A1(n46), .A2(n266), .B1(n263), .B2(n289), .ZN(n89) );
  INV_X1 U33 ( .A(DIN[10]), .ZN(n289) );
  OAI22_X1 U34 ( .A1(n47), .A2(n266), .B1(n263), .B2(n288), .ZN(n88) );
  INV_X1 U35 ( .A(DIN[11]), .ZN(n288) );
  OAI22_X1 U36 ( .A1(n48), .A2(n266), .B1(n263), .B2(n287), .ZN(n87) );
  INV_X1 U37 ( .A(DIN[12]), .ZN(n287) );
  OAI22_X1 U38 ( .A1(n49), .A2(n266), .B1(n263), .B2(n286), .ZN(n86) );
  INV_X1 U39 ( .A(DIN[13]), .ZN(n286) );
  OAI22_X1 U40 ( .A1(n50), .A2(n266), .B1(n263), .B2(n285), .ZN(n85) );
  INV_X1 U41 ( .A(DIN[14]), .ZN(n285) );
  OAI22_X1 U42 ( .A1(n51), .A2(n266), .B1(n263), .B2(n284), .ZN(n84) );
  INV_X1 U43 ( .A(DIN[15]), .ZN(n284) );
  OAI22_X1 U44 ( .A1(n52), .A2(n266), .B1(n263), .B2(n283), .ZN(n83) );
  INV_X1 U45 ( .A(DIN[16]), .ZN(n283) );
  OAI22_X1 U46 ( .A1(n53), .A2(n266), .B1(n263), .B2(n282), .ZN(n82) );
  INV_X1 U47 ( .A(DIN[17]), .ZN(n282) );
  OAI22_X1 U48 ( .A1(n54), .A2(n266), .B1(n263), .B2(n281), .ZN(n81) );
  INV_X1 U49 ( .A(DIN[18]), .ZN(n281) );
  OAI22_X1 U50 ( .A1(n55), .A2(n266), .B1(n263), .B2(n280), .ZN(n80) );
  INV_X1 U51 ( .A(DIN[19]), .ZN(n280) );
  OAI22_X1 U52 ( .A1(n56), .A2(n266), .B1(n263), .B2(n279), .ZN(n79) );
  INV_X1 U53 ( .A(DIN[20]), .ZN(n279) );
  OAI22_X1 U54 ( .A1(n57), .A2(n265), .B1(n262), .B2(n278), .ZN(n78) );
  INV_X1 U55 ( .A(DIN[21]), .ZN(n278) );
  OAI22_X1 U56 ( .A1(n58), .A2(n265), .B1(n262), .B2(n277), .ZN(n77) );
  INV_X1 U57 ( .A(DIN[22]), .ZN(n277) );
  OAI22_X1 U58 ( .A1(n59), .A2(n265), .B1(n262), .B2(n276), .ZN(n76) );
  INV_X1 U59 ( .A(DIN[23]), .ZN(n276) );
  OAI22_X1 U60 ( .A1(n60), .A2(n265), .B1(n262), .B2(n275), .ZN(n75) );
  INV_X1 U61 ( .A(DIN[24]), .ZN(n275) );
  OAI22_X1 U62 ( .A1(n61), .A2(n265), .B1(n262), .B2(n274), .ZN(n74) );
  INV_X1 U63 ( .A(DIN[25]), .ZN(n274) );
  OAI22_X1 U64 ( .A1(n62), .A2(n265), .B1(n262), .B2(n273), .ZN(n73) );
  INV_X1 U65 ( .A(DIN[26]), .ZN(n273) );
  OAI22_X1 U66 ( .A1(n63), .A2(n265), .B1(n262), .B2(n272), .ZN(n72) );
  INV_X1 U67 ( .A(DIN[27]), .ZN(n272) );
  OAI22_X1 U68 ( .A1(n64), .A2(n265), .B1(n262), .B2(n271), .ZN(n71) );
  INV_X1 U69 ( .A(DIN[28]), .ZN(n271) );
  OAI22_X1 U70 ( .A1(n65), .A2(n265), .B1(n262), .B2(n270), .ZN(n70) );
  INV_X1 U71 ( .A(DIN[29]), .ZN(n270) );
  OAI22_X1 U72 ( .A1(n66), .A2(n265), .B1(n262), .B2(n269), .ZN(n69) );
  INV_X1 U73 ( .A(DIN[30]), .ZN(n269) );
  OAI22_X1 U74 ( .A1(n67), .A2(n265), .B1(n262), .B2(n268), .ZN(n68) );
  INV_X1 U75 ( .A(DIN[31]), .ZN(n268) );
endmodule


module REGISTER_GENERIC_WIDTH32_1 ( CLK, RST, EN, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST, EN;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300;

  DFF_X1 \DOUT_reg[31]  ( .D(n68), .CK(CLK), .Q(DOUT[31]), .QN(n67) );
  DFF_X1 \DOUT_reg[30]  ( .D(n69), .CK(CLK), .Q(DOUT[30]), .QN(n66) );
  DFF_X1 \DOUT_reg[29]  ( .D(n70), .CK(CLK), .Q(DOUT[29]), .QN(n65) );
  DFF_X1 \DOUT_reg[28]  ( .D(n71), .CK(CLK), .Q(DOUT[28]), .QN(n64) );
  DFF_X1 \DOUT_reg[27]  ( .D(n72), .CK(CLK), .Q(DOUT[27]), .QN(n63) );
  DFF_X1 \DOUT_reg[26]  ( .D(n73), .CK(CLK), .Q(DOUT[26]), .QN(n62) );
  DFF_X1 \DOUT_reg[25]  ( .D(n74), .CK(CLK), .Q(DOUT[25]), .QN(n61) );
  DFF_X1 \DOUT_reg[24]  ( .D(n75), .CK(CLK), .Q(DOUT[24]), .QN(n60) );
  DFF_X1 \DOUT_reg[23]  ( .D(n76), .CK(CLK), .Q(DOUT[23]), .QN(n59) );
  DFF_X1 \DOUT_reg[22]  ( .D(n77), .CK(CLK), .Q(DOUT[22]), .QN(n58) );
  DFF_X1 \DOUT_reg[21]  ( .D(n78), .CK(CLK), .Q(DOUT[21]), .QN(n57) );
  DFF_X1 \DOUT_reg[20]  ( .D(n79), .CK(CLK), .Q(DOUT[20]), .QN(n56) );
  DFF_X1 \DOUT_reg[19]  ( .D(n80), .CK(CLK), .Q(DOUT[19]), .QN(n55) );
  DFF_X1 \DOUT_reg[18]  ( .D(n81), .CK(CLK), .Q(DOUT[18]), .QN(n54) );
  DFF_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .Q(DOUT[17]), .QN(n53) );
  DFF_X1 \DOUT_reg[16]  ( .D(n83), .CK(CLK), .Q(DOUT[16]), .QN(n52) );
  DFF_X1 \DOUT_reg[15]  ( .D(n84), .CK(CLK), .Q(DOUT[15]), .QN(n51) );
  DFF_X1 \DOUT_reg[14]  ( .D(n85), .CK(CLK), .Q(DOUT[14]), .QN(n50) );
  DFF_X1 \DOUT_reg[13]  ( .D(n86), .CK(CLK), .Q(DOUT[13]), .QN(n49) );
  DFF_X1 \DOUT_reg[12]  ( .D(n87), .CK(CLK), .Q(DOUT[12]), .QN(n48) );
  DFF_X1 \DOUT_reg[11]  ( .D(n88), .CK(CLK), .Q(DOUT[11]), .QN(n47) );
  DFF_X1 \DOUT_reg[10]  ( .D(n89), .CK(CLK), .Q(DOUT[10]), .QN(n46) );
  DFF_X1 \DOUT_reg[9]  ( .D(n90), .CK(CLK), .Q(DOUT[9]), .QN(n45) );
  DFF_X1 \DOUT_reg[8]  ( .D(n91), .CK(CLK), .Q(DOUT[8]), .QN(n44) );
  DFF_X1 \DOUT_reg[7]  ( .D(n92), .CK(CLK), .Q(DOUT[7]), .QN(n43) );
  DFF_X1 \DOUT_reg[6]  ( .D(n93), .CK(CLK), .Q(DOUT[6]), .QN(n42) );
  DFF_X1 \DOUT_reg[5]  ( .D(n94), .CK(CLK), .Q(DOUT[5]), .QN(n41) );
  DFF_X1 \DOUT_reg[4]  ( .D(n95), .CK(CLK), .Q(DOUT[4]), .QN(n40) );
  DFF_X1 \DOUT_reg[3]  ( .D(n96), .CK(CLK), .Q(DOUT[3]), .QN(n39) );
  DFF_X1 \DOUT_reg[2]  ( .D(n97), .CK(CLK), .Q(DOUT[2]), .QN(n38) );
  DFF_X1 \DOUT_reg[1]  ( .D(n98), .CK(CLK), .Q(DOUT[1]), .QN(n37) );
  DFF_X1 \DOUT_reg[0]  ( .D(n99), .CK(CLK), .Q(DOUT[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n264) );
  BUF_X1 U4 ( .A(n35), .Z(n263) );
  BUF_X1 U5 ( .A(n35), .Z(n262) );
  NAND2_X1 U6 ( .A1(RST), .A2(n265), .ZN(n35) );
  BUF_X1 U7 ( .A(n34), .Z(n267) );
  BUF_X1 U8 ( .A(n34), .Z(n265) );
  BUF_X1 U9 ( .A(n34), .Z(n266) );
  NAND2_X1 U10 ( .A1(n300), .A2(RST), .ZN(n34) );
  INV_X1 U11 ( .A(EN), .ZN(n300) );
  OAI22_X1 U12 ( .A1(n36), .A2(n267), .B1(n264), .B2(n299), .ZN(n99) );
  INV_X1 U13 ( .A(DIN[0]), .ZN(n299) );
  OAI22_X1 U14 ( .A1(n37), .A2(n267), .B1(n264), .B2(n298), .ZN(n98) );
  INV_X1 U15 ( .A(DIN[1]), .ZN(n298) );
  OAI22_X1 U16 ( .A1(n38), .A2(n267), .B1(n264), .B2(n297), .ZN(n97) );
  INV_X1 U17 ( .A(DIN[2]), .ZN(n297) );
  OAI22_X1 U18 ( .A1(n39), .A2(n267), .B1(n264), .B2(n296), .ZN(n96) );
  INV_X1 U19 ( .A(DIN[3]), .ZN(n296) );
  OAI22_X1 U20 ( .A1(n40), .A2(n267), .B1(n264), .B2(n295), .ZN(n95) );
  INV_X1 U21 ( .A(DIN[4]), .ZN(n295) );
  OAI22_X1 U22 ( .A1(n41), .A2(n267), .B1(n264), .B2(n294), .ZN(n94) );
  INV_X1 U23 ( .A(DIN[5]), .ZN(n294) );
  OAI22_X1 U24 ( .A1(n42), .A2(n267), .B1(n264), .B2(n293), .ZN(n93) );
  INV_X1 U25 ( .A(DIN[6]), .ZN(n293) );
  OAI22_X1 U26 ( .A1(n43), .A2(n267), .B1(n264), .B2(n292), .ZN(n92) );
  INV_X1 U27 ( .A(DIN[7]), .ZN(n292) );
  OAI22_X1 U28 ( .A1(n44), .A2(n267), .B1(n264), .B2(n291), .ZN(n91) );
  INV_X1 U29 ( .A(DIN[8]), .ZN(n291) );
  OAI22_X1 U30 ( .A1(n45), .A2(n266), .B1(n264), .B2(n290), .ZN(n90) );
  INV_X1 U31 ( .A(DIN[9]), .ZN(n290) );
  OAI22_X1 U32 ( .A1(n46), .A2(n266), .B1(n263), .B2(n289), .ZN(n89) );
  INV_X1 U33 ( .A(DIN[10]), .ZN(n289) );
  OAI22_X1 U34 ( .A1(n47), .A2(n266), .B1(n263), .B2(n288), .ZN(n88) );
  INV_X1 U35 ( .A(DIN[11]), .ZN(n288) );
  OAI22_X1 U36 ( .A1(n48), .A2(n266), .B1(n263), .B2(n287), .ZN(n87) );
  INV_X1 U37 ( .A(DIN[12]), .ZN(n287) );
  OAI22_X1 U38 ( .A1(n49), .A2(n266), .B1(n263), .B2(n286), .ZN(n86) );
  INV_X1 U39 ( .A(DIN[13]), .ZN(n286) );
  OAI22_X1 U40 ( .A1(n50), .A2(n266), .B1(n263), .B2(n285), .ZN(n85) );
  INV_X1 U41 ( .A(DIN[14]), .ZN(n285) );
  OAI22_X1 U42 ( .A1(n51), .A2(n266), .B1(n263), .B2(n284), .ZN(n84) );
  INV_X1 U43 ( .A(DIN[15]), .ZN(n284) );
  OAI22_X1 U44 ( .A1(n52), .A2(n266), .B1(n263), .B2(n283), .ZN(n83) );
  INV_X1 U45 ( .A(DIN[16]), .ZN(n283) );
  OAI22_X1 U46 ( .A1(n53), .A2(n266), .B1(n263), .B2(n282), .ZN(n82) );
  INV_X1 U47 ( .A(DIN[17]), .ZN(n282) );
  OAI22_X1 U48 ( .A1(n54), .A2(n266), .B1(n263), .B2(n281), .ZN(n81) );
  INV_X1 U49 ( .A(DIN[18]), .ZN(n281) );
  OAI22_X1 U50 ( .A1(n55), .A2(n266), .B1(n263), .B2(n280), .ZN(n80) );
  INV_X1 U51 ( .A(DIN[19]), .ZN(n280) );
  OAI22_X1 U52 ( .A1(n56), .A2(n266), .B1(n263), .B2(n279), .ZN(n79) );
  INV_X1 U53 ( .A(DIN[20]), .ZN(n279) );
  OAI22_X1 U54 ( .A1(n57), .A2(n265), .B1(n262), .B2(n278), .ZN(n78) );
  INV_X1 U55 ( .A(DIN[21]), .ZN(n278) );
  OAI22_X1 U56 ( .A1(n58), .A2(n265), .B1(n262), .B2(n277), .ZN(n77) );
  INV_X1 U57 ( .A(DIN[22]), .ZN(n277) );
  OAI22_X1 U58 ( .A1(n59), .A2(n265), .B1(n262), .B2(n276), .ZN(n76) );
  INV_X1 U59 ( .A(DIN[23]), .ZN(n276) );
  OAI22_X1 U60 ( .A1(n60), .A2(n265), .B1(n262), .B2(n275), .ZN(n75) );
  INV_X1 U61 ( .A(DIN[24]), .ZN(n275) );
  OAI22_X1 U62 ( .A1(n61), .A2(n265), .B1(n262), .B2(n274), .ZN(n74) );
  INV_X1 U63 ( .A(DIN[25]), .ZN(n274) );
  OAI22_X1 U64 ( .A1(n62), .A2(n265), .B1(n262), .B2(n273), .ZN(n73) );
  INV_X1 U65 ( .A(DIN[26]), .ZN(n273) );
  OAI22_X1 U66 ( .A1(n63), .A2(n265), .B1(n262), .B2(n272), .ZN(n72) );
  INV_X1 U67 ( .A(DIN[27]), .ZN(n272) );
  OAI22_X1 U68 ( .A1(n64), .A2(n265), .B1(n262), .B2(n271), .ZN(n71) );
  INV_X1 U69 ( .A(DIN[28]), .ZN(n271) );
  OAI22_X1 U70 ( .A1(n65), .A2(n265), .B1(n262), .B2(n270), .ZN(n70) );
  INV_X1 U71 ( .A(DIN[29]), .ZN(n270) );
  OAI22_X1 U72 ( .A1(n66), .A2(n265), .B1(n262), .B2(n269), .ZN(n69) );
  INV_X1 U73 ( .A(DIN[30]), .ZN(n269) );
  OAI22_X1 U74 ( .A1(n67), .A2(n265), .B1(n262), .B2(n268), .ZN(n68) );
  INV_X1 U75 ( .A(DIN[31]), .ZN(n268) );
endmodule


module MUX21_GENERIC_NBIT32_1 ( S1, S0, SEL, Y );
  input [31:0] S1;
  input [31:0] S0;
  output [31:0] Y;
  input SEL;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295;

  INV_X1 U1 ( .A(n295), .ZN(n285) );
  INV_X1 U2 ( .A(n295), .ZN(n286) );
  BUF_X1 U3 ( .A(n284), .Z(n293) );
  BUF_X1 U4 ( .A(n283), .Z(n292) );
  BUF_X1 U5 ( .A(n283), .Z(n290) );
  BUF_X1 U6 ( .A(n282), .Z(n289) );
  BUF_X1 U7 ( .A(n283), .Z(n291) );
  BUF_X1 U8 ( .A(n282), .Z(n288) );
  BUF_X1 U9 ( .A(n282), .Z(n287) );
  BUF_X1 U10 ( .A(n284), .Z(n295) );
  BUF_X1 U11 ( .A(n284), .Z(n294) );
  INV_X1 U12 ( .A(n65), .ZN(Y[0]) );
  AOI22_X1 U13 ( .A1(S0[0]), .A2(n285), .B1(S1[0]), .B2(n294), .ZN(n65) );
  INV_X1 U14 ( .A(n64), .ZN(Y[1]) );
  AOI22_X1 U15 ( .A1(S0[1]), .A2(n285), .B1(S1[1]), .B2(n294), .ZN(n64) );
  INV_X1 U16 ( .A(n63), .ZN(Y[2]) );
  AOI22_X1 U17 ( .A1(S0[2]), .A2(n285), .B1(S1[2]), .B2(n294), .ZN(n63) );
  INV_X1 U18 ( .A(n62), .ZN(Y[3]) );
  AOI22_X1 U19 ( .A1(S0[3]), .A2(n285), .B1(S1[3]), .B2(n293), .ZN(n62) );
  INV_X1 U20 ( .A(n61), .ZN(Y[4]) );
  AOI22_X1 U21 ( .A1(S0[4]), .A2(n285), .B1(S1[4]), .B2(n293), .ZN(n61) );
  INV_X1 U22 ( .A(n60), .ZN(Y[5]) );
  AOI22_X1 U23 ( .A1(S0[5]), .A2(n285), .B1(S1[5]), .B2(n293), .ZN(n60) );
  INV_X1 U24 ( .A(n59), .ZN(Y[6]) );
  AOI22_X1 U25 ( .A1(S0[6]), .A2(n285), .B1(S1[6]), .B2(n293), .ZN(n59) );
  INV_X1 U26 ( .A(n58), .ZN(Y[7]) );
  AOI22_X1 U27 ( .A1(S0[7]), .A2(n285), .B1(S1[7]), .B2(n292), .ZN(n58) );
  INV_X1 U28 ( .A(n57), .ZN(Y[8]) );
  AOI22_X1 U29 ( .A1(S0[8]), .A2(n285), .B1(S1[8]), .B2(n292), .ZN(n57) );
  INV_X1 U30 ( .A(n56), .ZN(Y[9]) );
  AOI22_X1 U31 ( .A1(S0[9]), .A2(n285), .B1(S1[9]), .B2(n292), .ZN(n56) );
  INV_X1 U32 ( .A(n55), .ZN(Y[10]) );
  AOI22_X1 U33 ( .A1(S0[10]), .A2(n285), .B1(S1[10]), .B2(n292), .ZN(n55) );
  INV_X1 U34 ( .A(n54), .ZN(Y[11]) );
  AOI22_X1 U35 ( .A1(S0[11]), .A2(n285), .B1(S1[11]), .B2(n291), .ZN(n54) );
  INV_X1 U36 ( .A(n53), .ZN(Y[12]) );
  AOI22_X1 U37 ( .A1(S0[12]), .A2(n286), .B1(S1[12]), .B2(n291), .ZN(n53) );
  INV_X1 U38 ( .A(n52), .ZN(Y[13]) );
  AOI22_X1 U39 ( .A1(S0[13]), .A2(n286), .B1(S1[13]), .B2(n291), .ZN(n52) );
  INV_X1 U40 ( .A(n51), .ZN(Y[14]) );
  AOI22_X1 U41 ( .A1(S0[14]), .A2(n286), .B1(S1[14]), .B2(n290), .ZN(n51) );
  INV_X1 U42 ( .A(n50), .ZN(Y[15]) );
  AOI22_X1 U43 ( .A1(S0[15]), .A2(n286), .B1(S1[15]), .B2(n290), .ZN(n50) );
  INV_X1 U44 ( .A(n49), .ZN(Y[16]) );
  AOI22_X1 U45 ( .A1(S0[16]), .A2(n286), .B1(S1[16]), .B2(n290), .ZN(n49) );
  INV_X1 U46 ( .A(n48), .ZN(Y[17]) );
  AOI22_X1 U47 ( .A1(S0[17]), .A2(n286), .B1(S1[17]), .B2(n290), .ZN(n48) );
  INV_X1 U48 ( .A(n47), .ZN(Y[18]) );
  AOI22_X1 U49 ( .A1(S0[18]), .A2(n286), .B1(S1[18]), .B2(n289), .ZN(n47) );
  INV_X1 U50 ( .A(n46), .ZN(Y[19]) );
  AOI22_X1 U51 ( .A1(S0[19]), .A2(n286), .B1(S1[19]), .B2(n289), .ZN(n46) );
  INV_X1 U52 ( .A(n45), .ZN(Y[20]) );
  AOI22_X1 U53 ( .A1(S0[20]), .A2(n286), .B1(S1[20]), .B2(n289), .ZN(n45) );
  INV_X1 U54 ( .A(n44), .ZN(Y[21]) );
  AOI22_X1 U55 ( .A1(S0[21]), .A2(n286), .B1(S1[21]), .B2(n289), .ZN(n44) );
  INV_X1 U56 ( .A(n43), .ZN(Y[22]) );
  AOI22_X1 U57 ( .A1(S0[22]), .A2(n286), .B1(S1[22]), .B2(n288), .ZN(n43) );
  INV_X1 U58 ( .A(n42), .ZN(Y[23]) );
  AOI22_X1 U59 ( .A1(S0[23]), .A2(n286), .B1(S1[23]), .B2(n291), .ZN(n42) );
  INV_X1 U60 ( .A(n34), .ZN(Y[31]) );
  AOI22_X1 U61 ( .A1(S0[31]), .A2(n285), .B1(n294), .B2(S1[31]), .ZN(n34) );
  INV_X1 U62 ( .A(n41), .ZN(Y[24]) );
  AOI22_X1 U63 ( .A1(S0[24]), .A2(n285), .B1(S1[24]), .B2(n288), .ZN(n41) );
  INV_X1 U64 ( .A(n40), .ZN(Y[25]) );
  AOI22_X1 U65 ( .A1(S0[25]), .A2(n286), .B1(S1[25]), .B2(n288), .ZN(n40) );
  INV_X1 U66 ( .A(n39), .ZN(Y[26]) );
  AOI22_X1 U67 ( .A1(S0[26]), .A2(n285), .B1(S1[26]), .B2(n288), .ZN(n39) );
  INV_X1 U68 ( .A(n38), .ZN(Y[27]) );
  AOI22_X1 U69 ( .A1(S0[27]), .A2(n285), .B1(S1[27]), .B2(n287), .ZN(n38) );
  INV_X1 U70 ( .A(n37), .ZN(Y[28]) );
  AOI22_X1 U71 ( .A1(S0[28]), .A2(n285), .B1(S1[28]), .B2(n287), .ZN(n37) );
  INV_X1 U72 ( .A(n36), .ZN(Y[29]) );
  AOI22_X1 U73 ( .A1(S0[29]), .A2(n286), .B1(S1[29]), .B2(n287), .ZN(n36) );
  INV_X1 U74 ( .A(n35), .ZN(Y[30]) );
  AOI22_X1 U75 ( .A1(S0[30]), .A2(n286), .B1(S1[30]), .B2(n287), .ZN(n35) );
  BUF_X1 U76 ( .A(SEL), .Z(n284) );
  BUF_X1 U77 ( .A(SEL), .Z(n283) );
  BUF_X1 U78 ( .A(SEL), .Z(n282) );
endmodule


module FORWARDING_UNIT_WIDTH32_LENGTH5 ( CLK, RST, RS1, RS2, RD3, RD4, RF_WE3, 
        RF_WE4, ForwardA, ForwardB, ForwardC, ForwardD );
  input [4:0] RS1;
  input [4:0] RS2;
  input [4:0] RD3;
  input [4:0] RD4;
  output [2:0] ForwardA;
  output [2:0] ForwardB;
  output [2:0] ForwardC;
  input CLK, RST, RF_WE3, RF_WE4;
  output ForwardD;
  wire   N4, N11, net87466, N18, n80, n92, n81, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n77, n78, n82, n83, n84, n85, n86, n88, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169;
  assign ForwardA[2] = N4;
  assign ForwardB[2] = N11;
  assign ForwardC[1] = net87466;
  assign ForwardC[2] = N18;

  DFFR_X1 \RS1_ID_reg[4]  ( .D(RS1[4]), .CK(CLK), .RN(n161), .QN(n73) );
  DFFR_X1 \RS1_ID_reg[3]  ( .D(RS1[3]), .CK(CLK), .RN(n161), .QN(n72) );
  DFFR_X1 \RS1_ID_reg[2]  ( .D(RS1[2]), .CK(CLK), .RN(n161), .QN(n78) );
  DFFR_X1 \RS1_ID_reg[1]  ( .D(RS1[1]), .CK(CLK), .RN(n161), .QN(n82) );
  DFFR_X1 \RS1_ID_reg[0]  ( .D(RS1[0]), .CK(CLK), .RN(n161), .QN(n158) );
  DFFR_X1 \RS2_ID_reg[4]  ( .D(RS2[4]), .CK(CLK), .RN(n161), .QN(n156) );
  DFF_X1 \RS2_EX_reg[4]  ( .D(n85), .CK(CLK), .QN(n83) );
  DFFR_X1 \RS2_ID_reg[3]  ( .D(RS2[3]), .CK(CLK), .RN(n161), .QN(n77) );
  DFF_X1 \RS2_EX_reg[3]  ( .D(n86), .CK(CLK), .QN(n157) );
  DFFR_X1 \RS2_ID_reg[2]  ( .D(RS2[2]), .CK(CLK), .RN(n161), .Q(n80) );
  DFF_X1 \RS2_EX_reg[2]  ( .D(n165), .CK(CLK), .Q(n81), .QN(n160) );
  DFFR_X1 \RS2_ID_reg[1]  ( .D(RS2[1]), .CK(CLK), .RN(n161), .QN(n75) );
  DFF_X1 \RS2_EX_reg[1]  ( .D(n88), .CK(CLK), .QN(n84) );
  DFFR_X1 \RS2_ID_reg[0]  ( .D(RS2[0]), .CK(CLK), .RN(n161), .Q(n74) );
  DFF_X1 \RS2_EX_reg[0]  ( .D(n166), .CK(CLK), .Q(n92), .QN(n159) );
  NAND3_X1 U70 ( .A1(n22), .A2(RF_WE4), .A3(n23), .ZN(n16) );
  XOR2_X1 U71 ( .A(RS1[4]), .B(RD4[4]), .Z(n31) );
  XOR2_X1 U72 ( .A(RS1[3]), .B(RD4[3]), .Z(n30) );
  XOR2_X1 U73 ( .A(RS1[2]), .B(RD4[2]), .Z(n29) );
  XOR2_X1 U74 ( .A(RS1[1]), .B(RD4[1]), .Z(n28) );
  XOR2_X1 U75 ( .A(RS1[0]), .B(RD4[0]), .Z(n32) );
  XOR2_X1 U76 ( .A(RS1[4]), .B(RD3[4]), .Z(n39) );
  XOR2_X1 U77 ( .A(RS1[1]), .B(RD3[1]), .Z(n38) );
  XOR2_X1 U78 ( .A(n80), .B(RD4[2]), .Z(n45) );
  XOR2_X1 U79 ( .A(n74), .B(RD4[0]), .Z(n44) );
  XOR2_X1 U80 ( .A(n80), .B(RD3[2]), .Z(n55) );
  XOR2_X1 U81 ( .A(n74), .B(RD3[0]), .Z(n54) );
  XOR2_X1 U82 ( .A(n77), .B(RD3[3]), .Z(n51) );
  XOR2_X1 U83 ( .A(n75), .B(RD3[1]), .Z(n50) );
  XOR2_X1 U84 ( .A(n72), .B(RD3[3]), .Z(n68) );
  XOR2_X1 U85 ( .A(n82), .B(RD3[1]), .Z(n67) );
  XOR2_X1 U86 ( .A(n78), .B(RD3[2]), .Z(n66) );
  OAI21_X1 U3 ( .B1(n21), .B2(RD4[3]), .A(n157), .ZN(n20) );
  NOR2_X1 U4 ( .A1(net87466), .A2(N18), .ZN(ForwardC[0]) );
  INV_X1 U5 ( .A(n162), .ZN(n161) );
  NOR2_X1 U6 ( .A1(n24), .A2(n25), .ZN(N18) );
  AND4_X1 U7 ( .A1(n24), .A2(n169), .A3(n26), .A4(n27), .ZN(net87466) );
  NOR2_X1 U8 ( .A1(n168), .A2(n32), .ZN(n26) );
  NOR4_X1 U9 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n27) );
  INV_X1 U10 ( .A(n25), .ZN(n169) );
  NOR2_X1 U11 ( .A1(n41), .A2(n164), .ZN(N11) );
  INV_X1 U12 ( .A(n40), .ZN(n164) );
  NOR2_X1 U13 ( .A1(n56), .A2(n163), .ZN(N4) );
  INV_X1 U14 ( .A(n57), .ZN(n163) );
  INV_X1 U15 ( .A(RST), .ZN(n162) );
  NOR2_X1 U16 ( .A1(N11), .A2(ForwardB[1]), .ZN(ForwardB[0]) );
  NOR2_X1 U17 ( .A1(N4), .A2(ForwardA[1]), .ZN(ForwardA[0]) );
  NOR4_X1 U18 ( .A1(RS1[3]), .A2(RS1[4]), .A3(RS1[2]), .A4(n33), .ZN(n25) );
  OR2_X1 U19 ( .A1(RS1[1]), .A2(RS1[0]), .ZN(n33) );
  NOR3_X1 U20 ( .A1(n38), .A2(n167), .A3(n39), .ZN(n37) );
  NAND4_X1 U21 ( .A1(n34), .A2(n35), .A3(n36), .A4(n37), .ZN(n24) );
  XNOR2_X1 U22 ( .A(RD3[2]), .B(RS1[2]), .ZN(n35) );
  XNOR2_X1 U23 ( .A(RD3[0]), .B(RS1[0]), .ZN(n34) );
  XNOR2_X1 U24 ( .A(RD3[3]), .B(RS1[3]), .ZN(n36) );
  INV_X1 U25 ( .A(RF_WE4), .ZN(n168) );
  INV_X1 U26 ( .A(RF_WE3), .ZN(n167) );
  OAI22_X1 U27 ( .A1(n77), .A2(n162), .B1(n161), .B2(n157), .ZN(n86) );
  OAI22_X1 U28 ( .A1(n75), .A2(n162), .B1(n84), .B2(n161), .ZN(n88) );
  OAI22_X1 U29 ( .A1(n162), .A2(n156), .B1(n83), .B2(n161), .ZN(n85) );
  INV_X1 U30 ( .A(n14), .ZN(n166) );
  AOI22_X1 U31 ( .A1(n161), .A2(n74), .B1(n162), .B2(n92), .ZN(n14) );
  INV_X1 U32 ( .A(n15), .ZN(n165) );
  AOI22_X1 U33 ( .A1(n161), .A2(n80), .B1(n162), .B2(n81), .ZN(n15) );
  NOR4_X1 U34 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(ForwardD) );
  XNOR2_X1 U35 ( .A(n83), .B(RD4[4]), .ZN(n19) );
  OAI21_X1 U36 ( .B1(RD4[3]), .B2(n157), .A(n20), .ZN(n17) );
  XNOR2_X1 U37 ( .A(n84), .B(RD4[1]), .ZN(n18) );
  XNOR2_X1 U38 ( .A(n82), .B(RD4[1]), .ZN(n60) );
  XNOR2_X1 U39 ( .A(n72), .B(RD4[3]), .ZN(n63) );
  AND4_X1 U40 ( .A1(n159), .A2(n160), .A3(n84), .A4(n83), .ZN(n21) );
  XNOR2_X1 U41 ( .A(n78), .B(RD4[2]), .ZN(n61) );
  NAND4_X1 U42 ( .A1(n75), .A2(n77), .A3(n49), .A4(n156), .ZN(n40) );
  NOR2_X1 U43 ( .A1(n74), .A2(n80), .ZN(n49) );
  XNOR2_X1 U44 ( .A(RD4[3]), .B(n77), .ZN(n48) );
  NAND4_X1 U45 ( .A1(n50), .A2(n51), .A3(RF_WE3), .A4(n52), .ZN(n41) );
  NOR3_X1 U46 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n52) );
  NAND4_X1 U47 ( .A1(n82), .A2(n158), .A3(n78), .A4(n65), .ZN(n57) );
  AND2_X1 U48 ( .A1(n73), .A2(n72), .ZN(n65) );
  NAND4_X1 U49 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(n56) );
  NOR3_X1 U50 ( .A1(n70), .A2(n71), .A3(n167), .ZN(n69) );
  XNOR2_X1 U51 ( .A(n81), .B(RD4[2]), .ZN(n22) );
  XNOR2_X1 U52 ( .A(n156), .B(RD4[4]), .ZN(n46) );
  XNOR2_X1 U53 ( .A(n158), .B(RD4[0]), .ZN(n62) );
  XNOR2_X1 U54 ( .A(RD3[4]), .B(n73), .ZN(n71) );
  XNOR2_X1 U55 ( .A(n92), .B(RD4[0]), .ZN(n23) );
  XNOR2_X1 U56 ( .A(n156), .B(RD3[4]), .ZN(n53) );
  XNOR2_X1 U57 ( .A(n158), .B(RD3[0]), .ZN(n70) );
  AND4_X1 U58 ( .A1(n56), .A2(n57), .A3(n58), .A4(n59), .ZN(ForwardA[1]) );
  NOR2_X1 U59 ( .A1(n63), .A2(n64), .ZN(n58) );
  NOR4_X1 U60 ( .A1(n60), .A2(n61), .A3(n168), .A4(n62), .ZN(n59) );
  XNOR2_X1 U61 ( .A(n73), .B(RD4[4]), .ZN(n64) );
  AND4_X1 U62 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(ForwardB[1]) );
  NOR2_X1 U63 ( .A1(n47), .A2(n48), .ZN(n42) );
  NOR4_X1 U64 ( .A1(n168), .A2(n44), .A3(n45), .A4(n46), .ZN(n43) );
  XNOR2_X1 U65 ( .A(RD4[1]), .B(n75), .ZN(n47) );
endmodule


module DLX_DP_WIDTH32_LENGTH5_RADIX4_OPCODE6_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n12, n13, n19,
         n21, n23, n25, n29, n30, n31, n34, n36, n37, n38, n43, n44, n45, n46,
         n49, n52, n53, n55, n57, n58, n59, n61, n62, n65, n68, n72, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2_X1 U22 ( .A(n19), .B(n187), .Z(SUM[31]) );
  XOR2_X1 U23 ( .A(n31), .B(n192), .Z(SUM[27]) );
  XOR2_X1 U24 ( .A(A[25]), .B(n194), .Z(SUM[25]) );
  XOR2_X1 U27 ( .A(A[29]), .B(n191), .Z(SUM[29]) );
  XOR2_X1 U28 ( .A(n4), .B(A[26]), .Z(SUM[26]) );
  XOR2_X1 U42 ( .A(n193), .B(n190), .Z(SUM[28]) );
  NAND3_X1 U94 ( .A1(A[26]), .A2(A[27]), .A3(A[25]), .ZN(n30) );
  NAND3_X1 U97 ( .A1(A[22]), .A2(A[23]), .A3(A[21]), .ZN(n37) );
  NOR2_X1 U2 ( .A1(n220), .A2(SUM[2]), .ZN(n52) );
  NOR2_X1 U3 ( .A1(n219), .A2(n57), .ZN(n12) );
  INV_X1 U4 ( .A(n52), .ZN(n219) );
  XNOR2_X1 U5 ( .A(n205), .B(n62), .ZN(SUM[14]) );
  NOR2_X1 U6 ( .A1(n215), .A2(n58), .ZN(n68) );
  INV_X1 U7 ( .A(n12), .ZN(n215) );
  NOR2_X1 U8 ( .A1(n207), .A2(n210), .ZN(n65) );
  INV_X1 U9 ( .A(n68), .ZN(n210) );
  AND4_X1 U10 ( .A1(n52), .A2(n53), .A3(n209), .A4(n55), .ZN(n1) );
  NOR2_X1 U11 ( .A1(n206), .A2(n59), .ZN(n53) );
  INV_X1 U12 ( .A(n58), .ZN(n209) );
  NOR2_X1 U13 ( .A1(n207), .A2(n57), .ZN(n55) );
  INV_X1 U14 ( .A(n36), .ZN(n198) );
  INV_X1 U15 ( .A(n29), .ZN(n194) );
  XNOR2_X1 U16 ( .A(n206), .B(n65), .ZN(SUM[13]) );
  XNOR2_X1 U17 ( .A(n204), .B(n61), .ZN(SUM[15]) );
  INV_X1 U18 ( .A(n21), .ZN(n188) );
  INV_X1 U19 ( .A(n23), .ZN(n191) );
  INV_X1 U20 ( .A(n25), .ZN(n193) );
  INV_X1 U21 ( .A(n34), .ZN(n195) );
  XNOR2_X1 U25 ( .A(n218), .B(n52), .ZN(SUM[4]) );
  XNOR2_X1 U26 ( .A(n217), .B(n6), .ZN(SUM[5]) );
  XNOR2_X1 U29 ( .A(n216), .B(n13), .ZN(SUM[6]) );
  XNOR2_X1 U30 ( .A(n214), .B(n7), .ZN(SUM[7]) );
  XNOR2_X1 U31 ( .A(n213), .B(n12), .ZN(SUM[8]) );
  XNOR2_X1 U32 ( .A(n208), .B(n72), .ZN(SUM[11]) );
  XNOR2_X1 U33 ( .A(n207), .B(n68), .ZN(SUM[12]) );
  XNOR2_X1 U34 ( .A(n1), .B(n203), .ZN(SUM[16]) );
  XNOR2_X1 U35 ( .A(n201), .B(n46), .ZN(SUM[18]) );
  XNOR2_X1 U36 ( .A(n199), .B(n8), .ZN(SUM[19]) );
  XNOR2_X1 U37 ( .A(n197), .B(n198), .ZN(SUM[21]) );
  XNOR2_X1 U38 ( .A(n5), .B(n196), .ZN(SUM[22]) );
  INV_X1 U39 ( .A(n2), .ZN(n200) );
  NAND4_X1 U40 ( .A1(A[11]), .A2(A[10]), .A3(A[9]), .A4(A[8]), .ZN(n58) );
  NAND4_X1 U41 ( .A1(A[4]), .A2(A[5]), .A3(A[6]), .A4(A[7]), .ZN(n57) );
  NOR2_X1 U43 ( .A1(n189), .A2(n23), .ZN(n21) );
  INV_X1 U44 ( .A(A[29]), .ZN(n189) );
  NOR2_X1 U45 ( .A1(n36), .A2(n37), .ZN(n34) );
  NOR2_X1 U46 ( .A1(n29), .A2(n30), .ZN(n25) );
  INV_X1 U47 ( .A(A[12]), .ZN(n207) );
  NAND2_X1 U48 ( .A1(n25), .A2(A[28]), .ZN(n23) );
  NAND2_X1 U49 ( .A1(n2), .A2(A[20]), .ZN(n36) );
  NAND2_X1 U50 ( .A1(n34), .A2(A[24]), .ZN(n29) );
  AND2_X1 U51 ( .A1(A[21]), .A2(n198), .ZN(n5) );
  AND2_X1 U52 ( .A1(n65), .A2(A[13]), .ZN(n62) );
  AND2_X1 U53 ( .A1(n1), .A2(n43), .ZN(n2) );
  NOR2_X1 U54 ( .A1(n44), .A2(n45), .ZN(n43) );
  NAND2_X1 U55 ( .A1(A[19]), .A2(A[18]), .ZN(n45) );
  NAND2_X1 U56 ( .A1(A[16]), .A2(A[17]), .ZN(n44) );
  INV_X1 U57 ( .A(A[13]), .ZN(n206) );
  INV_X1 U58 ( .A(A[3]), .ZN(n220) );
  AND2_X1 U59 ( .A1(A[25]), .A2(n194), .ZN(n4) );
  INV_X1 U60 ( .A(A[2]), .ZN(SUM[2]) );
  NAND2_X1 U61 ( .A1(A[22]), .A2(n5), .ZN(n38) );
  AND2_X1 U62 ( .A1(n62), .A2(A[14]), .ZN(n61) );
  NAND2_X1 U63 ( .A1(A[14]), .A2(A[15]), .ZN(n59) );
  NAND2_X1 U64 ( .A1(n21), .A2(A[30]), .ZN(n19) );
  XNOR2_X1 U65 ( .A(n188), .B(A[30]), .ZN(SUM[30]) );
  NAND2_X1 U66 ( .A1(A[26]), .A2(n4), .ZN(n31) );
  XNOR2_X1 U67 ( .A(n38), .B(A[23]), .ZN(SUM[23]) );
  NOR2_X1 U68 ( .A1(n49), .A2(n202), .ZN(n46) );
  INV_X1 U69 ( .A(A[17]), .ZN(n202) );
  NOR2_X1 U70 ( .A1(n3), .A2(n211), .ZN(n72) );
  INV_X1 U71 ( .A(A[10]), .ZN(n211) );
  NAND2_X1 U72 ( .A1(n12), .A2(A[8]), .ZN(n9) );
  NAND2_X1 U73 ( .A1(n1), .A2(A[16]), .ZN(n49) );
  AND2_X1 U74 ( .A1(n52), .A2(A[4]), .ZN(n6) );
  AND2_X1 U75 ( .A1(n6), .A2(A[5]), .ZN(n13) );
  OR2_X1 U76 ( .A1(n212), .A2(n9), .ZN(n3) );
  INV_X1 U77 ( .A(A[9]), .ZN(n212) );
  AND2_X1 U78 ( .A1(A[6]), .A2(n13), .ZN(n7) );
  AND2_X1 U79 ( .A1(A[18]), .A2(n46), .ZN(n8) );
  INV_X1 U80 ( .A(A[16]), .ZN(n203) );
  INV_X1 U81 ( .A(A[22]), .ZN(n196) );
  INV_X1 U82 ( .A(A[8]), .ZN(n213) );
  XNOR2_X1 U83 ( .A(n195), .B(A[24]), .ZN(SUM[24]) );
  INV_X1 U84 ( .A(A[6]), .ZN(n216) );
  INV_X1 U85 ( .A(A[18]), .ZN(n201) );
  INV_X1 U86 ( .A(A[5]), .ZN(n217) );
  INV_X1 U87 ( .A(A[14]), .ZN(n205) );
  INV_X1 U88 ( .A(A[4]), .ZN(n218) );
  INV_X1 U89 ( .A(A[7]), .ZN(n214) );
  INV_X1 U90 ( .A(A[21]), .ZN(n197) );
  INV_X1 U91 ( .A(A[15]), .ZN(n204) );
  INV_X1 U92 ( .A(A[19]), .ZN(n199) );
  INV_X1 U93 ( .A(A[11]), .ZN(n208) );
  XNOR2_X1 U95 ( .A(n220), .B(A[2]), .ZN(SUM[3]) );
  XNOR2_X1 U96 ( .A(n9), .B(A[9]), .ZN(SUM[9]) );
  XNOR2_X1 U98 ( .A(n3), .B(A[10]), .ZN(SUM[10]) );
  XNOR2_X1 U99 ( .A(n49), .B(A[17]), .ZN(SUM[17]) );
  XNOR2_X1 U100 ( .A(n200), .B(A[20]), .ZN(SUM[20]) );
  INV_X1 U101 ( .A(A[28]), .ZN(n190) );
  INV_X1 U102 ( .A(A[27]), .ZN(n192) );
  INV_X1 U103 ( .A(A[31]), .ZN(n187) );
endmodule


module DLX_DP_WIDTH32_LENGTH5_RADIX4_OPCODE6_DW01_add_5 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n63, n64, n65, n66, n140, n141, n142, n143,
         n144, n145, n147, n148, n149, n150, n151, n152, n153, n154;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2_X1 U60 ( .A(A[9]), .B(n78), .Z(SUM[9]) );
  XOR2_X1 U61 ( .A(A[6]), .B(n64), .Z(SUM[6]) );
  XOR2_X1 U62 ( .A(n84), .B(A[31]), .Z(SUM[31]) );
  NAND3_X1 U63 ( .A1(A[28]), .A2(n86), .A3(A[29]), .ZN(n85) );
  XOR2_X1 U64 ( .A(A[28]), .B(n65), .Z(SUM[28]) );
  NAND3_X1 U65 ( .A1(A[24]), .A2(n90), .A3(A[25]), .ZN(n88) );
  XOR2_X1 U66 ( .A(A[24]), .B(n90), .Z(SUM[24]) );
  NAND3_X1 U67 ( .A1(A[20]), .A2(n94), .A3(A[21]), .ZN(n92) );
  XOR2_X1 U68 ( .A(A[20]), .B(n94), .Z(SUM[20]) );
  NAND3_X1 U69 ( .A1(A[16]), .A2(n98), .A3(A[17]), .ZN(n96) );
  XOR2_X1 U70 ( .A(A[16]), .B(n98), .Z(SUM[16]) );
  NAND3_X1 U71 ( .A1(A[12]), .A2(n102), .A3(A[13]), .ZN(n100) );
  XOR2_X1 U72 ( .A(A[12]), .B(n102), .Z(SUM[12]) );
  NAND3_X1 U73 ( .A1(A[6]), .A2(n81), .A3(A[7]), .ZN(n79) );
  NAND3_X1 U38 ( .A1(A[28]), .A2(n65), .A3(A[29]), .ZN(n66) );
  NOR3_X1 U2 ( .A1(n150), .A2(n88), .A3(n143), .ZN(n65) );
  NOR3_X1 U3 ( .A1(n152), .A2(n92), .A3(n144), .ZN(n90) );
  NOR3_X1 U4 ( .A1(n142), .A2(n96), .A3(n148), .ZN(n94) );
  NOR3_X1 U5 ( .A1(n151), .A2(n104), .A3(n141), .ZN(n102) );
  NOR2_X1 U6 ( .A1(n100), .A2(n63), .ZN(n98) );
  OR2_X1 U7 ( .A1(n145), .A2(n153), .ZN(n63) );
  NOR3_X1 U8 ( .A1(n154), .A2(n83), .A3(n149), .ZN(n64) );
  NOR3_X1 U9 ( .A1(n154), .A2(n83), .A3(n149), .ZN(n81) );
  XNOR2_X1 U10 ( .A(n148), .B(n97), .ZN(SUM[19]) );
  NOR2_X1 U11 ( .A1(n96), .A2(n142), .ZN(n97) );
  XNOR2_X1 U12 ( .A(n144), .B(n93), .ZN(SUM[23]) );
  NOR2_X1 U13 ( .A1(n92), .A2(n152), .ZN(n93) );
  XNOR2_X1 U14 ( .A(n143), .B(n89), .ZN(SUM[27]) );
  NOR2_X1 U15 ( .A1(n88), .A2(n150), .ZN(n89) );
  NOR2_X1 U16 ( .A1(n85), .A2(n147), .ZN(n84) );
  NAND2_X1 U17 ( .A1(A[3]), .A2(A[2]), .ZN(n83) );
  NOR2_X1 U18 ( .A1(n79), .A2(n140), .ZN(n78) );
  INV_X1 U19 ( .A(A[8]), .ZN(n140) );
  XNOR2_X1 U20 ( .A(A[30]), .B(n66), .ZN(SUM[30]) );
  XNOR2_X1 U21 ( .A(A[22]), .B(n92), .ZN(SUM[22]) );
  NAND2_X1 U22 ( .A1(n78), .A2(A[9]), .ZN(n104) );
  XNOR2_X1 U23 ( .A(A[21]), .B(n95), .ZN(SUM[21]) );
  NAND2_X1 U24 ( .A1(A[20]), .A2(n94), .ZN(n95) );
  XNOR2_X1 U25 ( .A(A[25]), .B(n91), .ZN(SUM[25]) );
  NAND2_X1 U26 ( .A1(A[24]), .A2(n90), .ZN(n91) );
  NOR3_X1 U27 ( .A1(n150), .A2(n88), .A3(n143), .ZN(n86) );
  INV_X1 U28 ( .A(A[5]), .ZN(n149) );
  INV_X1 U29 ( .A(A[4]), .ZN(n154) );
  XNOR2_X1 U30 ( .A(A[29]), .B(n87), .ZN(SUM[29]) );
  NAND2_X1 U31 ( .A1(A[28]), .A2(n65), .ZN(n87) );
  INV_X1 U32 ( .A(A[11]), .ZN(n141) );
  INV_X1 U33 ( .A(A[10]), .ZN(n151) );
  INV_X1 U34 ( .A(A[15]), .ZN(n145) );
  INV_X1 U35 ( .A(A[14]), .ZN(n153) );
  XNOR2_X1 U36 ( .A(A[26]), .B(n88), .ZN(SUM[26]) );
  XNOR2_X1 U37 ( .A(A[18]), .B(n96), .ZN(SUM[18]) );
  XNOR2_X1 U39 ( .A(A[3]), .B(SUM[2]), .ZN(SUM[3]) );
  XNOR2_X1 U40 ( .A(A[4]), .B(n83), .ZN(SUM[4]) );
  XNOR2_X1 U41 ( .A(n149), .B(n82), .ZN(SUM[5]) );
  NOR2_X1 U42 ( .A1(n83), .A2(n154), .ZN(n82) );
  XNOR2_X1 U43 ( .A(A[7]), .B(n80), .ZN(SUM[7]) );
  NAND2_X1 U44 ( .A1(A[6]), .A2(n64), .ZN(n80) );
  XNOR2_X1 U45 ( .A(A[8]), .B(n79), .ZN(SUM[8]) );
  XNOR2_X1 U46 ( .A(n141), .B(n105), .ZN(SUM[11]) );
  NOR2_X1 U47 ( .A1(n104), .A2(n151), .ZN(n105) );
  XNOR2_X1 U48 ( .A(n145), .B(n101), .ZN(SUM[15]) );
  NOR2_X1 U49 ( .A1(n100), .A2(n153), .ZN(n101) );
  XNOR2_X1 U50 ( .A(A[17]), .B(n99), .ZN(SUM[17]) );
  NAND2_X1 U51 ( .A1(A[16]), .A2(n98), .ZN(n99) );
  INV_X1 U52 ( .A(A[27]), .ZN(n143) );
  INV_X1 U53 ( .A(A[26]), .ZN(n150) );
  INV_X1 U54 ( .A(A[2]), .ZN(SUM[2]) );
  INV_X1 U55 ( .A(A[19]), .ZN(n148) );
  INV_X1 U56 ( .A(A[23]), .ZN(n144) );
  INV_X1 U57 ( .A(A[18]), .ZN(n142) );
  INV_X1 U58 ( .A(A[22]), .ZN(n152) );
  XNOR2_X1 U59 ( .A(A[14]), .B(n100), .ZN(SUM[14]) );
  INV_X1 U74 ( .A(A[30]), .ZN(n147) );
  XNOR2_X1 U75 ( .A(A[10]), .B(n104), .ZN(SUM[10]) );
  XNOR2_X1 U76 ( .A(A[13]), .B(n103), .ZN(SUM[13]) );
  NAND2_X1 U77 ( .A1(A[12]), .A2(n102), .ZN(n103) );
endmodule


module DLX_DP_WIDTH32_LENGTH5_RADIX4_OPCODE6 ( CLK, RST, EN1, PC_IN, EN2, 
        RF_RD1, RF_RD2, MuxIMM_SEL, SIGN_EN, RD, RS1, RS2, IMM16, IMM26, EN3, 
        MuxA_SEL, MuxB_SEL, EQ_COND, JUMP_EN, RF_WE3, .ALU_OPCODE({
        \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , 
        \ALU_OPCODE[0] }), EN4, RF_WE4, SIGN_LD_EN, MuxLD_SEL, MuxSW_SEL, 
        NPC_OUT, DRAM_ADDR, DRAM_IN, DRAM_OUT, MuxWB_SEL, RF_WE, JUMP_LINK );
  input [31:0] PC_IN;
  input [4:0] RD;
  input [4:0] RS1;
  input [4:0] RS2;
  input [15:0] IMM16;
  input [25:0] IMM26;
  input [2:0] MuxLD_SEL;
  input [2:0] MuxSW_SEL;
  output [31:0] NPC_OUT;
  output [5:0] DRAM_ADDR;
  input [31:0] DRAM_IN;
  output [31:0] DRAM_OUT;
  input CLK, RST, EN1, EN2, RF_RD1, RF_RD2, MuxIMM_SEL, SIGN_EN, EN3, MuxA_SEL,
         MuxB_SEL, EQ_COND, JUMP_EN, RF_WE3, \ALU_OPCODE[4] , \ALU_OPCODE[3] ,
         \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] , EN4, RF_WE4,
         SIGN_LD_EN, MuxWB_SEL, RF_WE, JUMP_LINK;
  wire   Z, MuxMEM_SEL, FwdD_SEL, n27, n28, n29;
  wire   [4:0] ALU_OPCODE;
  wire   [31:0] NPC;
  wire   [31:0] NPC1;
  wire   [31:0] RetADDR;
  wire   [31:0] MuxWB_OUT;
  wire   [31:0] WR_DATA;
  wire   [31:0] RegA_IN;
  wire   [31:0] RegB_IN;
  wire   [4:0] RD4;
  wire   [31:0] RegA_OUT;
  wire   [31:0] RegB_OUT;
  wire   [31:0] IMMS16;
  wire   [31:0] IMMS26;
  wire   [31:0] IMM;
  wire   [31:0] RegIMM_OUT;
  wire   [4:0] RD2;
  wire   [31:0] NPC2;
  wire   [31:0] MuxA_OUT;
  wire   [31:0] MuxB_OUT;
  wire   [31:6] RegALU3_OUT;
  wire   [2:0] FwdA_SEL;
  wire   [31:0] A;
  wire   [2:0] FwdB_SEL;
  wire   [31:0] B;
  wire   [31:0] Y;
  wire   [2:0] FwdC_SEL;
  wire   [31:0] Z_IN;
  wire   [31:0] RegME_OUT;
  wire   [4:0] RD3;
  wire   [31:0] NPC3;
  wire   [31:0] RegLMD_OUT;
  wire   [31:0] LMD_8;
  wire   [31:0] LMD_16;
  wire   [31:0] MuxLD_OUT;
  wire   [31:0] MuxFWD_OUT;
  wire   [31:0] MEM_8;
  wire   [31:0] MEM_16;
  wire   [31:0] NPC4;
  wire   [31:0] RegALU4_OUT;

  REGISTER_GENERIC_WIDTH32_11 RegNPC1 ( .CLK(CLK), .RST(n28), .EN(EN1), .DIN(
        NPC), .DOUT(NPC1) );
  MUX21_GENERIC_NBIT32_0 MuxWR ( .S1(RetADDR), .S0(MuxWB_OUT), .SEL(JUMP_LINK), 
        .Y(WR_DATA) );
  REGISTER_FILE_WIDTH32_LENGTH5 RegFILE ( .CLK(CLK), .RST(n27), .EN(EN2), 
        .RD1(RF_RD1), .RD2(RF_RD2), .WR(RF_WE), .DATAIN(WR_DATA), .OUT1(
        RegA_IN), .OUT2(RegB_IN), .ADD_WR(RD4), .ADD_RD1(RS1), .ADD_RD2(RS2)
         );
  REGISTER_GENERIC_WIDTH32_10 RegA ( .CLK(CLK), .RST(n27), .EN(EN2), .DIN(
        RegA_IN), .DOUT(RegA_OUT) );
  REGISTER_GENERIC_WIDTH32_9 RegB ( .CLK(CLK), .RST(n27), .EN(EN2), .DIN(
        RegB_IN), .DOUT(RegB_OUT) );
  SIGN_EXTEND_WIDTH_IN16_WIDTH_OUT32_0 SignImm16 ( .A(IMM16), .S(SIGN_EN), .Y(
        IMMS16) );
  SIGN_EXTEND_WIDTH_IN26_WIDTH_OUT32 SignImm26 ( .A(IMM26), .S(1'b1), .Y(
        IMMS26) );
  MUX21_GENERIC_NBIT32_6 MuxIMM ( .S1(IMMS16), .S0(IMMS26), .SEL(MuxIMM_SEL), 
        .Y(IMM) );
  REGISTER_GENERIC_WIDTH32_8 RegIMM ( .CLK(CLK), .RST(n27), .EN(EN2), .DIN(IMM), .DOUT(RegIMM_OUT) );
  REGISTER_GENERIC_WIDTH5_0 RegRD2 ( .CLK(CLK), .RST(n29), .EN(EN2), .DIN(RD), 
        .DOUT(RD2) );
  REGISTER_GENERIC_WIDTH32_7 RegNPC2 ( .CLK(CLK), .RST(n27), .EN(EN2), .DIN(
        NPC1), .DOUT(NPC2) );
  MUX21_GENERIC_NBIT32_5 MuxA ( .S1(NPC2), .S0(RegA_OUT), .SEL(MuxA_SEL), .Y(
        MuxA_OUT) );
  MUX21_GENERIC_NBIT32_4 MuxB ( .S1(RegB_OUT), .S0(RegIMM_OUT), .SEL(MuxB_SEL), 
        .Y(MuxB_OUT) );
  MUX31_GENERIC_NBIT32_0 FwdA ( .S2({RegALU3_OUT, DRAM_ADDR}), .S1(MuxWB_OUT), 
        .S0(MuxA_OUT), .SEL(FwdA_SEL), .Y(A) );
  MUX31_GENERIC_NBIT32_4 FwdB ( .S2({RegALU3_OUT, DRAM_ADDR}), .S1(MuxWB_OUT), 
        .S0(MuxB_OUT), .SEL(FwdB_SEL), .Y(B) );
  ALU_WIDTH32_RADIX4 ALU0 ( .A(A), .B(B), .OP({\ALU_OPCODE[4] , 
        \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] }), 
        .Y(Y) );
  REGISTER_GENERIC_WIDTH32_6 RegALU3 ( .CLK(CLK), .RST(n28), .EN(EN3), .DIN(Y), 
        .DOUT({RegALU3_OUT, DRAM_ADDR}) );
  MUX31_GENERIC_NBIT32_3 FwdC ( .S2({RegALU3_OUT, DRAM_ADDR}), .S1(MuxWB_OUT), 
        .S0(RegA_OUT), .SEL(FwdC_SEL), .Y(Z_IN) );
  ZERO_DETECTOR_WIDTH32_0 ZERO ( .A(Z_IN), .Y(Z) );
  BRANCH_UNIT_WIDTH32 COND ( .Z(Z), .EQ_COND(EQ_COND), .JUMP_EN(JUMP_EN), 
        .BRANCH(MuxMEM_SEL) );
  REGISTER_GENERIC_WIDTH32_5 RegME ( .CLK(CLK), .RST(n28), .EN(EN3), .DIN(
        RegB_OUT), .DOUT(RegME_OUT) );
  REGISTER_GENERIC_WIDTH5_2 RegRD3 ( .CLK(CLK), .RST(n29), .EN(EN3), .DIN(RD2), 
        .DOUT(RD3) );
  REGISTER_GENERIC_WIDTH32_4 RegNPC3 ( .CLK(CLK), .RST(n28), .EN(EN3), .DIN(
        NPC2), .DOUT(NPC3) );
  SIGN_EXTEND_WIDTH_IN8_WIDTH_OUT32_0 SignLD8 ( .A(RegLMD_OUT[7:0]), .S(
        SIGN_LD_EN), .Y(LMD_8) );
  SIGN_EXTEND_WIDTH_IN16_WIDTH_OUT32_2 SignLD16 ( .A(RegLMD_OUT[15:0]), .S(
        SIGN_LD_EN), .Y(LMD_16) );
  MUX31_GENERIC_NBIT32_2 MuxLD ( .S2(LMD_8), .S1(LMD_16), .S0(RegLMD_OUT), 
        .SEL(MuxLD_SEL), .Y(MuxLD_OUT) );
  MUX21_GENERIC_NBIT32_3 MuxMEM ( .S1({RegALU3_OUT, DRAM_ADDR}), .S0(NPC3), 
        .SEL(MuxMEM_SEL), .Y(NPC_OUT) );
  MUX21_GENERIC_NBIT32_2 FwdD ( .S1(RegME_OUT), .S0(MuxWB_OUT), .SEL(FwdD_SEL), 
        .Y(MuxFWD_OUT) );
  SIGN_EXTEND_WIDTH_IN8_WIDTH_OUT32_1 SignSW8 ( .A(MuxFWD_OUT[31:24]), .S(1'b1), .Y(MEM_8) );
  SIGN_EXTEND_WIDTH_IN16_WIDTH_OUT32_1 SignSW16 ( .A(MuxFWD_OUT[31:16]), .S(
        1'b1), .Y(MEM_16) );
  MUX31_GENERIC_NBIT32_1 MuxSW ( .S2(MEM_8), .S1(MEM_16), .S0(MuxFWD_OUT), 
        .SEL(MuxSW_SEL), .Y(DRAM_OUT) );
  REGISTER_GENERIC_WIDTH32_3 RegLMD ( .CLK(CLK), .RST(n28), .EN(EN4), .DIN(
        DRAM_IN), .DOUT(RegLMD_OUT) );
  REGISTER_GENERIC_WIDTH5_1 RegRD4 ( .CLK(CLK), .RST(n29), .EN(EN4), .DIN(RD3), 
        .DOUT(RD4) );
  REGISTER_GENERIC_WIDTH32_2 RegNPC4 ( .CLK(CLK), .RST(n29), .EN(EN4), .DIN(
        NPC3), .DOUT(NPC4) );
  REGISTER_GENERIC_WIDTH32_1 RegALU4 ( .CLK(CLK), .RST(n29), .EN(EN4), .DIN({
        RegALU3_OUT, DRAM_ADDR}), .DOUT(RegALU4_OUT) );
  MUX21_GENERIC_NBIT32_1 MuxWB ( .S1(MuxLD_OUT), .S0(RegALU4_OUT), .SEL(
        MuxWB_SEL), .Y(MuxWB_OUT) );
  FORWARDING_UNIT_WIDTH32_LENGTH5 FU ( .CLK(CLK), .RST(n29), .RS1(RS1), .RS2(
        RS2), .RD3(RD3), .RD4(RD4), .RF_WE3(RF_WE3), .RF_WE4(RF_WE4), 
        .ForwardA(FwdA_SEL), .ForwardB(FwdB_SEL), .ForwardC(FwdC_SEL), 
        .ForwardD(FwdD_SEL) );
  DLX_DP_WIDTH32_LENGTH5_RADIX4_OPCODE6_DW01_add_3 add_440 ( .A(NPC4), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(
        RetADDR) );
  DLX_DP_WIDTH32_LENGTH5_RADIX4_OPCODE6_DW01_add_5 add_242 ( .A(PC_IN), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(NPC)
         );
  CLKBUF_X1 U3 ( .A(RST), .Z(n27) );
  CLKBUF_X1 U4 ( .A(RST), .Z(n28) );
  CLKBUF_X1 U5 ( .A(RST), .Z(n29) );
endmodule


module DLX_WIDTH32 ( CLK, RST, IRAM_EN, IRAM_ADDR, IRAM_DATA, DRAM_EN, DRAM_RW, 
        DRAM_ADDR, DRAM_DATA_IN, DRAM_DATA_OUT );
  output [5:0] IRAM_ADDR;
  input [31:0] IRAM_DATA;
  output [5:0] DRAM_ADDR;
  input [31:0] DRAM_DATA_IN;
  output [31:0] DRAM_DATA_OUT;
  input CLK, RST;
  output IRAM_EN, DRAM_EN, DRAM_RW;
  wire   w_EN2, w_RF_RD1, w_RF_RD2, w_MuxIMM_SEL, w_SIGN_EN, w_EN3, w_MuxA_SEL,
         w_MuxB_SEL, w_EQ_COND, w_JUMP_EN, w_RF_WE3, w_RF_WE4, w_SIGN_LD_EN,
         w_MuxWB_SEL, w_RF_WE, w_JUMP_LINK, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221;
  wire   [31:0] w_PC_IN;
  wire   [31:6] w_PC_OUT;
  wire   [31:0] w_IR_OUT;
  wire   [4:0] w_ALU_OPCODE;
  wire   [2:0] w_MuxLD_SEL;
  wire   [2:0] w_MuxSW_SEL;
  wire   [4:0] w_RD;
  wire   [4:0] w_RS2;
  wire   [15:0] w_IMM16;

  NOR4_X2 U248 ( .A1(n221), .A2(w_IR_OUT[26]), .A3(w_IR_OUT[27]), .A4(
        w_IR_OUT[30]), .ZN(n205) );
  REGISTER_GENERIC_WIDTH32_0 PC ( .CLK(CLK), .RST(RST), .EN(IRAM_EN), .DIN(
        w_PC_IN), .DOUT({w_PC_OUT, IRAM_ADDR}) );
  REGISTER_GENERIC_WIDTH32_12 IR ( .CLK(CLK), .RST(RST), .EN(IRAM_EN), .DIN(
        IRAM_DATA), .DOUT(w_IR_OUT) );
  DLX_CU_WIDTH32_LENGTH5 CU ( .CLK(CLK), .RST(RST), .IR_IN(w_IR_OUT), .EN1(
        IRAM_EN), .EN2(w_EN2), .RF_RD1(w_RF_RD1), .RF_RD2(w_RF_RD2), 
        .MuxIMM_SEL(w_MuxIMM_SEL), .SIGN_EN(w_SIGN_EN), .EN3(w_EN3), 
        .MuxA_SEL(w_MuxA_SEL), .MuxB_SEL(w_MuxB_SEL), .EQ_COND(w_EQ_COND), 
        .JUMP_EN(w_JUMP_EN), .RF_WE3(w_RF_WE3), .ALU_OPCODE(w_ALU_OPCODE), 
        .EN4(DRAM_EN), .RF_WE4(w_RF_WE4), .DRAM_WE(DRAM_RW), .SIGN_LD_EN(
        w_SIGN_LD_EN), .MuxLD_SEL(w_MuxLD_SEL), .MuxSW_SEL(w_MuxSW_SEL), 
        .MuxWB_SEL(w_MuxWB_SEL), .RF_WE(w_RF_WE), .JUMP_LINK(w_JUMP_LINK) );
  DLX_DP_WIDTH32_LENGTH5_RADIX4_OPCODE6 DP ( .CLK(CLK), .RST(RST), .EN1(
        IRAM_EN), .PC_IN({w_PC_OUT, IRAM_ADDR}), .EN2(w_EN2), .RF_RD1(w_RF_RD1), .RF_RD2(w_RF_RD2), .MuxIMM_SEL(w_MuxIMM_SEL), .SIGN_EN(w_SIGN_EN), .RD(w_RD), 
        .RS1(w_IR_OUT[25:21]), .RS2(w_RS2), .IMM16(w_IMM16), .IMM26(
        w_IR_OUT[25:0]), .EN3(w_EN3), .MuxA_SEL(w_MuxA_SEL), .MuxB_SEL(
        w_MuxB_SEL), .EQ_COND(w_EQ_COND), .JUMP_EN(w_JUMP_EN), .RF_WE3(
        w_RF_WE3), .ALU_OPCODE(w_ALU_OPCODE), .EN4(DRAM_EN), .RF_WE4(w_RF_WE4), 
        .SIGN_LD_EN(w_SIGN_LD_EN), .MuxLD_SEL(w_MuxLD_SEL), .MuxSW_SEL(
        w_MuxSW_SEL), .NPC_OUT(w_PC_IN), .DRAM_ADDR(DRAM_ADDR), .DRAM_IN(
        DRAM_DATA_IN), .DRAM_OUT(DRAM_DATA_OUT), .MuxWB_SEL(w_MuxWB_SEL), 
        .RF_WE(w_RF_WE), .JUMP_LINK(w_JUMP_LINK) );
  NOR2_X1 U281 ( .A1(n202), .A2(n211), .ZN(w_RS2[4]) );
  NOR2_X1 U282 ( .A1(n202), .A2(n212), .ZN(w_RS2[3]) );
  NOR2_X1 U283 ( .A1(n202), .A2(n215), .ZN(w_RS2[0]) );
  NOR2_X1 U284 ( .A1(n202), .A2(n213), .ZN(w_RS2[2]) );
  NOR2_X1 U285 ( .A1(n202), .A2(n214), .ZN(w_RS2[1]) );
  INV_X1 U286 ( .A(n205), .ZN(n208) );
  INV_X1 U287 ( .A(n206), .ZN(n209) );
  NOR2_X1 U288 ( .A1(n209), .A2(n216), .ZN(w_IMM16[15]) );
  NOR2_X1 U289 ( .A1(n209), .A2(n220), .ZN(w_IMM16[11]) );
  NOR2_X1 U290 ( .A1(n209), .A2(n219), .ZN(w_IMM16[12]) );
  NOR2_X1 U291 ( .A1(n209), .A2(n218), .ZN(w_IMM16[13]) );
  NOR2_X1 U292 ( .A1(n209), .A2(n217), .ZN(w_IMM16[14]) );
  INV_X1 U293 ( .A(n207), .ZN(n221) );
  NOR3_X1 U294 ( .A1(w_IR_OUT[29]), .A2(w_IR_OUT[31]), .A3(w_IR_OUT[28]), .ZN(
        n207) );
  AND2_X1 U295 ( .A1(n203), .A2(n208), .ZN(n202) );
  NAND4_X1 U296 ( .A1(w_IR_OUT[29]), .A2(w_IR_OUT[27]), .A3(w_IR_OUT[31]), 
        .A4(n204), .ZN(n203) );
  NOR3_X1 U297 ( .A1(n210), .A2(w_IR_OUT[30]), .A3(w_IR_OUT[28]), .ZN(n204) );
  INV_X1 U298 ( .A(w_IR_OUT[26]), .ZN(n210) );
  NAND3_X1 U299 ( .A1(w_IR_OUT[26]), .A2(n207), .A3(w_IR_OUT[27]), .ZN(n206)
         );
  OAI221_X1 U300 ( .B1(n205), .B2(n215), .C1(n208), .C2(n220), .A(n206), .ZN(
        w_RD[0]) );
  OAI221_X1 U301 ( .B1(n205), .B2(n214), .C1(n208), .C2(n219), .A(n206), .ZN(
        w_RD[1]) );
  OAI221_X1 U302 ( .B1(n205), .B2(n213), .C1(n208), .C2(n218), .A(n206), .ZN(
        w_RD[2]) );
  OAI221_X1 U303 ( .B1(n205), .B2(n212), .C1(n208), .C2(n217), .A(n206), .ZN(
        w_RD[3]) );
  OAI221_X1 U304 ( .B1(n205), .B2(n211), .C1(n208), .C2(n216), .A(n206), .ZN(
        w_RD[4]) );
  INV_X1 U305 ( .A(w_IR_OUT[11]), .ZN(n220) );
  INV_X1 U306 ( .A(w_IR_OUT[12]), .ZN(n219) );
  INV_X1 U307 ( .A(w_IR_OUT[13]), .ZN(n218) );
  INV_X1 U308 ( .A(w_IR_OUT[14]), .ZN(n217) );
  INV_X1 U309 ( .A(w_IR_OUT[15]), .ZN(n216) );
  INV_X1 U310 ( .A(w_IR_OUT[16]), .ZN(n215) );
  INV_X1 U311 ( .A(w_IR_OUT[17]), .ZN(n214) );
  INV_X1 U312 ( .A(w_IR_OUT[18]), .ZN(n213) );
  INV_X1 U313 ( .A(w_IR_OUT[19]), .ZN(n212) );
  INV_X1 U314 ( .A(w_IR_OUT[20]), .ZN(n211) );
  AND2_X1 U315 ( .A1(w_IR_OUT[2]), .A2(n206), .ZN(w_IMM16[2]) );
  AND2_X1 U316 ( .A1(w_IR_OUT[0]), .A2(n206), .ZN(w_IMM16[0]) );
  AND2_X1 U317 ( .A1(w_IR_OUT[1]), .A2(n206), .ZN(w_IMM16[1]) );
  AND2_X1 U318 ( .A1(w_IR_OUT[3]), .A2(n206), .ZN(w_IMM16[3]) );
  AND2_X1 U319 ( .A1(w_IR_OUT[4]), .A2(n206), .ZN(w_IMM16[4]) );
  AND2_X1 U320 ( .A1(w_IR_OUT[5]), .A2(n206), .ZN(w_IMM16[5]) );
  AND2_X1 U321 ( .A1(w_IR_OUT[6]), .A2(n206), .ZN(w_IMM16[6]) );
  AND2_X1 U322 ( .A1(w_IR_OUT[7]), .A2(n206), .ZN(w_IMM16[7]) );
  AND2_X1 U323 ( .A1(w_IR_OUT[8]), .A2(n206), .ZN(w_IMM16[8]) );
  AND2_X1 U324 ( .A1(w_IR_OUT[9]), .A2(n206), .ZN(w_IMM16[9]) );
  AND2_X1 U325 ( .A1(w_IR_OUT[10]), .A2(n206), .ZN(w_IMM16[10]) );
endmodule


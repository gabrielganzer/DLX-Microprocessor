
module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_0 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_31 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_30 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_29 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_28 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_27 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_26 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_25 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_24 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_23 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_22 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_21 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_20 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_19 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_18 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_17 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_16 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_15 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_14 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_13 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_12 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_11 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_10 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_9 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_8 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_7 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_6 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_5 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_4 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_3 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_2 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_1 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2386, net2388, net2390, net2391, net2394, net2397;
  assign net2386 = EN;
  assign net2388 = CLK;
  assign ENCLK = net2390;
  assign net2397 = TE;

  DLL_X1 latch ( .D(net2391), .GN(net2388), .Q(net2394) );
  OR2_X1 test_or ( .A1(net2386), .A2(net2397), .ZN(net2391) );
  AND2_X1 main_gate ( .A1(net2394), .A2(net2388), .ZN(net2390) );
endmodule


module REGISTER_FILE_WIDTH32_LENGTH5 ( CLK, RST, EN, RD1, RD2, WR, DATAIN, 
        OUT1, OUT2, ADD_WR, ADD_RD1, ADD_RD2 );
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input CLK, RST, EN, RD1, RD2, WR;
  wire   \REGISTERS[0][31] , \REGISTERS[0][30] , \REGISTERS[0][29] ,
         \REGISTERS[0][28] , \REGISTERS[0][27] , \REGISTERS[0][26] ,
         \REGISTERS[0][25] , \REGISTERS[0][24] , \REGISTERS[0][23] ,
         \REGISTERS[0][22] , \REGISTERS[0][21] , \REGISTERS[0][20] ,
         \REGISTERS[0][19] , \REGISTERS[0][18] , \REGISTERS[0][17] ,
         \REGISTERS[0][16] , \REGISTERS[0][15] , \REGISTERS[0][14] ,
         \REGISTERS[0][13] , \REGISTERS[0][12] , \REGISTERS[0][11] ,
         \REGISTERS[0][10] , \REGISTERS[0][9] , \REGISTERS[0][8] ,
         \REGISTERS[0][7] , \REGISTERS[0][6] , \REGISTERS[0][5] ,
         \REGISTERS[0][4] , \REGISTERS[0][3] , \REGISTERS[0][2] ,
         \REGISTERS[0][1] , \REGISTERS[0][0] , \REGISTERS[1][31] ,
         \REGISTERS[1][30] , \REGISTERS[1][29] , \REGISTERS[1][28] ,
         \REGISTERS[1][27] , \REGISTERS[1][26] , \REGISTERS[1][25] ,
         \REGISTERS[1][24] , \REGISTERS[1][23] , \REGISTERS[1][22] ,
         \REGISTERS[1][21] , \REGISTERS[1][20] , \REGISTERS[1][19] ,
         \REGISTERS[1][18] , \REGISTERS[1][17] , \REGISTERS[1][16] ,
         \REGISTERS[1][15] , \REGISTERS[1][14] , \REGISTERS[1][13] ,
         \REGISTERS[1][12] , \REGISTERS[1][11] , \REGISTERS[1][10] ,
         \REGISTERS[1][9] , \REGISTERS[1][8] , \REGISTERS[1][7] ,
         \REGISTERS[1][6] , \REGISTERS[1][5] , \REGISTERS[1][4] ,
         \REGISTERS[1][3] , \REGISTERS[1][2] , \REGISTERS[1][1] ,
         \REGISTERS[1][0] , \REGISTERS[2][31] , \REGISTERS[2][30] ,
         \REGISTERS[2][29] , \REGISTERS[2][28] , \REGISTERS[2][27] ,
         \REGISTERS[2][26] , \REGISTERS[2][25] , \REGISTERS[2][24] ,
         \REGISTERS[2][23] , \REGISTERS[2][22] , \REGISTERS[2][21] ,
         \REGISTERS[2][20] , \REGISTERS[2][19] , \REGISTERS[2][18] ,
         \REGISTERS[2][17] , \REGISTERS[2][16] , \REGISTERS[2][15] ,
         \REGISTERS[2][14] , \REGISTERS[2][13] , \REGISTERS[2][12] ,
         \REGISTERS[2][11] , \REGISTERS[2][10] , \REGISTERS[2][9] ,
         \REGISTERS[2][8] , \REGISTERS[2][7] , \REGISTERS[2][6] ,
         \REGISTERS[2][5] , \REGISTERS[2][4] , \REGISTERS[2][3] ,
         \REGISTERS[2][2] , \REGISTERS[2][1] , \REGISTERS[2][0] ,
         \REGISTERS[3][31] , \REGISTERS[3][30] , \REGISTERS[3][29] ,
         \REGISTERS[3][28] , \REGISTERS[3][27] , \REGISTERS[3][26] ,
         \REGISTERS[3][25] , \REGISTERS[3][24] , \REGISTERS[3][23] ,
         \REGISTERS[3][22] , \REGISTERS[3][21] , \REGISTERS[3][20] ,
         \REGISTERS[3][19] , \REGISTERS[3][18] , \REGISTERS[3][17] ,
         \REGISTERS[3][16] , \REGISTERS[3][15] , \REGISTERS[3][14] ,
         \REGISTERS[3][13] , \REGISTERS[3][12] , \REGISTERS[3][11] ,
         \REGISTERS[3][10] , \REGISTERS[3][9] , \REGISTERS[3][8] ,
         \REGISTERS[3][7] , \REGISTERS[3][6] , \REGISTERS[3][5] ,
         \REGISTERS[3][4] , \REGISTERS[3][3] , \REGISTERS[3][2] ,
         \REGISTERS[3][1] , \REGISTERS[3][0] , \REGISTERS[4][31] ,
         \REGISTERS[4][30] , \REGISTERS[4][29] , \REGISTERS[4][28] ,
         \REGISTERS[4][27] , \REGISTERS[4][26] , \REGISTERS[4][25] ,
         \REGISTERS[4][24] , \REGISTERS[4][23] , \REGISTERS[4][22] ,
         \REGISTERS[4][21] , \REGISTERS[4][20] , \REGISTERS[4][19] ,
         \REGISTERS[4][18] , \REGISTERS[4][17] , \REGISTERS[4][16] ,
         \REGISTERS[4][15] , \REGISTERS[4][14] , \REGISTERS[4][13] ,
         \REGISTERS[4][12] , \REGISTERS[4][11] , \REGISTERS[4][10] ,
         \REGISTERS[4][9] , \REGISTERS[4][8] , \REGISTERS[4][7] ,
         \REGISTERS[4][6] , \REGISTERS[4][5] , \REGISTERS[4][4] ,
         \REGISTERS[4][3] , \REGISTERS[4][2] , \REGISTERS[4][1] ,
         \REGISTERS[4][0] , \REGISTERS[5][31] , \REGISTERS[5][30] ,
         \REGISTERS[5][29] , \REGISTERS[5][28] , \REGISTERS[5][27] ,
         \REGISTERS[5][26] , \REGISTERS[5][25] , \REGISTERS[5][24] ,
         \REGISTERS[5][23] , \REGISTERS[5][22] , \REGISTERS[5][21] ,
         \REGISTERS[5][20] , \REGISTERS[5][19] , \REGISTERS[5][18] ,
         \REGISTERS[5][17] , \REGISTERS[5][16] , \REGISTERS[5][15] ,
         \REGISTERS[5][14] , \REGISTERS[5][13] , \REGISTERS[5][12] ,
         \REGISTERS[5][11] , \REGISTERS[5][10] , \REGISTERS[5][9] ,
         \REGISTERS[5][8] , \REGISTERS[5][7] , \REGISTERS[5][6] ,
         \REGISTERS[5][5] , \REGISTERS[5][4] , \REGISTERS[5][3] ,
         \REGISTERS[5][2] , \REGISTERS[5][1] , \REGISTERS[5][0] ,
         \REGISTERS[6][31] , \REGISTERS[6][30] , \REGISTERS[6][29] ,
         \REGISTERS[6][28] , \REGISTERS[6][27] , \REGISTERS[6][26] ,
         \REGISTERS[6][25] , \REGISTERS[6][24] , \REGISTERS[6][23] ,
         \REGISTERS[6][22] , \REGISTERS[6][21] , \REGISTERS[6][20] ,
         \REGISTERS[6][19] , \REGISTERS[6][18] , \REGISTERS[6][17] ,
         \REGISTERS[6][16] , \REGISTERS[6][15] , \REGISTERS[6][14] ,
         \REGISTERS[6][13] , \REGISTERS[6][12] , \REGISTERS[6][11] ,
         \REGISTERS[6][10] , \REGISTERS[6][9] , \REGISTERS[6][8] ,
         \REGISTERS[6][7] , \REGISTERS[6][6] , \REGISTERS[6][5] ,
         \REGISTERS[6][4] , \REGISTERS[6][3] , \REGISTERS[6][2] ,
         \REGISTERS[6][1] , \REGISTERS[6][0] , \REGISTERS[7][31] ,
         \REGISTERS[7][30] , \REGISTERS[7][29] , \REGISTERS[7][28] ,
         \REGISTERS[7][27] , \REGISTERS[7][26] , \REGISTERS[7][25] ,
         \REGISTERS[7][24] , \REGISTERS[7][23] , \REGISTERS[7][22] ,
         \REGISTERS[7][21] , \REGISTERS[7][20] , \REGISTERS[7][19] ,
         \REGISTERS[7][18] , \REGISTERS[7][17] , \REGISTERS[7][16] ,
         \REGISTERS[7][15] , \REGISTERS[7][14] , \REGISTERS[7][13] ,
         \REGISTERS[7][12] , \REGISTERS[7][11] , \REGISTERS[7][10] ,
         \REGISTERS[7][9] , \REGISTERS[7][8] , \REGISTERS[7][7] ,
         \REGISTERS[7][6] , \REGISTERS[7][5] , \REGISTERS[7][4] ,
         \REGISTERS[7][3] , \REGISTERS[7][2] , \REGISTERS[7][1] ,
         \REGISTERS[7][0] , \REGISTERS[8][31] , \REGISTERS[8][30] ,
         \REGISTERS[8][29] , \REGISTERS[8][28] , \REGISTERS[8][27] ,
         \REGISTERS[8][26] , \REGISTERS[8][25] , \REGISTERS[8][24] ,
         \REGISTERS[8][23] , \REGISTERS[8][22] , \REGISTERS[8][21] ,
         \REGISTERS[8][20] , \REGISTERS[8][19] , \REGISTERS[8][18] ,
         \REGISTERS[8][17] , \REGISTERS[8][16] , \REGISTERS[8][15] ,
         \REGISTERS[8][14] , \REGISTERS[8][13] , \REGISTERS[8][12] ,
         \REGISTERS[8][11] , \REGISTERS[8][10] , \REGISTERS[8][9] ,
         \REGISTERS[8][8] , \REGISTERS[8][7] , \REGISTERS[8][6] ,
         \REGISTERS[8][5] , \REGISTERS[8][4] , \REGISTERS[8][3] ,
         \REGISTERS[8][2] , \REGISTERS[8][1] , \REGISTERS[8][0] ,
         \REGISTERS[9][31] , \REGISTERS[9][30] , \REGISTERS[9][29] ,
         \REGISTERS[9][28] , \REGISTERS[9][27] , \REGISTERS[9][26] ,
         \REGISTERS[9][25] , \REGISTERS[9][24] , \REGISTERS[9][23] ,
         \REGISTERS[9][22] , \REGISTERS[9][21] , \REGISTERS[9][20] ,
         \REGISTERS[9][19] , \REGISTERS[9][18] , \REGISTERS[9][17] ,
         \REGISTERS[9][16] , \REGISTERS[9][15] , \REGISTERS[9][14] ,
         \REGISTERS[9][13] , \REGISTERS[9][12] , \REGISTERS[9][11] ,
         \REGISTERS[9][10] , \REGISTERS[9][9] , \REGISTERS[9][8] ,
         \REGISTERS[9][7] , \REGISTERS[9][6] , \REGISTERS[9][5] ,
         \REGISTERS[9][4] , \REGISTERS[9][3] , \REGISTERS[9][2] ,
         \REGISTERS[9][1] , \REGISTERS[9][0] , \REGISTERS[10][31] ,
         \REGISTERS[10][30] , \REGISTERS[10][29] , \REGISTERS[10][28] ,
         \REGISTERS[10][27] , \REGISTERS[10][26] , \REGISTERS[10][25] ,
         \REGISTERS[10][24] , \REGISTERS[10][23] , \REGISTERS[10][22] ,
         \REGISTERS[10][21] , \REGISTERS[10][20] , \REGISTERS[10][19] ,
         \REGISTERS[10][18] , \REGISTERS[10][17] , \REGISTERS[10][16] ,
         \REGISTERS[10][15] , \REGISTERS[10][14] , \REGISTERS[10][13] ,
         \REGISTERS[10][12] , \REGISTERS[10][11] , \REGISTERS[10][10] ,
         \REGISTERS[10][9] , \REGISTERS[10][8] , \REGISTERS[10][7] ,
         \REGISTERS[10][6] , \REGISTERS[10][5] , \REGISTERS[10][4] ,
         \REGISTERS[10][3] , \REGISTERS[10][2] , \REGISTERS[10][1] ,
         \REGISTERS[10][0] , \REGISTERS[11][31] , \REGISTERS[11][30] ,
         \REGISTERS[11][29] , \REGISTERS[11][28] , \REGISTERS[11][27] ,
         \REGISTERS[11][26] , \REGISTERS[11][25] , \REGISTERS[11][24] ,
         \REGISTERS[11][23] , \REGISTERS[11][22] , \REGISTERS[11][21] ,
         \REGISTERS[11][20] , \REGISTERS[11][19] , \REGISTERS[11][18] ,
         \REGISTERS[11][17] , \REGISTERS[11][16] , \REGISTERS[11][15] ,
         \REGISTERS[11][14] , \REGISTERS[11][13] , \REGISTERS[11][12] ,
         \REGISTERS[11][11] , \REGISTERS[11][10] , \REGISTERS[11][9] ,
         \REGISTERS[11][8] , \REGISTERS[11][7] , \REGISTERS[11][6] ,
         \REGISTERS[11][5] , \REGISTERS[11][4] , \REGISTERS[11][3] ,
         \REGISTERS[11][2] , \REGISTERS[11][1] , \REGISTERS[11][0] ,
         \REGISTERS[12][31] , \REGISTERS[12][30] , \REGISTERS[12][29] ,
         \REGISTERS[12][28] , \REGISTERS[12][27] , \REGISTERS[12][26] ,
         \REGISTERS[12][25] , \REGISTERS[12][24] , \REGISTERS[12][23] ,
         \REGISTERS[12][22] , \REGISTERS[12][21] , \REGISTERS[12][20] ,
         \REGISTERS[12][19] , \REGISTERS[12][18] , \REGISTERS[12][17] ,
         \REGISTERS[12][16] , \REGISTERS[12][15] , \REGISTERS[12][14] ,
         \REGISTERS[12][13] , \REGISTERS[12][12] , \REGISTERS[12][11] ,
         \REGISTERS[12][10] , \REGISTERS[12][9] , \REGISTERS[12][8] ,
         \REGISTERS[12][7] , \REGISTERS[12][6] , \REGISTERS[12][5] ,
         \REGISTERS[12][4] , \REGISTERS[12][3] , \REGISTERS[12][2] ,
         \REGISTERS[12][1] , \REGISTERS[12][0] , \REGISTERS[13][31] ,
         \REGISTERS[13][30] , \REGISTERS[13][29] , \REGISTERS[13][28] ,
         \REGISTERS[13][27] , \REGISTERS[13][26] , \REGISTERS[13][25] ,
         \REGISTERS[13][24] , \REGISTERS[13][23] , \REGISTERS[13][22] ,
         \REGISTERS[13][21] , \REGISTERS[13][20] , \REGISTERS[13][19] ,
         \REGISTERS[13][18] , \REGISTERS[13][17] , \REGISTERS[13][16] ,
         \REGISTERS[13][15] , \REGISTERS[13][14] , \REGISTERS[13][13] ,
         \REGISTERS[13][12] , \REGISTERS[13][11] , \REGISTERS[13][10] ,
         \REGISTERS[13][9] , \REGISTERS[13][8] , \REGISTERS[13][7] ,
         \REGISTERS[13][6] , \REGISTERS[13][5] , \REGISTERS[13][4] ,
         \REGISTERS[13][3] , \REGISTERS[13][2] , \REGISTERS[13][1] ,
         \REGISTERS[13][0] , \REGISTERS[14][31] , \REGISTERS[14][30] ,
         \REGISTERS[14][29] , \REGISTERS[14][28] , \REGISTERS[14][27] ,
         \REGISTERS[14][26] , \REGISTERS[14][25] , \REGISTERS[14][24] ,
         \REGISTERS[14][23] , \REGISTERS[14][22] , \REGISTERS[14][21] ,
         \REGISTERS[14][20] , \REGISTERS[14][19] , \REGISTERS[14][18] ,
         \REGISTERS[14][17] , \REGISTERS[14][16] , \REGISTERS[14][15] ,
         \REGISTERS[14][14] , \REGISTERS[14][13] , \REGISTERS[14][12] ,
         \REGISTERS[14][11] , \REGISTERS[14][10] , \REGISTERS[14][9] ,
         \REGISTERS[14][8] , \REGISTERS[14][7] , \REGISTERS[14][6] ,
         \REGISTERS[14][5] , \REGISTERS[14][4] , \REGISTERS[14][3] ,
         \REGISTERS[14][2] , \REGISTERS[14][1] , \REGISTERS[14][0] ,
         \REGISTERS[15][31] , \REGISTERS[15][30] , \REGISTERS[15][29] ,
         \REGISTERS[15][28] , \REGISTERS[15][27] , \REGISTERS[15][26] ,
         \REGISTERS[15][25] , \REGISTERS[15][24] , \REGISTERS[15][23] ,
         \REGISTERS[15][22] , \REGISTERS[15][21] , \REGISTERS[15][20] ,
         \REGISTERS[15][19] , \REGISTERS[15][18] , \REGISTERS[15][17] ,
         \REGISTERS[15][16] , \REGISTERS[15][15] , \REGISTERS[15][14] ,
         \REGISTERS[15][13] , \REGISTERS[15][12] , \REGISTERS[15][11] ,
         \REGISTERS[15][10] , \REGISTERS[15][9] , \REGISTERS[15][8] ,
         \REGISTERS[15][7] , \REGISTERS[15][6] , \REGISTERS[15][5] ,
         \REGISTERS[15][4] , \REGISTERS[15][3] , \REGISTERS[15][2] ,
         \REGISTERS[15][1] , \REGISTERS[15][0] , \REGISTERS[16][31] ,
         \REGISTERS[16][30] , \REGISTERS[16][29] , \REGISTERS[16][28] ,
         \REGISTERS[16][27] , \REGISTERS[16][26] , \REGISTERS[16][25] ,
         \REGISTERS[16][24] , \REGISTERS[16][23] , \REGISTERS[16][22] ,
         \REGISTERS[16][21] , \REGISTERS[16][20] , \REGISTERS[16][19] ,
         \REGISTERS[16][18] , \REGISTERS[16][17] , \REGISTERS[16][16] ,
         \REGISTERS[16][15] , \REGISTERS[16][14] , \REGISTERS[16][13] ,
         \REGISTERS[16][12] , \REGISTERS[16][11] , \REGISTERS[16][10] ,
         \REGISTERS[16][9] , \REGISTERS[16][8] , \REGISTERS[16][7] ,
         \REGISTERS[16][6] , \REGISTERS[16][5] , \REGISTERS[16][4] ,
         \REGISTERS[16][3] , \REGISTERS[16][2] , \REGISTERS[16][1] ,
         \REGISTERS[16][0] , \REGISTERS[17][31] , \REGISTERS[17][30] ,
         \REGISTERS[17][29] , \REGISTERS[17][28] , \REGISTERS[17][27] ,
         \REGISTERS[17][26] , \REGISTERS[17][25] , \REGISTERS[17][24] ,
         \REGISTERS[17][23] , \REGISTERS[17][22] , \REGISTERS[17][21] ,
         \REGISTERS[17][20] , \REGISTERS[17][19] , \REGISTERS[17][18] ,
         \REGISTERS[17][17] , \REGISTERS[17][16] , \REGISTERS[17][15] ,
         \REGISTERS[17][14] , \REGISTERS[17][13] , \REGISTERS[17][12] ,
         \REGISTERS[17][11] , \REGISTERS[17][10] , \REGISTERS[17][9] ,
         \REGISTERS[17][8] , \REGISTERS[17][7] , \REGISTERS[17][6] ,
         \REGISTERS[17][5] , \REGISTERS[17][4] , \REGISTERS[17][3] ,
         \REGISTERS[17][2] , \REGISTERS[17][1] , \REGISTERS[17][0] ,
         \REGISTERS[18][31] , \REGISTERS[18][30] , \REGISTERS[18][29] ,
         \REGISTERS[18][28] , \REGISTERS[18][27] , \REGISTERS[18][26] ,
         \REGISTERS[18][25] , \REGISTERS[18][24] , \REGISTERS[18][23] ,
         \REGISTERS[18][22] , \REGISTERS[18][21] , \REGISTERS[18][20] ,
         \REGISTERS[18][19] , \REGISTERS[18][18] , \REGISTERS[18][17] ,
         \REGISTERS[18][16] , \REGISTERS[18][15] , \REGISTERS[18][14] ,
         \REGISTERS[18][13] , \REGISTERS[18][12] , \REGISTERS[18][11] ,
         \REGISTERS[18][10] , \REGISTERS[18][9] , \REGISTERS[18][8] ,
         \REGISTERS[18][7] , \REGISTERS[18][6] , \REGISTERS[18][5] ,
         \REGISTERS[18][4] , \REGISTERS[18][3] , \REGISTERS[18][2] ,
         \REGISTERS[18][1] , \REGISTERS[18][0] , \REGISTERS[19][31] ,
         \REGISTERS[19][30] , \REGISTERS[19][29] , \REGISTERS[19][28] ,
         \REGISTERS[19][27] , \REGISTERS[19][26] , \REGISTERS[19][25] ,
         \REGISTERS[19][24] , \REGISTERS[19][23] , \REGISTERS[19][22] ,
         \REGISTERS[19][21] , \REGISTERS[19][20] , \REGISTERS[19][19] ,
         \REGISTERS[19][18] , \REGISTERS[19][17] , \REGISTERS[19][16] ,
         \REGISTERS[19][15] , \REGISTERS[19][14] , \REGISTERS[19][13] ,
         \REGISTERS[19][12] , \REGISTERS[19][11] , \REGISTERS[19][10] ,
         \REGISTERS[19][9] , \REGISTERS[19][8] , \REGISTERS[19][7] ,
         \REGISTERS[19][6] , \REGISTERS[19][5] , \REGISTERS[19][4] ,
         \REGISTERS[19][3] , \REGISTERS[19][2] , \REGISTERS[19][1] ,
         \REGISTERS[19][0] , \REGISTERS[20][31] , \REGISTERS[20][30] ,
         \REGISTERS[20][29] , \REGISTERS[20][28] , \REGISTERS[20][27] ,
         \REGISTERS[20][26] , \REGISTERS[20][25] , \REGISTERS[20][24] ,
         \REGISTERS[20][23] , \REGISTERS[20][22] , \REGISTERS[20][21] ,
         \REGISTERS[20][20] , \REGISTERS[20][19] , \REGISTERS[20][18] ,
         \REGISTERS[20][17] , \REGISTERS[20][16] , \REGISTERS[20][15] ,
         \REGISTERS[20][14] , \REGISTERS[20][13] , \REGISTERS[20][12] ,
         \REGISTERS[20][11] , \REGISTERS[20][10] , \REGISTERS[20][9] ,
         \REGISTERS[20][8] , \REGISTERS[20][7] , \REGISTERS[20][6] ,
         \REGISTERS[20][5] , \REGISTERS[20][4] , \REGISTERS[20][3] ,
         \REGISTERS[20][2] , \REGISTERS[20][1] , \REGISTERS[20][0] ,
         \REGISTERS[21][31] , \REGISTERS[21][30] , \REGISTERS[21][29] ,
         \REGISTERS[21][28] , \REGISTERS[21][27] , \REGISTERS[21][26] ,
         \REGISTERS[21][25] , \REGISTERS[21][24] , \REGISTERS[21][23] ,
         \REGISTERS[21][22] , \REGISTERS[21][21] , \REGISTERS[21][20] ,
         \REGISTERS[21][19] , \REGISTERS[21][18] , \REGISTERS[21][17] ,
         \REGISTERS[21][16] , \REGISTERS[21][15] , \REGISTERS[21][14] ,
         \REGISTERS[21][13] , \REGISTERS[21][12] , \REGISTERS[21][11] ,
         \REGISTERS[21][10] , \REGISTERS[21][9] , \REGISTERS[21][8] ,
         \REGISTERS[21][7] , \REGISTERS[21][6] , \REGISTERS[21][5] ,
         \REGISTERS[21][4] , \REGISTERS[21][3] , \REGISTERS[21][2] ,
         \REGISTERS[21][1] , \REGISTERS[21][0] , \REGISTERS[22][31] ,
         \REGISTERS[22][30] , \REGISTERS[22][29] , \REGISTERS[22][28] ,
         \REGISTERS[22][27] , \REGISTERS[22][26] , \REGISTERS[22][25] ,
         \REGISTERS[22][24] , \REGISTERS[22][23] , \REGISTERS[22][22] ,
         \REGISTERS[22][21] , \REGISTERS[22][20] , \REGISTERS[22][19] ,
         \REGISTERS[22][18] , \REGISTERS[22][17] , \REGISTERS[22][16] ,
         \REGISTERS[22][15] , \REGISTERS[22][14] , \REGISTERS[22][13] ,
         \REGISTERS[22][12] , \REGISTERS[22][11] , \REGISTERS[22][10] ,
         \REGISTERS[22][9] , \REGISTERS[22][8] , \REGISTERS[22][7] ,
         \REGISTERS[22][6] , \REGISTERS[22][5] , \REGISTERS[22][4] ,
         \REGISTERS[22][3] , \REGISTERS[22][2] , \REGISTERS[22][1] ,
         \REGISTERS[22][0] , \REGISTERS[23][31] , \REGISTERS[23][30] ,
         \REGISTERS[23][29] , \REGISTERS[23][28] , \REGISTERS[23][27] ,
         \REGISTERS[23][26] , \REGISTERS[23][25] , \REGISTERS[23][24] ,
         \REGISTERS[23][23] , \REGISTERS[23][22] , \REGISTERS[23][21] ,
         \REGISTERS[23][20] , \REGISTERS[23][19] , \REGISTERS[23][18] ,
         \REGISTERS[23][17] , \REGISTERS[23][16] , \REGISTERS[23][15] ,
         \REGISTERS[23][14] , \REGISTERS[23][13] , \REGISTERS[23][12] ,
         \REGISTERS[23][11] , \REGISTERS[23][10] , \REGISTERS[23][9] ,
         \REGISTERS[23][8] , \REGISTERS[23][7] , \REGISTERS[23][6] ,
         \REGISTERS[23][5] , \REGISTERS[23][4] , \REGISTERS[23][3] ,
         \REGISTERS[23][2] , \REGISTERS[23][1] , \REGISTERS[23][0] ,
         \REGISTERS[24][31] , \REGISTERS[24][30] , \REGISTERS[24][29] ,
         \REGISTERS[24][28] , \REGISTERS[24][27] , \REGISTERS[24][26] ,
         \REGISTERS[24][25] , \REGISTERS[24][24] , \REGISTERS[24][23] ,
         \REGISTERS[24][22] , \REGISTERS[24][21] , \REGISTERS[24][20] ,
         \REGISTERS[24][19] , \REGISTERS[24][18] , \REGISTERS[24][17] ,
         \REGISTERS[24][16] , \REGISTERS[24][15] , \REGISTERS[24][14] ,
         \REGISTERS[24][13] , \REGISTERS[24][12] , \REGISTERS[24][11] ,
         \REGISTERS[24][10] , \REGISTERS[24][9] , \REGISTERS[24][8] ,
         \REGISTERS[24][7] , \REGISTERS[24][6] , \REGISTERS[24][5] ,
         \REGISTERS[24][4] , \REGISTERS[24][3] , \REGISTERS[24][2] ,
         \REGISTERS[24][1] , \REGISTERS[24][0] , \REGISTERS[25][31] ,
         \REGISTERS[25][30] , \REGISTERS[25][29] , \REGISTERS[25][28] ,
         \REGISTERS[25][27] , \REGISTERS[25][26] , \REGISTERS[25][25] ,
         \REGISTERS[25][24] , \REGISTERS[25][23] , \REGISTERS[25][22] ,
         \REGISTERS[25][21] , \REGISTERS[25][20] , \REGISTERS[25][19] ,
         \REGISTERS[25][18] , \REGISTERS[25][17] , \REGISTERS[25][16] ,
         \REGISTERS[25][15] , \REGISTERS[25][14] , \REGISTERS[25][13] ,
         \REGISTERS[25][12] , \REGISTERS[25][11] , \REGISTERS[25][10] ,
         \REGISTERS[25][9] , \REGISTERS[25][8] , \REGISTERS[25][7] ,
         \REGISTERS[25][6] , \REGISTERS[25][5] , \REGISTERS[25][4] ,
         \REGISTERS[25][3] , \REGISTERS[25][2] , \REGISTERS[25][1] ,
         \REGISTERS[25][0] , \REGISTERS[26][31] , \REGISTERS[26][30] ,
         \REGISTERS[26][29] , \REGISTERS[26][28] , \REGISTERS[26][27] ,
         \REGISTERS[26][26] , \REGISTERS[26][25] , \REGISTERS[26][24] ,
         \REGISTERS[26][23] , \REGISTERS[26][22] , \REGISTERS[26][21] ,
         \REGISTERS[26][20] , \REGISTERS[26][19] , \REGISTERS[26][18] ,
         \REGISTERS[26][17] , \REGISTERS[26][16] , \REGISTERS[26][15] ,
         \REGISTERS[26][14] , \REGISTERS[26][13] , \REGISTERS[26][12] ,
         \REGISTERS[26][11] , \REGISTERS[26][10] , \REGISTERS[26][9] ,
         \REGISTERS[26][8] , \REGISTERS[26][7] , \REGISTERS[26][6] ,
         \REGISTERS[26][5] , \REGISTERS[26][4] , \REGISTERS[26][3] ,
         \REGISTERS[26][2] , \REGISTERS[26][1] , \REGISTERS[26][0] ,
         \REGISTERS[27][31] , \REGISTERS[27][30] , \REGISTERS[27][29] ,
         \REGISTERS[27][28] , \REGISTERS[27][27] , \REGISTERS[27][26] ,
         \REGISTERS[27][25] , \REGISTERS[27][24] , \REGISTERS[27][23] ,
         \REGISTERS[27][22] , \REGISTERS[27][21] , \REGISTERS[27][20] ,
         \REGISTERS[27][19] , \REGISTERS[27][18] , \REGISTERS[27][17] ,
         \REGISTERS[27][16] , \REGISTERS[27][15] , \REGISTERS[27][14] ,
         \REGISTERS[27][13] , \REGISTERS[27][12] , \REGISTERS[27][11] ,
         \REGISTERS[27][10] , \REGISTERS[27][9] , \REGISTERS[27][8] ,
         \REGISTERS[27][7] , \REGISTERS[27][6] , \REGISTERS[27][5] ,
         \REGISTERS[27][4] , \REGISTERS[27][3] , \REGISTERS[27][2] ,
         \REGISTERS[27][1] , \REGISTERS[27][0] , \REGISTERS[28][31] ,
         \REGISTERS[28][30] , \REGISTERS[28][29] , \REGISTERS[28][28] ,
         \REGISTERS[28][27] , \REGISTERS[28][26] , \REGISTERS[28][25] ,
         \REGISTERS[28][24] , \REGISTERS[28][23] , \REGISTERS[28][22] ,
         \REGISTERS[28][21] , \REGISTERS[28][20] , \REGISTERS[28][19] ,
         \REGISTERS[28][18] , \REGISTERS[28][17] , \REGISTERS[28][16] ,
         \REGISTERS[28][15] , \REGISTERS[28][14] , \REGISTERS[28][13] ,
         \REGISTERS[28][12] , \REGISTERS[28][11] , \REGISTERS[28][10] ,
         \REGISTERS[28][9] , \REGISTERS[28][8] , \REGISTERS[28][7] ,
         \REGISTERS[28][6] , \REGISTERS[28][5] , \REGISTERS[28][4] ,
         \REGISTERS[28][3] , \REGISTERS[28][2] , \REGISTERS[28][1] ,
         \REGISTERS[28][0] , \REGISTERS[29][31] , \REGISTERS[29][30] ,
         \REGISTERS[29][29] , \REGISTERS[29][28] , \REGISTERS[29][27] ,
         \REGISTERS[29][26] , \REGISTERS[29][25] , \REGISTERS[29][24] ,
         \REGISTERS[29][23] , \REGISTERS[29][22] , \REGISTERS[29][21] ,
         \REGISTERS[29][20] , \REGISTERS[29][19] , \REGISTERS[29][18] ,
         \REGISTERS[29][17] , \REGISTERS[29][16] , \REGISTERS[29][15] ,
         \REGISTERS[29][14] , \REGISTERS[29][13] , \REGISTERS[29][12] ,
         \REGISTERS[29][11] , \REGISTERS[29][10] , \REGISTERS[29][9] ,
         \REGISTERS[29][8] , \REGISTERS[29][7] , \REGISTERS[29][6] ,
         \REGISTERS[29][5] , \REGISTERS[29][4] , \REGISTERS[29][3] ,
         \REGISTERS[29][2] , \REGISTERS[29][1] , \REGISTERS[29][0] ,
         \REGISTERS[30][31] , \REGISTERS[30][30] , \REGISTERS[30][29] ,
         \REGISTERS[30][28] , \REGISTERS[30][27] , \REGISTERS[30][26] ,
         \REGISTERS[30][25] , \REGISTERS[30][24] , \REGISTERS[30][23] ,
         \REGISTERS[30][22] , \REGISTERS[30][21] , \REGISTERS[30][20] ,
         \REGISTERS[30][19] , \REGISTERS[30][18] , \REGISTERS[30][17] ,
         \REGISTERS[30][16] , \REGISTERS[30][15] , \REGISTERS[30][14] ,
         \REGISTERS[30][13] , \REGISTERS[30][12] , \REGISTERS[30][11] ,
         \REGISTERS[30][10] , \REGISTERS[30][9] , \REGISTERS[30][8] ,
         \REGISTERS[30][7] , \REGISTERS[30][6] , \REGISTERS[30][5] ,
         \REGISTERS[30][4] , \REGISTERS[30][3] , \REGISTERS[30][2] ,
         \REGISTERS[30][1] , \REGISTERS[30][0] , \REGISTERS[31][31] ,
         \REGISTERS[31][30] , \REGISTERS[31][29] , \REGISTERS[31][28] ,
         \REGISTERS[31][27] , \REGISTERS[31][26] , \REGISTERS[31][25] ,
         \REGISTERS[31][24] , \REGISTERS[31][23] , \REGISTERS[31][22] ,
         \REGISTERS[31][21] , \REGISTERS[31][20] , \REGISTERS[31][19] ,
         \REGISTERS[31][18] , \REGISTERS[31][17] , \REGISTERS[31][16] ,
         \REGISTERS[31][15] , \REGISTERS[31][14] , \REGISTERS[31][13] ,
         \REGISTERS[31][12] , \REGISTERS[31][11] , \REGISTERS[31][10] ,
         \REGISTERS[31][9] , \REGISTERS[31][8] , \REGISTERS[31][7] ,
         \REGISTERS[31][6] , \REGISTERS[31][5] , \REGISTERS[31][4] ,
         \REGISTERS[31][3] , \REGISTERS[31][2] , \REGISTERS[31][1] ,
         \REGISTERS[31][0] , N81, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, net2402, net2408, net2413, net2418, net2423, net2428,
         net2433, net2438, net2443, net2448, net2453, net2458, net2463,
         net2468, net2473, net2478, net2483, net2488, net2493, net2498,
         net2503, net2508, net2513, net2518, net2523, net2528, net2533,
         net2538, net2543, net2548, net2553, net2558, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n107, n108, n109, n110, n111,
         n112, n113, n114, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678;

  DLH_X1 \OUT1_reg[31]  ( .G(N411), .D(N278), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(N411), .D(N277), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(N411), .D(N276), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(N411), .D(N275), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(N411), .D(N274), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(N411), .D(N273), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(N411), .D(N272), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(N411), .D(N271), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(N411), .D(N270), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(N411), .D(N269), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(N411), .D(N268), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(N411), .D(N267), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(N411), .D(N266), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(N411), .D(N265), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(N411), .D(N264), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(N411), .D(N263), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(N411), .D(N262), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(N411), .D(N261), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(N411), .D(N260), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(N411), .D(N259), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(N411), .D(N258), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(N411), .D(N257), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(N411), .D(N256), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(N411), .D(N255), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(N411), .D(N254), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(N411), .D(N253), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(N411), .D(N252), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(N411), .D(N251), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(N411), .D(N250), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(N411), .D(N249), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(N411), .D(N248), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(N411), .D(N247), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(N412), .D(N410), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(N412), .D(N409), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(N412), .D(N408), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(N412), .D(N407), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(N412), .D(N406), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(N412), .D(N405), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(N412), .D(N404), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(N412), .D(N403), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(N412), .D(N402), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(N412), .D(N401), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(N412), .D(N400), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(N412), .D(N399), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(N412), .D(N398), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(N412), .D(N397), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(N412), .D(N396), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(N412), .D(N395), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(N412), .D(N394), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(N412), .D(N393), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(N412), .D(N392), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(N412), .D(N391), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(N412), .D(N390), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(N412), .D(N389), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(N412), .D(N388), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(N412), .D(N387), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(N412), .D(N386), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(N412), .D(N385), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(N412), .D(N384), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(N412), .D(N383), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(N412), .D(N382), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(N412), .D(N381), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(N412), .D(N380), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(N412), .D(N379), .Q(OUT2[0]) );
  INV_X1 U23 ( .A(n88), .ZN(n87) );
  INV_X1 U42 ( .A(n90), .ZN(n89) );
  AND2_X1 U55 ( .A1(RD1), .A2(EN), .ZN(N411) );
  AND2_X1 U56 ( .A1(EN), .A2(RD2), .ZN(N412) );
  INV_X1 U57 ( .A(DATAIN[11]), .ZN(n114) );
  BUF_X1 U58 ( .A(n842), .Z(n2) );
  BUF_X1 U59 ( .A(n883), .Z(n31) );
  BUF_X1 U60 ( .A(n867), .Z(n19) );
  BUF_X1 U61 ( .A(n865), .Z(n17) );
  BUF_X1 U62 ( .A(n857), .Z(n13) );
  BUF_X1 U63 ( .A(n847), .Z(n7) );
  INV_X1 U64 ( .A(DATAIN[25]), .ZN(n86) );
  BUF_X1 U65 ( .A(n877), .Z(n25) );
  BUF_X1 U66 ( .A(n858), .Z(n14) );
  BUF_X1 U67 ( .A(n854), .Z(n10) );
  BUF_X1 U68 ( .A(n846), .Z(n6) );
  BUF_X1 U69 ( .A(n871), .Z(n23) );
  BUF_X1 U70 ( .A(n844), .Z(n4) );
  BUF_X1 U71 ( .A(n878), .Z(n26) );
  BUF_X1 U72 ( .A(n845), .Z(n5) );
  BUF_X1 U73 ( .A(n843), .Z(n3) );
  BUF_X1 U74 ( .A(n859), .Z(n15) );
  BUF_X1 U75 ( .A(n882), .Z(n30) );
  BUF_X1 U76 ( .A(n853), .Z(n9) );
  BUF_X1 U77 ( .A(n879), .Z(n27) );
  BUF_X1 U78 ( .A(n848), .Z(n8) );
  INV_X1 U79 ( .A(n36), .ZN(n34) );
  BUF_X1 U80 ( .A(n881), .Z(n29) );
  BUF_X1 U81 ( .A(n872), .Z(n24) );
  BUF_X1 U82 ( .A(n855), .Z(n11) );
  BUF_X1 U83 ( .A(n869), .Z(n21) );
  BUF_X1 U84 ( .A(n841), .Z(n1) );
  BUF_X1 U85 ( .A(n866), .Z(n18) );
  BUF_X1 U86 ( .A(n868), .Z(n20) );
  BUF_X1 U87 ( .A(n860), .Z(n16) );
  BUF_X1 U88 ( .A(n870), .Z(n22) );
  BUF_X1 U89 ( .A(n856), .Z(n12) );
  BUF_X1 U90 ( .A(n884), .Z(n32) );
  BUF_X1 U91 ( .A(n880), .Z(n28) );
  INV_X1 U93 ( .A(n35), .ZN(n33) );
  BUF_X1 U94 ( .A(n36), .Z(n35) );
  INV_X1 U95 ( .A(n894), .ZN(n36) );
  NOR3_X1 U96 ( .A1(n171), .A2(n170), .A3(n169), .ZN(n894) );
  INV_X1 U97 ( .A(DATAIN[27]), .ZN(n82) );
  BUF_X1 U98 ( .A(n1603), .Z(n57) );
  BUF_X1 U99 ( .A(n1617), .Z(n67) );
  INV_X1 U100 ( .A(n72), .ZN(n70) );
  BUF_X1 U101 ( .A(n1581), .Z(n43) );
  BUF_X1 U102 ( .A(n1613), .Z(n63) );
  BUF_X1 U103 ( .A(n1604), .Z(n58) );
  BUF_X1 U104 ( .A(n1605), .Z(n59) );
  BUF_X1 U105 ( .A(n1606), .Z(n60) );
  BUF_X1 U106 ( .A(n1616), .Z(n66) );
  BUF_X1 U107 ( .A(n1578), .Z(n40) );
  BUF_X1 U108 ( .A(n1580), .Z(n42) );
  BUF_X1 U109 ( .A(n1593), .Z(n51) );
  BUF_X1 U110 ( .A(n1611), .Z(n61) );
  BUF_X1 U111 ( .A(n1587), .Z(n45) );
  BUF_X1 U112 ( .A(n1590), .Z(n48) );
  BUF_X1 U113 ( .A(n1576), .Z(n38) );
  BUF_X1 U114 ( .A(n1601), .Z(n55) );
  BUF_X1 U115 ( .A(n1591), .Z(n49) );
  BUF_X1 U116 ( .A(n1612), .Z(n62) );
  BUF_X1 U117 ( .A(n1589), .Z(n47) );
  BUF_X1 U118 ( .A(n1614), .Z(n64) );
  BUF_X1 U119 ( .A(n1602), .Z(n56) );
  BUF_X1 U120 ( .A(n1600), .Z(n54) );
  BUF_X1 U121 ( .A(n1599), .Z(n53) );
  BUF_X1 U122 ( .A(n1615), .Z(n65) );
  BUF_X1 U123 ( .A(n1618), .Z(n68) );
  BUF_X1 U124 ( .A(n1592), .Z(n50) );
  BUF_X1 U125 ( .A(n1594), .Z(n52) );
  BUF_X1 U126 ( .A(n1577), .Z(n39) );
  BUF_X1 U127 ( .A(n1579), .Z(n41) );
  BUF_X1 U128 ( .A(n1588), .Z(n46) );
  BUF_X1 U129 ( .A(n1575), .Z(n37) );
  BUF_X1 U130 ( .A(n1582), .Z(n44) );
  INV_X1 U131 ( .A(n71), .ZN(n69) );
  BUF_X1 U132 ( .A(n72), .Z(n71) );
  INV_X1 U133 ( .A(n1628), .ZN(n72) );
  NOR3_X1 U134 ( .A1(n904), .A2(n903), .A3(n902), .ZN(n1628) );
  INV_X1 U135 ( .A(ADD_WR[0]), .ZN(n900) );
  INV_X1 U136 ( .A(ADD_WR[2]), .ZN(n901) );
  INV_X1 U137 ( .A(ADD_WR[1]), .ZN(n897) );
  INV_X1 U138 ( .A(ADD_WR[3]), .ZN(n898) );
  INV_X1 U139 ( .A(ADD_WR[4]), .ZN(n895) );
  INV_X1 U140 ( .A(ADD_RD2[4]), .ZN(n913) );
  INV_X1 U141 ( .A(DATAIN[1]), .ZN(n134) );
  INV_X1 U145 ( .A(DATAIN[5]), .ZN(n126) );
  INV_X1 U146 ( .A(DATAIN[6]), .ZN(n124) );
  INV_X1 U147 ( .A(DATAIN[7]), .ZN(n122) );
  INV_X1 U152 ( .A(DATAIN[13]), .ZN(n110) );
  INV_X1 U153 ( .A(DATAIN[14]), .ZN(n108) );
  INV_X1 U157 ( .A(DATAIN[18]), .ZN(n100) );
  INV_X1 U159 ( .A(DATAIN[20]), .ZN(n96) );
  INV_X1 U162 ( .A(DATAIN[26]), .ZN(n84) );
  INV_X1 U167 ( .A(DATAIN[23]), .ZN(n90) );
  INV_X1 U168 ( .A(DATAIN[24]), .ZN(n88) );
  NAND4_X1 U169 ( .A1(ADD_WR[3]), .A2(WR), .A3(ADD_WR[4]), .A4(EN), .ZN(n1630)
         );
  NAND3_X1 U170 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n900), .ZN(n159) );
  OAI21_X1 U171 ( .B1(n1630), .B2(n159), .A(RST), .ZN(N114) );
  NAND3_X1 U172 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n897), .ZN(n160) );
  OAI21_X1 U173 ( .B1(n1630), .B2(n160), .A(RST), .ZN(N115) );
  NAND3_X1 U174 ( .A1(ADD_WR[2]), .A2(n900), .A3(n897), .ZN(n161) );
  OAI21_X1 U175 ( .B1(n1630), .B2(n161), .A(RST), .ZN(N116) );
  NAND3_X1 U176 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(n901), .ZN(n162) );
  OAI21_X1 U177 ( .B1(n1630), .B2(n162), .A(RST), .ZN(N117) );
  NAND3_X1 U178 ( .A1(ADD_WR[1]), .A2(n900), .A3(n901), .ZN(n163) );
  OAI21_X1 U179 ( .B1(n1630), .B2(n163), .A(RST), .ZN(N118) );
  NAND3_X1 U180 ( .A1(ADD_WR[0]), .A2(n897), .A3(n901), .ZN(n164) );
  OAI21_X1 U181 ( .B1(n1630), .B2(n164), .A(RST), .ZN(N119) );
  NAND3_X1 U182 ( .A1(n900), .A2(n897), .A3(n901), .ZN(n166) );
  OAI21_X1 U183 ( .B1(n1630), .B2(n166), .A(RST), .ZN(N120) );
  NAND3_X1 U184 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(ADD_WR[2]), .ZN(n1629)
         );
  NAND4_X1 U185 ( .A1(WR), .A2(ADD_WR[4]), .A3(EN), .A4(n898), .ZN(n157) );
  OAI21_X1 U186 ( .B1(n1629), .B2(n157), .A(RST), .ZN(N121) );
  OAI21_X1 U187 ( .B1(n159), .B2(n157), .A(RST), .ZN(N122) );
  OAI21_X1 U188 ( .B1(n160), .B2(n157), .A(RST), .ZN(N123) );
  OAI21_X1 U189 ( .B1(n161), .B2(n157), .A(RST), .ZN(N124) );
  OAI21_X1 U190 ( .B1(n162), .B2(n157), .A(n151), .ZN(N125) );
  OAI21_X1 U191 ( .B1(n163), .B2(n157), .A(n144), .ZN(N126) );
  OAI21_X1 U192 ( .B1(n164), .B2(n157), .A(n154), .ZN(N127) );
  OAI21_X1 U193 ( .B1(n166), .B2(n157), .A(n141), .ZN(N128) );
  NAND4_X1 U194 ( .A1(WR), .A2(ADD_WR[3]), .A3(EN), .A4(n895), .ZN(n158) );
  OAI21_X1 U195 ( .B1(n1629), .B2(n158), .A(n139), .ZN(N129) );
  OAI21_X1 U196 ( .B1(n159), .B2(n158), .A(n138), .ZN(N130) );
  OAI21_X1 U197 ( .B1(n160), .B2(n158), .A(n137), .ZN(N131) );
  OAI21_X1 U198 ( .B1(n161), .B2(n158), .A(RST), .ZN(N132) );
  OAI21_X1 U199 ( .B1(n162), .B2(n158), .A(n140), .ZN(N133) );
  OAI21_X1 U200 ( .B1(n163), .B2(n158), .A(n147), .ZN(N134) );
  OAI21_X1 U201 ( .B1(n164), .B2(n158), .A(n142), .ZN(N135) );
  OAI21_X1 U202 ( .B1(n166), .B2(n158), .A(RST), .ZN(N136) );
  NAND4_X1 U203 ( .A1(WR), .A2(EN), .A3(n898), .A4(n895), .ZN(n165) );
  OAI21_X1 U204 ( .B1(n1629), .B2(n165), .A(RST), .ZN(N137) );
  OAI21_X1 U205 ( .B1(n159), .B2(n165), .A(n151), .ZN(N138) );
  OAI21_X1 U206 ( .B1(n160), .B2(n165), .A(n155), .ZN(N139) );
  OAI21_X1 U207 ( .B1(n161), .B2(n165), .A(RST), .ZN(N140) );
  OAI21_X1 U208 ( .B1(n162), .B2(n165), .A(RST), .ZN(N141) );
  OAI21_X1 U209 ( .B1(n163), .B2(n165), .A(RST), .ZN(N142) );
  OAI21_X1 U210 ( .B1(n164), .B2(n165), .A(RST), .ZN(N143) );
  OAI21_X1 U211 ( .B1(n166), .B2(n165), .A(n148), .ZN(N144) );
  INV_X1 U212 ( .A(ADD_RD1[1]), .ZN(n173) );
  OAI221_X1 U213 ( .B1(ADD_WR[1]), .B2(n173), .C1(n897), .C2(ADD_RD1[1]), .A(
        WR), .ZN(n171) );
  AOI22_X1 U214 ( .A1(n901), .A2(ADD_RD1[2]), .B1(ADD_RD1[4]), .B2(n895), .ZN(
        n167) );
  OAI221_X1 U215 ( .B1(n901), .B2(ADD_RD1[2]), .C1(n895), .C2(ADD_RD1[4]), .A(
        n167), .ZN(n170) );
  AOI22_X1 U216 ( .A1(n898), .A2(ADD_RD1[3]), .B1(ADD_RD1[0]), .B2(n900), .ZN(
        n168) );
  OAI221_X1 U217 ( .B1(n898), .B2(ADD_RD1[3]), .C1(n900), .C2(ADD_RD1[0]), .A(
        n168), .ZN(n169) );
  NAND2_X1 U218 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n201) );
  INV_X1 U219 ( .A(ADD_RD1[3]), .ZN(n174) );
  INV_X1 U220 ( .A(ADD_RD1[4]), .ZN(n179) );
  NAND3_X1 U221 ( .A1(ADD_RD1[0]), .A2(n174), .A3(n179), .ZN(n194) );
  NOR2_X1 U222 ( .A1(n201), .A2(n194), .ZN(n878) );
  INV_X1 U223 ( .A(ADD_RD1[0]), .ZN(n180) );
  NAND3_X1 U224 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n180), .ZN(n186) );
  NOR2_X1 U225 ( .A1(n201), .A2(n186), .ZN(n880) );
  AOI22_X1 U226 ( .A1(\REGISTERS[7][0] ), .A2(n878), .B1(\REGISTERS[30][0] ), 
        .B2(n28), .ZN(n178) );
  INV_X1 U227 ( .A(ADD_RD1[2]), .ZN(n172) );
  NAND2_X1 U228 ( .A1(ADD_RD1[1]), .A2(n172), .ZN(n196) );
  NOR2_X1 U229 ( .A1(n186), .A2(n196), .ZN(n879) );
  NAND3_X1 U230 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n179), .ZN(n199) );
  NAND2_X1 U231 ( .A1(ADD_RD1[2]), .A2(n173), .ZN(n193) );
  NOR2_X1 U232 ( .A1(n199), .A2(n193), .ZN(n884) );
  AOI22_X1 U233 ( .A1(\REGISTERS[26][0] ), .A2(n879), .B1(\REGISTERS[13][0] ), 
        .B2(n32), .ZN(n177) );
  NAND2_X1 U234 ( .A1(n173), .A2(n172), .ZN(n198) );
  NAND3_X1 U235 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[0]), .A3(ADD_RD1[4]), .ZN(n200)
         );
  NOR2_X1 U236 ( .A1(n198), .A2(n200), .ZN(n882) );
  NOR2_X1 U237 ( .A1(n186), .A2(n193), .ZN(n856) );
  AOI22_X1 U238 ( .A1(\REGISTERS[25][0] ), .A2(n882), .B1(\REGISTERS[28][0] ), 
        .B2(n12), .ZN(n176) );
  NAND3_X1 U239 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n174), .ZN(n187) );
  NOR2_X1 U240 ( .A1(n198), .A2(n187), .ZN(n854) );
  NOR2_X1 U241 ( .A1(n193), .A2(n187), .ZN(n870) );
  AOI22_X1 U242 ( .A1(\REGISTERS[17][0] ), .A2(n854), .B1(\REGISTERS[21][0] ), 
        .B2(n22), .ZN(n175) );
  NAND4_X1 U243 ( .A1(n178), .A2(n177), .A3(n176), .A4(n175), .ZN(n209) );
  NOR2_X1 U244 ( .A1(n193), .A2(n200), .ZN(n858) );
  NOR2_X1 U245 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[0]), .ZN(n185) );
  NAND2_X1 U246 ( .A1(n185), .A2(n179), .ZN(n195) );
  NOR2_X1 U247 ( .A1(n201), .A2(n195), .ZN(n860) );
  AOI22_X1 U248 ( .A1(\REGISTERS[29][0] ), .A2(n858), .B1(\REGISTERS[6][0] ), 
        .B2(n16), .ZN(n184) );
  NAND3_X1 U249 ( .A1(ADD_RD1[3]), .A2(n180), .A3(n179), .ZN(n192) );
  NOR2_X1 U250 ( .A1(n196), .A2(n192), .ZN(n883) );
  NOR2_X1 U251 ( .A1(n198), .A2(n192), .ZN(n868) );
  AOI22_X1 U252 ( .A1(\REGISTERS[10][0] ), .A2(n883), .B1(\REGISTERS[8][0] ), 
        .B2(n20), .ZN(n183) );
  NOR2_X1 U253 ( .A1(n201), .A2(n199), .ZN(n877) );
  NOR2_X1 U254 ( .A1(n201), .A2(n192), .ZN(n866) );
  AOI22_X1 U255 ( .A1(\REGISTERS[15][0] ), .A2(n877), .B1(\REGISTERS[14][0] ), 
        .B2(n18), .ZN(n182) );
  NOR2_X1 U256 ( .A1(n201), .A2(n187), .ZN(n842) );
  NOR2_X1 U257 ( .A1(n198), .A2(n195), .ZN(n841) );
  AOI22_X1 U258 ( .A1(\REGISTERS[23][0] ), .A2(n842), .B1(\REGISTERS[0][0] ), 
        .B2(n1), .ZN(n181) );
  NAND4_X1 U259 ( .A1(n184), .A2(n183), .A3(n182), .A4(n181), .ZN(n208) );
  NOR2_X1 U260 ( .A1(n194), .A2(n198), .ZN(n848) );
  NAND2_X1 U261 ( .A1(ADD_RD1[4]), .A2(n185), .ZN(n197) );
  NOR2_X1 U262 ( .A1(n196), .A2(n197), .ZN(n869) );
  AOI22_X1 U263 ( .A1(\REGISTERS[1][0] ), .A2(n848), .B1(\REGISTERS[18][0] ), 
        .B2(n21), .ZN(n191) );
  NOR2_X1 U264 ( .A1(n196), .A2(n200), .ZN(n844) );
  NOR2_X1 U265 ( .A1(n193), .A2(n197), .ZN(n865) );
  AOI22_X1 U266 ( .A1(\REGISTERS[27][0] ), .A2(n844), .B1(\REGISTERS[20][0] ), 
        .B2(n865), .ZN(n190) );
  NOR2_X1 U267 ( .A1(n186), .A2(n198), .ZN(n846) );
  NOR2_X1 U268 ( .A1(n194), .A2(n196), .ZN(n855) );
  AOI22_X1 U269 ( .A1(\REGISTERS[24][0] ), .A2(n846), .B1(\REGISTERS[3][0] ), 
        .B2(n11), .ZN(n189) );
  NOR2_X1 U270 ( .A1(n196), .A2(n187), .ZN(n847) );
  NOR2_X1 U271 ( .A1(n193), .A2(n195), .ZN(n867) );
  AOI22_X1 U272 ( .A1(\REGISTERS[19][0] ), .A2(n847), .B1(\REGISTERS[4][0] ), 
        .B2(n867), .ZN(n188) );
  NAND4_X1 U273 ( .A1(n191), .A2(n190), .A3(n189), .A4(n188), .ZN(n207) );
  NOR2_X1 U274 ( .A1(n193), .A2(n192), .ZN(n857) );
  NOR2_X1 U275 ( .A1(n194), .A2(n193), .ZN(n872) );
  AOI22_X1 U276 ( .A1(\REGISTERS[12][0] ), .A2(n857), .B1(\REGISTERS[5][0] ), 
        .B2(n24), .ZN(n205) );
  NOR2_X1 U277 ( .A1(n196), .A2(n195), .ZN(n843) );
  NOR2_X1 U278 ( .A1(n196), .A2(n199), .ZN(n881) );
  AOI22_X1 U279 ( .A1(\REGISTERS[2][0] ), .A2(n843), .B1(\REGISTERS[11][0] ), 
        .B2(n29), .ZN(n204) );
  NOR2_X1 U280 ( .A1(n201), .A2(n197), .ZN(n859) );
  NOR2_X1 U281 ( .A1(n198), .A2(n197), .ZN(n871) );
  AOI22_X1 U282 ( .A1(\REGISTERS[22][0] ), .A2(n859), .B1(\REGISTERS[16][0] ), 
        .B2(n871), .ZN(n203) );
  NOR2_X1 U283 ( .A1(n199), .A2(n198), .ZN(n853) );
  NOR2_X1 U284 ( .A1(n201), .A2(n200), .ZN(n845) );
  AOI22_X1 U285 ( .A1(\REGISTERS[9][0] ), .A2(n853), .B1(\REGISTERS[31][0] ), 
        .B2(n845), .ZN(n202) );
  NAND4_X1 U286 ( .A1(n205), .A2(n204), .A3(n203), .A4(n202), .ZN(n206) );
  NOR4_X1 U287 ( .A1(n209), .A2(n208), .A3(n207), .A4(n206), .ZN(n210) );
  AOI22_X1 U288 ( .A1(n33), .A2(n2677), .B1(n210), .B2(n36), .ZN(N247) );
  AOI22_X1 U289 ( .A1(n842), .A2(\REGISTERS[23][1] ), .B1(n8), .B2(
        \REGISTERS[1][1] ), .ZN(n214) );
  AOI22_X1 U290 ( .A1(n27), .A2(\REGISTERS[26][1] ), .B1(n21), .B2(
        \REGISTERS[18][1] ), .ZN(n213) );
  AOI22_X1 U291 ( .A1(n855), .A2(\REGISTERS[3][1] ), .B1(n857), .B2(
        \REGISTERS[12][1] ), .ZN(n212) );
  AOI22_X1 U292 ( .A1(n868), .A2(\REGISTERS[8][1] ), .B1(n872), .B2(
        \REGISTERS[5][1] ), .ZN(n211) );
  NAND4_X1 U293 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(n230) );
  AOI22_X1 U294 ( .A1(n883), .A2(\REGISTERS[10][1] ), .B1(n18), .B2(
        \REGISTERS[14][1] ), .ZN(n218) );
  AOI22_X1 U295 ( .A1(n12), .A2(\REGISTERS[28][1] ), .B1(n847), .B2(
        \REGISTERS[19][1] ), .ZN(n217) );
  AOI22_X1 U296 ( .A1(n860), .A2(\REGISTERS[6][1] ), .B1(n865), .B2(
        \REGISTERS[20][1] ), .ZN(n216) );
  AOI22_X1 U297 ( .A1(n867), .A2(\REGISTERS[4][1] ), .B1(n9), .B2(
        \REGISTERS[9][1] ), .ZN(n215) );
  NAND4_X1 U298 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(n229) );
  AOI22_X1 U299 ( .A1(n30), .A2(\REGISTERS[25][1] ), .B1(n15), .B2(
        \REGISTERS[22][1] ), .ZN(n222) );
  AOI22_X1 U300 ( .A1(n870), .A2(\REGISTERS[21][1] ), .B1(n881), .B2(
        \REGISTERS[11][1] ), .ZN(n221) );
  AOI22_X1 U301 ( .A1(n3), .A2(\REGISTERS[2][1] ), .B1(n5), .B2(
        \REGISTERS[31][1] ), .ZN(n220) );
  AOI22_X1 U302 ( .A1(n26), .A2(\REGISTERS[7][1] ), .B1(n4), .B2(
        \REGISTERS[27][1] ), .ZN(n219) );
  NAND4_X1 U303 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(n228) );
  AOI22_X1 U304 ( .A1(n841), .A2(\REGISTERS[0][1] ), .B1(n23), .B2(
        \REGISTERS[16][1] ), .ZN(n226) );
  AOI22_X1 U305 ( .A1(n32), .A2(\REGISTERS[13][1] ), .B1(n6), .B2(
        \REGISTERS[24][1] ), .ZN(n225) );
  AOI22_X1 U306 ( .A1(n28), .A2(\REGISTERS[30][1] ), .B1(n10), .B2(
        \REGISTERS[17][1] ), .ZN(n224) );
  AOI22_X1 U307 ( .A1(n14), .A2(\REGISTERS[29][1] ), .B1(n25), .B2(
        \REGISTERS[15][1] ), .ZN(n223) );
  NAND4_X1 U308 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(n227) );
  NOR4_X1 U309 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(n231) );
  AOI22_X1 U310 ( .A1(n34), .A2(n134), .B1(n231), .B2(n35), .ZN(N248) );
  AOI22_X1 U311 ( .A1(n7), .A2(\REGISTERS[19][2] ), .B1(n13), .B2(
        \REGISTERS[12][2] ), .ZN(n235) );
  AOI22_X1 U312 ( .A1(n10), .A2(\REGISTERS[17][2] ), .B1(n853), .B2(
        \REGISTERS[9][2] ), .ZN(n234) );
  AOI22_X1 U313 ( .A1(n12), .A2(\REGISTERS[28][2] ), .B1(n15), .B2(
        \REGISTERS[22][2] ), .ZN(n233) );
  AOI22_X1 U314 ( .A1(n16), .A2(\REGISTERS[6][2] ), .B1(n23), .B2(
        \REGISTERS[16][2] ), .ZN(n232) );
  NAND4_X1 U315 ( .A1(n235), .A2(n234), .A3(n233), .A4(n232), .ZN(n251) );
  AOI22_X1 U316 ( .A1(n30), .A2(\REGISTERS[25][2] ), .B1(n24), .B2(
        \REGISTERS[5][2] ), .ZN(n239) );
  AOI22_X1 U317 ( .A1(n22), .A2(\REGISTERS[21][2] ), .B1(n21), .B2(
        \REGISTERS[18][2] ), .ZN(n238) );
  AOI22_X1 U318 ( .A1(n848), .A2(\REGISTERS[1][2] ), .B1(n17), .B2(
        \REGISTERS[20][2] ), .ZN(n237) );
  AOI22_X1 U319 ( .A1(n20), .A2(\REGISTERS[8][2] ), .B1(n18), .B2(
        \REGISTERS[14][2] ), .ZN(n236) );
  NAND4_X1 U320 ( .A1(n239), .A2(n238), .A3(n237), .A4(n236), .ZN(n250) );
  AOI22_X1 U321 ( .A1(n27), .A2(\REGISTERS[26][2] ), .B1(n6), .B2(
        \REGISTERS[24][2] ), .ZN(n243) );
  AOI22_X1 U322 ( .A1(n878), .A2(\REGISTERS[7][2] ), .B1(n19), .B2(
        \REGISTERS[4][2] ), .ZN(n242) );
  AOI22_X1 U323 ( .A1(n1), .A2(\REGISTERS[0][2] ), .B1(n4), .B2(
        \REGISTERS[27][2] ), .ZN(n241) );
  AOI22_X1 U324 ( .A1(n843), .A2(\REGISTERS[2][2] ), .B1(n29), .B2(
        \REGISTERS[11][2] ), .ZN(n240) );
  NAND4_X1 U325 ( .A1(n243), .A2(n242), .A3(n241), .A4(n240), .ZN(n249) );
  AOI22_X1 U326 ( .A1(n31), .A2(\REGISTERS[10][2] ), .B1(n2), .B2(
        \REGISTERS[23][2] ), .ZN(n247) );
  AOI22_X1 U327 ( .A1(n28), .A2(\REGISTERS[30][2] ), .B1(n845), .B2(
        \REGISTERS[31][2] ), .ZN(n246) );
  AOI22_X1 U328 ( .A1(n877), .A2(\REGISTERS[15][2] ), .B1(n855), .B2(
        \REGISTERS[3][2] ), .ZN(n245) );
  AOI22_X1 U329 ( .A1(n32), .A2(\REGISTERS[13][2] ), .B1(n14), .B2(
        \REGISTERS[29][2] ), .ZN(n244) );
  NAND4_X1 U330 ( .A1(n247), .A2(n246), .A3(n245), .A4(n244), .ZN(n248) );
  NOR4_X1 U331 ( .A1(n251), .A2(n250), .A3(n249), .A4(n248), .ZN(n252) );
  AOI22_X1 U332 ( .A1(n34), .A2(n2669), .B1(n252), .B2(n36), .ZN(N249) );
  AOI22_X1 U333 ( .A1(n841), .A2(\REGISTERS[0][3] ), .B1(n9), .B2(
        \REGISTERS[9][3] ), .ZN(n256) );
  AOI22_X1 U334 ( .A1(n28), .A2(\REGISTERS[30][3] ), .B1(n22), .B2(
        \REGISTERS[21][3] ), .ZN(n255) );
  AOI22_X1 U335 ( .A1(n16), .A2(\REGISTERS[6][3] ), .B1(n29), .B2(
        \REGISTERS[11][3] ), .ZN(n254) );
  AOI22_X1 U336 ( .A1(n19), .A2(\REGISTERS[4][3] ), .B1(n23), .B2(
        \REGISTERS[16][3] ), .ZN(n253) );
  NAND4_X1 U337 ( .A1(n256), .A2(n255), .A3(n254), .A4(n253), .ZN(n272) );
  AOI22_X1 U338 ( .A1(n21), .A2(\REGISTERS[18][3] ), .B1(n11), .B2(
        \REGISTERS[3][3] ), .ZN(n260) );
  AOI22_X1 U339 ( .A1(n26), .A2(\REGISTERS[7][3] ), .B1(n4), .B2(
        \REGISTERS[27][3] ), .ZN(n259) );
  AOI22_X1 U340 ( .A1(n854), .A2(\REGISTERS[17][3] ), .B1(n5), .B2(
        \REGISTERS[31][3] ), .ZN(n258) );
  AOI22_X1 U341 ( .A1(n30), .A2(\REGISTERS[25][3] ), .B1(n12), .B2(
        \REGISTERS[28][3] ), .ZN(n257) );
  NAND4_X1 U342 ( .A1(n260), .A2(n259), .A3(n258), .A4(n257), .ZN(n271) );
  AOI22_X1 U343 ( .A1(n868), .A2(\REGISTERS[8][3] ), .B1(n25), .B2(
        \REGISTERS[15][3] ), .ZN(n264) );
  AOI22_X1 U344 ( .A1(n872), .A2(\REGISTERS[5][3] ), .B1(n3), .B2(
        \REGISTERS[2][3] ), .ZN(n263) );
  AOI22_X1 U345 ( .A1(n883), .A2(\REGISTERS[10][3] ), .B1(n17), .B2(
        \REGISTERS[20][3] ), .ZN(n262) );
  AOI22_X1 U346 ( .A1(n866), .A2(\REGISTERS[14][3] ), .B1(n8), .B2(
        \REGISTERS[1][3] ), .ZN(n261) );
  NAND4_X1 U347 ( .A1(n264), .A2(n263), .A3(n262), .A4(n261), .ZN(n270) );
  AOI22_X1 U348 ( .A1(n14), .A2(\REGISTERS[29][3] ), .B1(n13), .B2(
        \REGISTERS[12][3] ), .ZN(n268) );
  AOI22_X1 U349 ( .A1(n884), .A2(\REGISTERS[13][3] ), .B1(n15), .B2(
        \REGISTERS[22][3] ), .ZN(n267) );
  AOI22_X1 U350 ( .A1(n842), .A2(\REGISTERS[23][3] ), .B1(n6), .B2(
        \REGISTERS[24][3] ), .ZN(n266) );
  AOI22_X1 U351 ( .A1(n27), .A2(\REGISTERS[26][3] ), .B1(n7), .B2(
        \REGISTERS[19][3] ), .ZN(n265) );
  NAND4_X1 U352 ( .A1(n268), .A2(n267), .A3(n266), .A4(n265), .ZN(n269) );
  NOR4_X1 U353 ( .A1(n272), .A2(n271), .A3(n270), .A4(n269), .ZN(n273) );
  AOI22_X1 U354 ( .A1(n34), .A2(n2670), .B1(n273), .B2(n35), .ZN(N250) );
  AOI22_X1 U355 ( .A1(n27), .A2(\REGISTERS[26][4] ), .B1(n19), .B2(
        \REGISTERS[4][4] ), .ZN(n277) );
  AOI22_X1 U356 ( .A1(n869), .A2(\REGISTERS[18][4] ), .B1(n11), .B2(
        \REGISTERS[3][4] ), .ZN(n276) );
  AOI22_X1 U357 ( .A1(n856), .A2(\REGISTERS[28][4] ), .B1(n22), .B2(
        \REGISTERS[21][4] ), .ZN(n275) );
  AOI22_X1 U358 ( .A1(n18), .A2(\REGISTERS[14][4] ), .B1(n853), .B2(
        \REGISTERS[9][4] ), .ZN(n274) );
  NAND4_X1 U359 ( .A1(n277), .A2(n276), .A3(n275), .A4(n274), .ZN(n293) );
  AOI22_X1 U360 ( .A1(n25), .A2(\REGISTERS[15][4] ), .B1(n29), .B2(
        \REGISTERS[11][4] ), .ZN(n281) );
  AOI22_X1 U361 ( .A1(n878), .A2(\REGISTERS[7][4] ), .B1(n1), .B2(
        \REGISTERS[0][4] ), .ZN(n280) );
  AOI22_X1 U362 ( .A1(n865), .A2(\REGISTERS[20][4] ), .B1(n13), .B2(
        \REGISTERS[12][4] ), .ZN(n279) );
  AOI22_X1 U363 ( .A1(n14), .A2(\REGISTERS[29][4] ), .B1(n23), .B2(
        \REGISTERS[16][4] ), .ZN(n278) );
  NAND4_X1 U364 ( .A1(n281), .A2(n280), .A3(n279), .A4(n278), .ZN(n292) );
  AOI22_X1 U365 ( .A1(n2), .A2(\REGISTERS[23][4] ), .B1(n24), .B2(
        \REGISTERS[5][4] ), .ZN(n285) );
  AOI22_X1 U366 ( .A1(n4), .A2(\REGISTERS[27][4] ), .B1(n6), .B2(
        \REGISTERS[24][4] ), .ZN(n284) );
  AOI22_X1 U367 ( .A1(n10), .A2(\REGISTERS[17][4] ), .B1(n7), .B2(
        \REGISTERS[19][4] ), .ZN(n283) );
  AOI22_X1 U368 ( .A1(n32), .A2(\REGISTERS[13][4] ), .B1(n30), .B2(
        \REGISTERS[25][4] ), .ZN(n282) );
  NAND4_X1 U369 ( .A1(n285), .A2(n284), .A3(n283), .A4(n282), .ZN(n291) );
  AOI22_X1 U370 ( .A1(n28), .A2(\REGISTERS[30][4] ), .B1(n15), .B2(
        \REGISTERS[22][4] ), .ZN(n289) );
  AOI22_X1 U371 ( .A1(n20), .A2(\REGISTERS[8][4] ), .B1(n8), .B2(
        \REGISTERS[1][4] ), .ZN(n288) );
  AOI22_X1 U372 ( .A1(n31), .A2(\REGISTERS[10][4] ), .B1(n845), .B2(
        \REGISTERS[31][4] ), .ZN(n287) );
  AOI22_X1 U373 ( .A1(n860), .A2(\REGISTERS[6][4] ), .B1(n3), .B2(
        \REGISTERS[2][4] ), .ZN(n286) );
  NAND4_X1 U374 ( .A1(n289), .A2(n288), .A3(n287), .A4(n286), .ZN(n290) );
  NOR4_X1 U375 ( .A1(n293), .A2(n292), .A3(n291), .A4(n290), .ZN(n294) );
  AOI22_X1 U376 ( .A1(n34), .A2(n2676), .B1(n294), .B2(n36), .ZN(N251) );
  AOI22_X1 U377 ( .A1(n14), .A2(\REGISTERS[29][5] ), .B1(n11), .B2(
        \REGISTERS[3][5] ), .ZN(n298) );
  AOI22_X1 U378 ( .A1(n1), .A2(\REGISTERS[0][5] ), .B1(n17), .B2(
        \REGISTERS[20][5] ), .ZN(n297) );
  AOI22_X1 U379 ( .A1(n846), .A2(\REGISTERS[24][5] ), .B1(n9), .B2(
        \REGISTERS[9][5] ), .ZN(n296) );
  AOI22_X1 U380 ( .A1(n879), .A2(\REGISTERS[26][5] ), .B1(n2), .B2(
        \REGISTERS[23][5] ), .ZN(n295) );
  NAND4_X1 U381 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(n314) );
  AOI22_X1 U382 ( .A1(n30), .A2(\REGISTERS[25][5] ), .B1(n12), .B2(
        \REGISTERS[28][5] ), .ZN(n302) );
  AOI22_X1 U383 ( .A1(n28), .A2(\REGISTERS[30][5] ), .B1(n10), .B2(
        \REGISTERS[17][5] ), .ZN(n301) );
  AOI22_X1 U384 ( .A1(n881), .A2(\REGISTERS[11][5] ), .B1(n23), .B2(
        \REGISTERS[16][5] ), .ZN(n300) );
  AOI22_X1 U385 ( .A1(n22), .A2(\REGISTERS[21][5] ), .B1(n31), .B2(
        \REGISTERS[10][5] ), .ZN(n299) );
  NAND4_X1 U386 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(n313) );
  AOI22_X1 U387 ( .A1(n844), .A2(\REGISTERS[27][5] ), .B1(n24), .B2(
        \REGISTERS[5][5] ), .ZN(n306) );
  AOI22_X1 U388 ( .A1(n16), .A2(\REGISTERS[6][5] ), .B1(n8), .B2(
        \REGISTERS[1][5] ), .ZN(n305) );
  AOI22_X1 U389 ( .A1(n32), .A2(\REGISTERS[13][5] ), .B1(n25), .B2(
        \REGISTERS[15][5] ), .ZN(n304) );
  AOI22_X1 U390 ( .A1(n26), .A2(\REGISTERS[7][5] ), .B1(n15), .B2(
        \REGISTERS[22][5] ), .ZN(n303) );
  NAND4_X1 U391 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(n312) );
  AOI22_X1 U392 ( .A1(n20), .A2(\REGISTERS[8][5] ), .B1(n5), .B2(
        \REGISTERS[31][5] ), .ZN(n310) );
  AOI22_X1 U393 ( .A1(n866), .A2(\REGISTERS[14][5] ), .B1(n3), .B2(
        \REGISTERS[2][5] ), .ZN(n309) );
  AOI22_X1 U394 ( .A1(n869), .A2(\REGISTERS[18][5] ), .B1(n7), .B2(
        \REGISTERS[19][5] ), .ZN(n308) );
  AOI22_X1 U395 ( .A1(n867), .A2(\REGISTERS[4][5] ), .B1(n13), .B2(
        \REGISTERS[12][5] ), .ZN(n307) );
  NAND4_X1 U396 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(n311) );
  NOR4_X1 U397 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(n315) );
  AOI22_X1 U398 ( .A1(n34), .A2(n2662), .B1(n315), .B2(n35), .ZN(N252) );
  AOI22_X1 U399 ( .A1(n841), .A2(\REGISTERS[0][6] ), .B1(n21), .B2(
        \REGISTERS[18][6] ), .ZN(n319) );
  AOI22_X1 U400 ( .A1(n22), .A2(\REGISTERS[21][6] ), .B1(n845), .B2(
        \REGISTERS[31][6] ), .ZN(n318) );
  AOI22_X1 U401 ( .A1(n881), .A2(\REGISTERS[11][6] ), .B1(n23), .B2(
        \REGISTERS[16][6] ), .ZN(n317) );
  AOI22_X1 U402 ( .A1(n30), .A2(\REGISTERS[25][6] ), .B1(n7), .B2(
        \REGISTERS[19][6] ), .ZN(n316) );
  NAND4_X1 U403 ( .A1(n319), .A2(n318), .A3(n317), .A4(n316), .ZN(n335) );
  AOI22_X1 U404 ( .A1(n878), .A2(\REGISTERS[7][6] ), .B1(n25), .B2(
        \REGISTERS[15][6] ), .ZN(n323) );
  AOI22_X1 U405 ( .A1(n854), .A2(\REGISTERS[17][6] ), .B1(n8), .B2(
        \REGISTERS[1][6] ), .ZN(n322) );
  AOI22_X1 U406 ( .A1(n11), .A2(\REGISTERS[3][6] ), .B1(n24), .B2(
        \REGISTERS[5][6] ), .ZN(n321) );
  AOI22_X1 U407 ( .A1(n856), .A2(\REGISTERS[28][6] ), .B1(n16), .B2(
        \REGISTERS[6][6] ), .ZN(n320) );
  NAND4_X1 U408 ( .A1(n323), .A2(n322), .A3(n321), .A4(n320), .ZN(n334) );
  AOI22_X1 U409 ( .A1(n18), .A2(\REGISTERS[14][6] ), .B1(n2), .B2(
        \REGISTERS[23][6] ), .ZN(n327) );
  AOI22_X1 U410 ( .A1(n32), .A2(\REGISTERS[13][6] ), .B1(n4), .B2(
        \REGISTERS[27][6] ), .ZN(n326) );
  AOI22_X1 U411 ( .A1(n28), .A2(\REGISTERS[30][6] ), .B1(n20), .B2(
        \REGISTERS[8][6] ), .ZN(n325) );
  AOI22_X1 U412 ( .A1(n865), .A2(\REGISTERS[20][6] ), .B1(n19), .B2(
        \REGISTERS[4][6] ), .ZN(n324) );
  NAND4_X1 U413 ( .A1(n327), .A2(n326), .A3(n325), .A4(n324), .ZN(n333) );
  AOI22_X1 U414 ( .A1(n27), .A2(\REGISTERS[26][6] ), .B1(n6), .B2(
        \REGISTERS[24][6] ), .ZN(n331) );
  AOI22_X1 U415 ( .A1(n3), .A2(\REGISTERS[2][6] ), .B1(n853), .B2(
        \REGISTERS[9][6] ), .ZN(n330) );
  AOI22_X1 U416 ( .A1(n14), .A2(\REGISTERS[29][6] ), .B1(n13), .B2(
        \REGISTERS[12][6] ), .ZN(n329) );
  AOI22_X1 U417 ( .A1(n883), .A2(\REGISTERS[10][6] ), .B1(n15), .B2(
        \REGISTERS[22][6] ), .ZN(n328) );
  NAND4_X1 U418 ( .A1(n331), .A2(n330), .A3(n329), .A4(n328), .ZN(n332) );
  NOR4_X1 U419 ( .A1(n335), .A2(n334), .A3(n333), .A4(n332), .ZN(n336) );
  AOI22_X1 U420 ( .A1(n894), .A2(n2659), .B1(n336), .B2(n35), .ZN(N253) );
  AOI22_X1 U421 ( .A1(n12), .A2(\REGISTERS[28][7] ), .B1(n853), .B2(
        \REGISTERS[9][7] ), .ZN(n340) );
  AOI22_X1 U422 ( .A1(n16), .A2(\REGISTERS[6][7] ), .B1(n2), .B2(
        \REGISTERS[23][7] ), .ZN(n339) );
  AOI22_X1 U423 ( .A1(n14), .A2(\REGISTERS[29][7] ), .B1(n23), .B2(
        \REGISTERS[16][7] ), .ZN(n338) );
  AOI22_X1 U424 ( .A1(n6), .A2(\REGISTERS[24][7] ), .B1(n7), .B2(
        \REGISTERS[19][7] ), .ZN(n337) );
  NAND4_X1 U425 ( .A1(n340), .A2(n339), .A3(n338), .A4(n337), .ZN(n356) );
  AOI22_X1 U426 ( .A1(n869), .A2(\REGISTERS[18][7] ), .B1(n24), .B2(
        \REGISTERS[5][7] ), .ZN(n344) );
  AOI22_X1 U427 ( .A1(n28), .A2(\REGISTERS[30][7] ), .B1(n3), .B2(
        \REGISTERS[2][7] ), .ZN(n343) );
  AOI22_X1 U428 ( .A1(n884), .A2(\REGISTERS[13][7] ), .B1(n17), .B2(
        \REGISTERS[20][7] ), .ZN(n342) );
  AOI22_X1 U429 ( .A1(n10), .A2(\REGISTERS[17][7] ), .B1(n13), .B2(
        \REGISTERS[12][7] ), .ZN(n341) );
  NAND4_X1 U430 ( .A1(n344), .A2(n343), .A3(n342), .A4(n341), .ZN(n355) );
  AOI22_X1 U431 ( .A1(n20), .A2(\REGISTERS[8][7] ), .B1(n4), .B2(
        \REGISTERS[27][7] ), .ZN(n348) );
  AOI22_X1 U432 ( .A1(n882), .A2(\REGISTERS[25][7] ), .B1(n22), .B2(
        \REGISTERS[21][7] ), .ZN(n347) );
  AOI22_X1 U433 ( .A1(n31), .A2(\REGISTERS[10][7] ), .B1(n8), .B2(
        \REGISTERS[1][7] ), .ZN(n346) );
  AOI22_X1 U434 ( .A1(n27), .A2(\REGISTERS[26][7] ), .B1(n1), .B2(
        \REGISTERS[0][7] ), .ZN(n345) );
  NAND4_X1 U435 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .ZN(n354) );
  AOI22_X1 U436 ( .A1(n877), .A2(\REGISTERS[15][7] ), .B1(n29), .B2(
        \REGISTERS[11][7] ), .ZN(n352) );
  AOI22_X1 U437 ( .A1(n878), .A2(\REGISTERS[7][7] ), .B1(n15), .B2(
        \REGISTERS[22][7] ), .ZN(n351) );
  AOI22_X1 U438 ( .A1(n19), .A2(\REGISTERS[4][7] ), .B1(n845), .B2(
        \REGISTERS[31][7] ), .ZN(n350) );
  AOI22_X1 U439 ( .A1(n18), .A2(\REGISTERS[14][7] ), .B1(n11), .B2(
        \REGISTERS[3][7] ), .ZN(n349) );
  NAND4_X1 U440 ( .A1(n352), .A2(n351), .A3(n350), .A4(n349), .ZN(n353) );
  NOR4_X1 U441 ( .A1(n356), .A2(n355), .A3(n354), .A4(n353), .ZN(n357) );
  AOI22_X1 U442 ( .A1(n894), .A2(n122), .B1(n357), .B2(n36), .ZN(N254) );
  AOI22_X1 U443 ( .A1(n878), .A2(\REGISTERS[7][8] ), .B1(n18), .B2(
        \REGISTERS[14][8] ), .ZN(n361) );
  AOI22_X1 U444 ( .A1(n880), .A2(\REGISTERS[30][8] ), .B1(n32), .B2(
        \REGISTERS[13][8] ), .ZN(n360) );
  AOI22_X1 U445 ( .A1(n27), .A2(\REGISTERS[26][8] ), .B1(n30), .B2(
        \REGISTERS[25][8] ), .ZN(n359) );
  AOI22_X1 U446 ( .A1(n12), .A2(\REGISTERS[28][8] ), .B1(n1), .B2(
        \REGISTERS[0][8] ), .ZN(n358) );
  NAND4_X1 U447 ( .A1(n361), .A2(n360), .A3(n359), .A4(n358), .ZN(n377) );
  AOI22_X1 U448 ( .A1(n20), .A2(\REGISTERS[8][8] ), .B1(n19), .B2(
        \REGISTERS[4][8] ), .ZN(n365) );
  AOI22_X1 U449 ( .A1(n858), .A2(\REGISTERS[29][8] ), .B1(n7), .B2(
        \REGISTERS[19][8] ), .ZN(n364) );
  AOI22_X1 U450 ( .A1(n8), .A2(\REGISTERS[1][8] ), .B1(n845), .B2(
        \REGISTERS[31][8] ), .ZN(n363) );
  AOI22_X1 U451 ( .A1(n844), .A2(\REGISTERS[27][8] ), .B1(n11), .B2(
        \REGISTERS[3][8] ), .ZN(n362) );
  NAND4_X1 U452 ( .A1(n365), .A2(n364), .A3(n363), .A4(n362), .ZN(n376) );
  AOI22_X1 U453 ( .A1(n870), .A2(\REGISTERS[21][8] ), .B1(n3), .B2(
        \REGISTERS[2][8] ), .ZN(n369) );
  AOI22_X1 U454 ( .A1(n6), .A2(\REGISTERS[24][8] ), .B1(n13), .B2(
        \REGISTERS[12][8] ), .ZN(n368) );
  AOI22_X1 U455 ( .A1(n16), .A2(\REGISTERS[6][8] ), .B1(n23), .B2(
        \REGISTERS[16][8] ), .ZN(n367) );
  AOI22_X1 U456 ( .A1(n10), .A2(\REGISTERS[17][8] ), .B1(n24), .B2(
        \REGISTERS[5][8] ), .ZN(n366) );
  NAND4_X1 U457 ( .A1(n369), .A2(n368), .A3(n367), .A4(n366), .ZN(n375) );
  AOI22_X1 U458 ( .A1(n869), .A2(\REGISTERS[18][8] ), .B1(n853), .B2(
        \REGISTERS[9][8] ), .ZN(n373) );
  AOI22_X1 U459 ( .A1(n25), .A2(\REGISTERS[15][8] ), .B1(n17), .B2(
        \REGISTERS[20][8] ), .ZN(n372) );
  AOI22_X1 U460 ( .A1(n842), .A2(\REGISTERS[23][8] ), .B1(n15), .B2(
        \REGISTERS[22][8] ), .ZN(n371) );
  AOI22_X1 U461 ( .A1(n31), .A2(\REGISTERS[10][8] ), .B1(n29), .B2(
        \REGISTERS[11][8] ), .ZN(n370) );
  NAND4_X1 U462 ( .A1(n373), .A2(n372), .A3(n371), .A4(n370), .ZN(n374) );
  NOR4_X1 U463 ( .A1(n377), .A2(n376), .A3(n375), .A4(n374), .ZN(n378) );
  AOI22_X1 U464 ( .A1(n894), .A2(n2675), .B1(n378), .B2(n36), .ZN(N255) );
  AOI22_X1 U465 ( .A1(n20), .A2(\REGISTERS[8][9] ), .B1(n18), .B2(
        \REGISTERS[14][9] ), .ZN(n382) );
  AOI22_X1 U466 ( .A1(n865), .A2(\REGISTERS[20][9] ), .B1(n15), .B2(
        \REGISTERS[22][9] ), .ZN(n381) );
  AOI22_X1 U467 ( .A1(n22), .A2(\REGISTERS[21][9] ), .B1(n21), .B2(
        \REGISTERS[18][9] ), .ZN(n380) );
  AOI22_X1 U468 ( .A1(n31), .A2(\REGISTERS[10][9] ), .B1(n25), .B2(
        \REGISTERS[15][9] ), .ZN(n379) );
  NAND4_X1 U469 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(n398) );
  AOI22_X1 U470 ( .A1(n858), .A2(\REGISTERS[29][9] ), .B1(n16), .B2(
        \REGISTERS[6][9] ), .ZN(n386) );
  AOI22_X1 U471 ( .A1(n872), .A2(\REGISTERS[5][9] ), .B1(n845), .B2(
        \REGISTERS[31][9] ), .ZN(n385) );
  AOI22_X1 U472 ( .A1(n855), .A2(\REGISTERS[3][9] ), .B1(n853), .B2(
        \REGISTERS[9][9] ), .ZN(n384) );
  AOI22_X1 U473 ( .A1(n841), .A2(\REGISTERS[0][9] ), .B1(n7), .B2(
        \REGISTERS[19][9] ), .ZN(n383) );
  NAND4_X1 U474 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(n397) );
  AOI22_X1 U475 ( .A1(n880), .A2(\REGISTERS[30][9] ), .B1(n3), .B2(
        \REGISTERS[2][9] ), .ZN(n390) );
  AOI22_X1 U476 ( .A1(n844), .A2(\REGISTERS[27][9] ), .B1(n29), .B2(
        \REGISTERS[11][9] ), .ZN(n389) );
  AOI22_X1 U477 ( .A1(n879), .A2(\REGISTERS[26][9] ), .B1(n19), .B2(
        \REGISTERS[4][9] ), .ZN(n388) );
  AOI22_X1 U478 ( .A1(n848), .A2(\REGISTERS[1][9] ), .B1(n6), .B2(
        \REGISTERS[24][9] ), .ZN(n387) );
  NAND4_X1 U479 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(n396) );
  AOI22_X1 U480 ( .A1(n10), .A2(\REGISTERS[17][9] ), .B1(n13), .B2(
        \REGISTERS[12][9] ), .ZN(n394) );
  AOI22_X1 U481 ( .A1(n12), .A2(\REGISTERS[28][9] ), .B1(n2), .B2(
        \REGISTERS[23][9] ), .ZN(n393) );
  AOI22_X1 U482 ( .A1(n878), .A2(\REGISTERS[7][9] ), .B1(n23), .B2(
        \REGISTERS[16][9] ), .ZN(n392) );
  AOI22_X1 U483 ( .A1(n32), .A2(\REGISTERS[13][9] ), .B1(n30), .B2(
        \REGISTERS[25][9] ), .ZN(n391) );
  NAND4_X1 U484 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(n395) );
  NOR4_X1 U485 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(n399) );
  AOI22_X1 U486 ( .A1(n894), .A2(n2674), .B1(n399), .B2(n35), .ZN(N256) );
  AOI22_X1 U487 ( .A1(n848), .A2(\REGISTERS[1][10] ), .B1(n859), .B2(
        \REGISTERS[22][10] ), .ZN(n403) );
  AOI22_X1 U488 ( .A1(n846), .A2(\REGISTERS[24][10] ), .B1(n845), .B2(
        \REGISTERS[31][10] ), .ZN(n402) );
  AOI22_X1 U489 ( .A1(n18), .A2(\REGISTERS[14][10] ), .B1(n857), .B2(
        \REGISTERS[12][10] ), .ZN(n401) );
  AOI22_X1 U490 ( .A1(n22), .A2(\REGISTERS[21][10] ), .B1(n871), .B2(
        \REGISTERS[16][10] ), .ZN(n400) );
  NAND4_X1 U491 ( .A1(n403), .A2(n402), .A3(n401), .A4(n400), .ZN(n419) );
  AOI22_X1 U492 ( .A1(n31), .A2(\REGISTERS[10][10] ), .B1(n24), .B2(
        \REGISTERS[5][10] ), .ZN(n407) );
  AOI22_X1 U493 ( .A1(n25), .A2(\REGISTERS[15][10] ), .B1(n2), .B2(
        \REGISTERS[23][10] ), .ZN(n406) );
  AOI22_X1 U494 ( .A1(n844), .A2(\REGISTERS[27][10] ), .B1(n17), .B2(
        \REGISTERS[20][10] ), .ZN(n405) );
  AOI22_X1 U495 ( .A1(n882), .A2(\REGISTERS[25][10] ), .B1(n3), .B2(
        \REGISTERS[2][10] ), .ZN(n404) );
  NAND4_X1 U496 ( .A1(n407), .A2(n406), .A3(n405), .A4(n404), .ZN(n418) );
  AOI22_X1 U497 ( .A1(n10), .A2(\REGISTERS[17][10] ), .B1(n16), .B2(
        \REGISTERS[6][10] ), .ZN(n411) );
  AOI22_X1 U498 ( .A1(n28), .A2(\REGISTERS[30][10] ), .B1(n19), .B2(
        \REGISTERS[4][10] ), .ZN(n410) );
  AOI22_X1 U499 ( .A1(n12), .A2(\REGISTERS[28][10] ), .B1(n29), .B2(
        \REGISTERS[11][10] ), .ZN(n409) );
  AOI22_X1 U500 ( .A1(n878), .A2(\REGISTERS[7][10] ), .B1(n11), .B2(
        \REGISTERS[3][10] ), .ZN(n408) );
  NAND4_X1 U501 ( .A1(n411), .A2(n410), .A3(n409), .A4(n408), .ZN(n417) );
  AOI22_X1 U502 ( .A1(n32), .A2(\REGISTERS[13][10] ), .B1(n7), .B2(
        \REGISTERS[19][10] ), .ZN(n415) );
  AOI22_X1 U503 ( .A1(n841), .A2(\REGISTERS[0][10] ), .B1(n853), .B2(
        \REGISTERS[9][10] ), .ZN(n414) );
  AOI22_X1 U504 ( .A1(n27), .A2(\REGISTERS[26][10] ), .B1(n14), .B2(
        \REGISTERS[29][10] ), .ZN(n413) );
  AOI22_X1 U505 ( .A1(n20), .A2(\REGISTERS[8][10] ), .B1(n21), .B2(
        \REGISTERS[18][10] ), .ZN(n412) );
  NAND4_X1 U506 ( .A1(n415), .A2(n414), .A3(n413), .A4(n412), .ZN(n416) );
  NOR4_X1 U507 ( .A1(n419), .A2(n418), .A3(n417), .A4(n416), .ZN(n420) );
  AOI22_X1 U508 ( .A1(n894), .A2(n2661), .B1(n420), .B2(n36), .ZN(N257) );
  AOI22_X1 U509 ( .A1(n10), .A2(\REGISTERS[17][11] ), .B1(n13), .B2(
        \REGISTERS[12][11] ), .ZN(n424) );
  AOI22_X1 U510 ( .A1(n14), .A2(\REGISTERS[29][11] ), .B1(n853), .B2(
        \REGISTERS[9][11] ), .ZN(n423) );
  AOI22_X1 U511 ( .A1(n31), .A2(\REGISTERS[10][11] ), .B1(n2), .B2(
        \REGISTERS[23][11] ), .ZN(n422) );
  AOI22_X1 U512 ( .A1(n22), .A2(\REGISTERS[21][11] ), .B1(n21), .B2(
        \REGISTERS[18][11] ), .ZN(n421) );
  NAND4_X1 U513 ( .A1(n424), .A2(n423), .A3(n422), .A4(n421), .ZN(n440) );
  AOI22_X1 U514 ( .A1(n19), .A2(\REGISTERS[4][11] ), .B1(n871), .B2(
        \REGISTERS[16][11] ), .ZN(n428) );
  AOI22_X1 U515 ( .A1(n12), .A2(\REGISTERS[28][11] ), .B1(n847), .B2(
        \REGISTERS[19][11] ), .ZN(n427) );
  AOI22_X1 U516 ( .A1(n27), .A2(\REGISTERS[26][11] ), .B1(n11), .B2(
        \REGISTERS[3][11] ), .ZN(n426) );
  AOI22_X1 U517 ( .A1(n30), .A2(\REGISTERS[25][11] ), .B1(n8), .B2(
        \REGISTERS[1][11] ), .ZN(n425) );
  NAND4_X1 U518 ( .A1(n428), .A2(n427), .A3(n426), .A4(n425), .ZN(n439) );
  AOI22_X1 U519 ( .A1(n878), .A2(\REGISTERS[7][11] ), .B1(n32), .B2(
        \REGISTERS[13][11] ), .ZN(n432) );
  AOI22_X1 U520 ( .A1(n28), .A2(\REGISTERS[30][11] ), .B1(n16), .B2(
        \REGISTERS[6][11] ), .ZN(n431) );
  AOI22_X1 U521 ( .A1(n20), .A2(\REGISTERS[8][11] ), .B1(n845), .B2(
        \REGISTERS[31][11] ), .ZN(n430) );
  AOI22_X1 U522 ( .A1(n844), .A2(\REGISTERS[27][11] ), .B1(n17), .B2(
        \REGISTERS[20][11] ), .ZN(n429) );
  NAND4_X1 U523 ( .A1(n432), .A2(n431), .A3(n430), .A4(n429), .ZN(n438) );
  AOI22_X1 U524 ( .A1(n841), .A2(\REGISTERS[0][11] ), .B1(n3), .B2(
        \REGISTERS[2][11] ), .ZN(n436) );
  AOI22_X1 U525 ( .A1(n25), .A2(\REGISTERS[15][11] ), .B1(n29), .B2(
        \REGISTERS[11][11] ), .ZN(n435) );
  AOI22_X1 U526 ( .A1(n872), .A2(\REGISTERS[5][11] ), .B1(n859), .B2(
        \REGISTERS[22][11] ), .ZN(n434) );
  AOI22_X1 U527 ( .A1(n866), .A2(\REGISTERS[14][11] ), .B1(n6), .B2(
        \REGISTERS[24][11] ), .ZN(n433) );
  NAND4_X1 U528 ( .A1(n436), .A2(n435), .A3(n434), .A4(n433), .ZN(n437) );
  NOR4_X1 U529 ( .A1(n440), .A2(n439), .A3(n438), .A4(n437), .ZN(n441) );
  AOI22_X1 U530 ( .A1(n894), .A2(n114), .B1(n441), .B2(n35), .ZN(N258) );
  AOI22_X1 U531 ( .A1(n22), .A2(\REGISTERS[21][12] ), .B1(n17), .B2(
        \REGISTERS[20][12] ), .ZN(n445) );
  AOI22_X1 U532 ( .A1(n27), .A2(\REGISTERS[26][12] ), .B1(n5), .B2(
        \REGISTERS[31][12] ), .ZN(n444) );
  AOI22_X1 U533 ( .A1(n28), .A2(\REGISTERS[30][12] ), .B1(n11), .B2(
        \REGISTERS[3][12] ), .ZN(n443) );
  AOI22_X1 U534 ( .A1(n30), .A2(\REGISTERS[25][12] ), .B1(n1), .B2(
        \REGISTERS[0][12] ), .ZN(n442) );
  NAND4_X1 U535 ( .A1(n445), .A2(n444), .A3(n443), .A4(n442), .ZN(n461) );
  AOI22_X1 U536 ( .A1(n16), .A2(\REGISTERS[6][12] ), .B1(n3), .B2(
        \REGISTERS[2][12] ), .ZN(n449) );
  AOI22_X1 U537 ( .A1(n844), .A2(\REGISTERS[27][12] ), .B1(n881), .B2(
        \REGISTERS[11][12] ), .ZN(n448) );
  AOI22_X1 U538 ( .A1(n10), .A2(\REGISTERS[17][12] ), .B1(n18), .B2(
        \REGISTERS[14][12] ), .ZN(n447) );
  AOI22_X1 U539 ( .A1(n848), .A2(\REGISTERS[1][12] ), .B1(n9), .B2(
        \REGISTERS[9][12] ), .ZN(n446) );
  NAND4_X1 U540 ( .A1(n449), .A2(n448), .A3(n447), .A4(n446), .ZN(n460) );
  AOI22_X1 U541 ( .A1(n25), .A2(\REGISTERS[15][12] ), .B1(n847), .B2(
        \REGISTERS[19][12] ), .ZN(n453) );
  AOI22_X1 U542 ( .A1(n867), .A2(\REGISTERS[4][12] ), .B1(n23), .B2(
        \REGISTERS[16][12] ), .ZN(n452) );
  AOI22_X1 U543 ( .A1(n32), .A2(\REGISTERS[13][12] ), .B1(n6), .B2(
        \REGISTERS[24][12] ), .ZN(n451) );
  AOI22_X1 U544 ( .A1(n20), .A2(\REGISTERS[8][12] ), .B1(n2), .B2(
        \REGISTERS[23][12] ), .ZN(n450) );
  NAND4_X1 U545 ( .A1(n453), .A2(n452), .A3(n451), .A4(n450), .ZN(n459) );
  AOI22_X1 U546 ( .A1(n14), .A2(\REGISTERS[29][12] ), .B1(n21), .B2(
        \REGISTERS[18][12] ), .ZN(n457) );
  AOI22_X1 U547 ( .A1(n12), .A2(\REGISTERS[28][12] ), .B1(n31), .B2(
        \REGISTERS[10][12] ), .ZN(n456) );
  AOI22_X1 U548 ( .A1(n26), .A2(\REGISTERS[7][12] ), .B1(n15), .B2(
        \REGISTERS[22][12] ), .ZN(n455) );
  AOI22_X1 U549 ( .A1(n857), .A2(\REGISTERS[12][12] ), .B1(n24), .B2(
        \REGISTERS[5][12] ), .ZN(n454) );
  NAND4_X1 U550 ( .A1(n457), .A2(n456), .A3(n455), .A4(n454), .ZN(n458) );
  NOR4_X1 U551 ( .A1(n461), .A2(n460), .A3(n459), .A4(n458), .ZN(n462) );
  AOI22_X1 U552 ( .A1(n33), .A2(n2666), .B1(n462), .B2(n36), .ZN(N259) );
  AOI22_X1 U553 ( .A1(n846), .A2(\REGISTERS[24][13] ), .B1(n857), .B2(
        \REGISTERS[12][13] ), .ZN(n466) );
  AOI22_X1 U554 ( .A1(n10), .A2(\REGISTERS[17][13] ), .B1(n31), .B2(
        \REGISTERS[10][13] ), .ZN(n465) );
  AOI22_X1 U555 ( .A1(n30), .A2(\REGISTERS[25][13] ), .B1(n23), .B2(
        \REGISTERS[16][13] ), .ZN(n464) );
  AOI22_X1 U556 ( .A1(n12), .A2(\REGISTERS[28][13] ), .B1(n1), .B2(
        \REGISTERS[0][13] ), .ZN(n463) );
  NAND4_X1 U557 ( .A1(n466), .A2(n465), .A3(n464), .A4(n463), .ZN(n482) );
  AOI22_X1 U558 ( .A1(n843), .A2(\REGISTERS[2][13] ), .B1(n5), .B2(
        \REGISTERS[31][13] ), .ZN(n470) );
  AOI22_X1 U559 ( .A1(n2), .A2(\REGISTERS[23][13] ), .B1(n15), .B2(
        \REGISTERS[22][13] ), .ZN(n469) );
  AOI22_X1 U560 ( .A1(n32), .A2(\REGISTERS[13][13] ), .B1(n881), .B2(
        \REGISTERS[11][13] ), .ZN(n468) );
  AOI22_X1 U561 ( .A1(n847), .A2(\REGISTERS[19][13] ), .B1(n9), .B2(
        \REGISTERS[9][13] ), .ZN(n467) );
  NAND4_X1 U562 ( .A1(n470), .A2(n469), .A3(n468), .A4(n467), .ZN(n481) );
  AOI22_X1 U563 ( .A1(n877), .A2(\REGISTERS[15][13] ), .B1(n4), .B2(
        \REGISTERS[27][13] ), .ZN(n474) );
  AOI22_X1 U564 ( .A1(n868), .A2(\REGISTERS[8][13] ), .B1(n872), .B2(
        \REGISTERS[5][13] ), .ZN(n473) );
  AOI22_X1 U565 ( .A1(n14), .A2(\REGISTERS[29][13] ), .B1(n865), .B2(
        \REGISTERS[20][13] ), .ZN(n472) );
  AOI22_X1 U566 ( .A1(n860), .A2(\REGISTERS[6][13] ), .B1(n18), .B2(
        \REGISTERS[14][13] ), .ZN(n471) );
  NAND4_X1 U567 ( .A1(n474), .A2(n473), .A3(n472), .A4(n471), .ZN(n480) );
  AOI22_X1 U568 ( .A1(n848), .A2(\REGISTERS[1][13] ), .B1(n855), .B2(
        \REGISTERS[3][13] ), .ZN(n478) );
  AOI22_X1 U569 ( .A1(n26), .A2(\REGISTERS[7][13] ), .B1(n19), .B2(
        \REGISTERS[4][13] ), .ZN(n477) );
  AOI22_X1 U570 ( .A1(n27), .A2(\REGISTERS[26][13] ), .B1(n21), .B2(
        \REGISTERS[18][13] ), .ZN(n476) );
  AOI22_X1 U571 ( .A1(n28), .A2(\REGISTERS[30][13] ), .B1(n22), .B2(
        \REGISTERS[21][13] ), .ZN(n475) );
  NAND4_X1 U572 ( .A1(n478), .A2(n477), .A3(n476), .A4(n475), .ZN(n479) );
  NOR4_X1 U573 ( .A1(n482), .A2(n481), .A3(n480), .A4(n479), .ZN(n483) );
  AOI22_X1 U574 ( .A1(n33), .A2(n110), .B1(n483), .B2(n35), .ZN(N260) );
  AOI22_X1 U575 ( .A1(n10), .A2(\REGISTERS[17][14] ), .B1(n23), .B2(
        \REGISTERS[16][14] ), .ZN(n487) );
  AOI22_X1 U576 ( .A1(n30), .A2(\REGISTERS[25][14] ), .B1(n865), .B2(
        \REGISTERS[20][14] ), .ZN(n486) );
  AOI22_X1 U577 ( .A1(n14), .A2(\REGISTERS[29][14] ), .B1(n1), .B2(
        \REGISTERS[0][14] ), .ZN(n485) );
  AOI22_X1 U578 ( .A1(n7), .A2(\REGISTERS[19][14] ), .B1(n13), .B2(
        \REGISTERS[12][14] ), .ZN(n484) );
  NAND4_X1 U579 ( .A1(n487), .A2(n486), .A3(n485), .A4(n484), .ZN(n503) );
  AOI22_X1 U580 ( .A1(n867), .A2(\REGISTERS[4][14] ), .B1(n15), .B2(
        \REGISTERS[22][14] ), .ZN(n491) );
  AOI22_X1 U581 ( .A1(n27), .A2(\REGISTERS[26][14] ), .B1(n25), .B2(
        \REGISTERS[15][14] ), .ZN(n490) );
  AOI22_X1 U582 ( .A1(n860), .A2(\REGISTERS[6][14] ), .B1(n6), .B2(
        \REGISTERS[24][14] ), .ZN(n489) );
  AOI22_X1 U583 ( .A1(n881), .A2(\REGISTERS[11][14] ), .B1(n9), .B2(
        \REGISTERS[9][14] ), .ZN(n488) );
  NAND4_X1 U584 ( .A1(n491), .A2(n490), .A3(n489), .A4(n488), .ZN(n502) );
  AOI22_X1 U585 ( .A1(n12), .A2(\REGISTERS[28][14] ), .B1(n8), .B2(
        \REGISTERS[1][14] ), .ZN(n495) );
  AOI22_X1 U586 ( .A1(n843), .A2(\REGISTERS[2][14] ), .B1(n5), .B2(
        \REGISTERS[31][14] ), .ZN(n494) );
  AOI22_X1 U587 ( .A1(n26), .A2(\REGISTERS[7][14] ), .B1(n2), .B2(
        \REGISTERS[23][14] ), .ZN(n493) );
  AOI22_X1 U588 ( .A1(n28), .A2(\REGISTERS[30][14] ), .B1(n4), .B2(
        \REGISTERS[27][14] ), .ZN(n492) );
  NAND4_X1 U589 ( .A1(n495), .A2(n494), .A3(n493), .A4(n492), .ZN(n501) );
  AOI22_X1 U590 ( .A1(n31), .A2(\REGISTERS[10][14] ), .B1(n20), .B2(
        \REGISTERS[8][14] ), .ZN(n499) );
  AOI22_X1 U591 ( .A1(n869), .A2(\REGISTERS[18][14] ), .B1(n872), .B2(
        \REGISTERS[5][14] ), .ZN(n498) );
  AOI22_X1 U592 ( .A1(n870), .A2(\REGISTERS[21][14] ), .B1(n18), .B2(
        \REGISTERS[14][14] ), .ZN(n497) );
  AOI22_X1 U593 ( .A1(n32), .A2(\REGISTERS[13][14] ), .B1(n855), .B2(
        \REGISTERS[3][14] ), .ZN(n496) );
  NAND4_X1 U594 ( .A1(n499), .A2(n498), .A3(n497), .A4(n496), .ZN(n500) );
  NOR4_X1 U595 ( .A1(n503), .A2(n502), .A3(n501), .A4(n500), .ZN(n504) );
  AOI22_X1 U596 ( .A1(n33), .A2(n2660), .B1(n504), .B2(n36), .ZN(N261) );
  AOI22_X1 U597 ( .A1(n4), .A2(\REGISTERS[27][15] ), .B1(n17), .B2(
        \REGISTERS[20][15] ), .ZN(n508) );
  AOI22_X1 U598 ( .A1(n30), .A2(\REGISTERS[25][15] ), .B1(n14), .B2(
        \REGISTERS[29][15] ), .ZN(n507) );
  AOI22_X1 U599 ( .A1(n855), .A2(\REGISTERS[3][15] ), .B1(n13), .B2(
        \REGISTERS[12][15] ), .ZN(n506) );
  AOI22_X1 U600 ( .A1(n32), .A2(\REGISTERS[13][15] ), .B1(n12), .B2(
        \REGISTERS[28][15] ), .ZN(n505) );
  NAND4_X1 U601 ( .A1(n508), .A2(n507), .A3(n506), .A4(n505), .ZN(n524) );
  AOI22_X1 U602 ( .A1(n877), .A2(\REGISTERS[15][15] ), .B1(n21), .B2(
        \REGISTERS[18][15] ), .ZN(n512) );
  AOI22_X1 U603 ( .A1(n847), .A2(\REGISTERS[19][15] ), .B1(n9), .B2(
        \REGISTERS[9][15] ), .ZN(n511) );
  AOI22_X1 U604 ( .A1(n859), .A2(\REGISTERS[22][15] ), .B1(n23), .B2(
        \REGISTERS[16][15] ), .ZN(n510) );
  AOI22_X1 U605 ( .A1(n841), .A2(\REGISTERS[0][15] ), .B1(n8), .B2(
        \REGISTERS[1][15] ), .ZN(n509) );
  NAND4_X1 U606 ( .A1(n512), .A2(n511), .A3(n510), .A4(n509), .ZN(n523) );
  AOI22_X1 U607 ( .A1(n26), .A2(\REGISTERS[7][15] ), .B1(n18), .B2(
        \REGISTERS[14][15] ), .ZN(n516) );
  AOI22_X1 U608 ( .A1(n22), .A2(\REGISTERS[21][15] ), .B1(n16), .B2(
        \REGISTERS[6][15] ), .ZN(n515) );
  AOI22_X1 U609 ( .A1(n846), .A2(\REGISTERS[24][15] ), .B1(n24), .B2(
        \REGISTERS[5][15] ), .ZN(n514) );
  AOI22_X1 U610 ( .A1(n10), .A2(\REGISTERS[17][15] ), .B1(n843), .B2(
        \REGISTERS[2][15] ), .ZN(n513) );
  NAND4_X1 U611 ( .A1(n516), .A2(n515), .A3(n514), .A4(n513), .ZN(n522) );
  AOI22_X1 U612 ( .A1(n868), .A2(\REGISTERS[8][15] ), .B1(n5), .B2(
        \REGISTERS[31][15] ), .ZN(n520) );
  AOI22_X1 U613 ( .A1(n28), .A2(\REGISTERS[30][15] ), .B1(n2), .B2(
        \REGISTERS[23][15] ), .ZN(n519) );
  AOI22_X1 U614 ( .A1(n867), .A2(\REGISTERS[4][15] ), .B1(n29), .B2(
        \REGISTERS[11][15] ), .ZN(n518) );
  AOI22_X1 U615 ( .A1(n27), .A2(\REGISTERS[26][15] ), .B1(n31), .B2(
        \REGISTERS[10][15] ), .ZN(n517) );
  NAND4_X1 U616 ( .A1(n520), .A2(n519), .A3(n518), .A4(n517), .ZN(n521) );
  NOR4_X1 U617 ( .A1(n524), .A2(n523), .A3(n522), .A4(n521), .ZN(n525) );
  AOI22_X1 U618 ( .A1(n33), .A2(n2658), .B1(n525), .B2(n35), .ZN(N262) );
  AOI22_X1 U619 ( .A1(n854), .A2(\REGISTERS[17][16] ), .B1(n23), .B2(
        \REGISTERS[16][16] ), .ZN(n529) );
  AOI22_X1 U620 ( .A1(n30), .A2(\REGISTERS[25][16] ), .B1(n13), .B2(
        \REGISTERS[12][16] ), .ZN(n528) );
  AOI22_X1 U621 ( .A1(n26), .A2(\REGISTERS[7][16] ), .B1(n869), .B2(
        \REGISTERS[18][16] ), .ZN(n527) );
  AOI22_X1 U622 ( .A1(n867), .A2(\REGISTERS[4][16] ), .B1(n5), .B2(
        \REGISTERS[31][16] ), .ZN(n526) );
  NAND4_X1 U623 ( .A1(n529), .A2(n528), .A3(n527), .A4(n526), .ZN(n545) );
  AOI22_X1 U624 ( .A1(n860), .A2(\REGISTERS[6][16] ), .B1(n9), .B2(
        \REGISTERS[9][16] ), .ZN(n533) );
  AOI22_X1 U625 ( .A1(n32), .A2(\REGISTERS[13][16] ), .B1(n843), .B2(
        \REGISTERS[2][16] ), .ZN(n532) );
  AOI22_X1 U626 ( .A1(n14), .A2(\REGISTERS[29][16] ), .B1(n4), .B2(
        \REGISTERS[27][16] ), .ZN(n531) );
  AOI22_X1 U627 ( .A1(n866), .A2(\REGISTERS[14][16] ), .B1(n7), .B2(
        \REGISTERS[19][16] ), .ZN(n530) );
  NAND4_X1 U628 ( .A1(n533), .A2(n532), .A3(n531), .A4(n530), .ZN(n544) );
  AOI22_X1 U629 ( .A1(n877), .A2(\REGISTERS[15][16] ), .B1(n17), .B2(
        \REGISTERS[20][16] ), .ZN(n537) );
  AOI22_X1 U630 ( .A1(n2), .A2(\REGISTERS[23][16] ), .B1(n29), .B2(
        \REGISTERS[11][16] ), .ZN(n536) );
  AOI22_X1 U631 ( .A1(n31), .A2(\REGISTERS[10][16] ), .B1(n1), .B2(
        \REGISTERS[0][16] ), .ZN(n535) );
  AOI22_X1 U632 ( .A1(n8), .A2(\REGISTERS[1][16] ), .B1(n15), .B2(
        \REGISTERS[22][16] ), .ZN(n534) );
  NAND4_X1 U633 ( .A1(n537), .A2(n536), .A3(n535), .A4(n534), .ZN(n543) );
  AOI22_X1 U634 ( .A1(n28), .A2(\REGISTERS[30][16] ), .B1(n20), .B2(
        \REGISTERS[8][16] ), .ZN(n541) );
  AOI22_X1 U635 ( .A1(n27), .A2(\REGISTERS[26][16] ), .B1(n24), .B2(
        \REGISTERS[5][16] ), .ZN(n540) );
  AOI22_X1 U636 ( .A1(n12), .A2(\REGISTERS[28][16] ), .B1(n22), .B2(
        \REGISTERS[21][16] ), .ZN(n539) );
  AOI22_X1 U637 ( .A1(n846), .A2(\REGISTERS[24][16] ), .B1(n11), .B2(
        \REGISTERS[3][16] ), .ZN(n538) );
  NAND4_X1 U638 ( .A1(n541), .A2(n540), .A3(n539), .A4(n538), .ZN(n542) );
  NOR4_X1 U639 ( .A1(n545), .A2(n544), .A3(n543), .A4(n542), .ZN(n546) );
  AOI22_X1 U640 ( .A1(n33), .A2(n2668), .B1(n546), .B2(n36), .ZN(N263) );
  AOI22_X1 U641 ( .A1(n877), .A2(\REGISTERS[15][17] ), .B1(n24), .B2(
        \REGISTERS[5][17] ), .ZN(n550) );
  AOI22_X1 U642 ( .A1(n32), .A2(\REGISTERS[13][17] ), .B1(n3), .B2(
        \REGISTERS[2][17] ), .ZN(n549) );
  AOI22_X1 U643 ( .A1(n860), .A2(\REGISTERS[6][17] ), .B1(n5), .B2(
        \REGISTERS[31][17] ), .ZN(n548) );
  AOI22_X1 U644 ( .A1(n869), .A2(\REGISTERS[18][17] ), .B1(n6), .B2(
        \REGISTERS[24][17] ), .ZN(n547) );
  NAND4_X1 U645 ( .A1(n550), .A2(n549), .A3(n548), .A4(n547), .ZN(n566) );
  AOI22_X1 U646 ( .A1(n855), .A2(\REGISTERS[3][17] ), .B1(n15), .B2(
        \REGISTERS[22][17] ), .ZN(n554) );
  AOI22_X1 U647 ( .A1(n14), .A2(\REGISTERS[29][17] ), .B1(n18), .B2(
        \REGISTERS[14][17] ), .ZN(n553) );
  AOI22_X1 U648 ( .A1(n1), .A2(\REGISTERS[0][17] ), .B1(n23), .B2(
        \REGISTERS[16][17] ), .ZN(n552) );
  AOI22_X1 U649 ( .A1(n854), .A2(\REGISTERS[17][17] ), .B1(n31), .B2(
        \REGISTERS[10][17] ), .ZN(n551) );
  NAND4_X1 U650 ( .A1(n554), .A2(n553), .A3(n552), .A4(n551), .ZN(n565) );
  AOI22_X1 U651 ( .A1(n870), .A2(\REGISTERS[21][17] ), .B1(n9), .B2(
        \REGISTERS[9][17] ), .ZN(n558) );
  AOI22_X1 U652 ( .A1(n28), .A2(\REGISTERS[30][17] ), .B1(n27), .B2(
        \REGISTERS[26][17] ), .ZN(n557) );
  AOI22_X1 U653 ( .A1(n844), .A2(\REGISTERS[27][17] ), .B1(n19), .B2(
        \REGISTERS[4][17] ), .ZN(n556) );
  AOI22_X1 U654 ( .A1(n30), .A2(\REGISTERS[25][17] ), .B1(n7), .B2(
        \REGISTERS[19][17] ), .ZN(n555) );
  NAND4_X1 U655 ( .A1(n558), .A2(n557), .A3(n556), .A4(n555), .ZN(n564) );
  AOI22_X1 U656 ( .A1(n856), .A2(\REGISTERS[28][17] ), .B1(n29), .B2(
        \REGISTERS[11][17] ), .ZN(n562) );
  AOI22_X1 U657 ( .A1(n26), .A2(\REGISTERS[7][17] ), .B1(n17), .B2(
        \REGISTERS[20][17] ), .ZN(n561) );
  AOI22_X1 U658 ( .A1(n868), .A2(\REGISTERS[8][17] ), .B1(n2), .B2(
        \REGISTERS[23][17] ), .ZN(n560) );
  AOI22_X1 U659 ( .A1(n848), .A2(\REGISTERS[1][17] ), .B1(n13), .B2(
        \REGISTERS[12][17] ), .ZN(n559) );
  NAND4_X1 U660 ( .A1(n562), .A2(n561), .A3(n560), .A4(n559), .ZN(n563) );
  NOR4_X1 U661 ( .A1(n566), .A2(n565), .A3(n564), .A4(n563), .ZN(n567) );
  AOI22_X1 U662 ( .A1(n33), .A2(n2667), .B1(n567), .B2(n35), .ZN(N264) );
  AOI22_X1 U663 ( .A1(n860), .A2(\REGISTERS[6][18] ), .B1(n29), .B2(
        \REGISTERS[11][18] ), .ZN(n571) );
  AOI22_X1 U664 ( .A1(n884), .A2(\REGISTERS[13][18] ), .B1(n1), .B2(
        \REGISTERS[0][18] ), .ZN(n570) );
  AOI22_X1 U665 ( .A1(n872), .A2(\REGISTERS[5][18] ), .B1(n15), .B2(
        \REGISTERS[22][18] ), .ZN(n569) );
  AOI22_X1 U666 ( .A1(n14), .A2(\REGISTERS[29][18] ), .B1(n6), .B2(
        \REGISTERS[24][18] ), .ZN(n568) );
  NAND4_X1 U667 ( .A1(n571), .A2(n570), .A3(n569), .A4(n568), .ZN(n587) );
  AOI22_X1 U668 ( .A1(n28), .A2(\REGISTERS[30][18] ), .B1(n12), .B2(
        \REGISTERS[28][18] ), .ZN(n575) );
  AOI22_X1 U669 ( .A1(n866), .A2(\REGISTERS[14][18] ), .B1(n13), .B2(
        \REGISTERS[12][18] ), .ZN(n574) );
  AOI22_X1 U670 ( .A1(n868), .A2(\REGISTERS[8][18] ), .B1(n23), .B2(
        \REGISTERS[16][18] ), .ZN(n573) );
  AOI22_X1 U671 ( .A1(n842), .A2(\REGISTERS[23][18] ), .B1(n9), .B2(
        \REGISTERS[9][18] ), .ZN(n572) );
  NAND4_X1 U672 ( .A1(n575), .A2(n574), .A3(n573), .A4(n572), .ZN(n586) );
  AOI22_X1 U673 ( .A1(n855), .A2(\REGISTERS[3][18] ), .B1(n5), .B2(
        \REGISTERS[31][18] ), .ZN(n579) );
  AOI22_X1 U674 ( .A1(n31), .A2(\REGISTERS[10][18] ), .B1(n7), .B2(
        \REGISTERS[19][18] ), .ZN(n578) );
  AOI22_X1 U675 ( .A1(n26), .A2(\REGISTERS[7][18] ), .B1(n25), .B2(
        \REGISTERS[15][18] ), .ZN(n577) );
  AOI22_X1 U676 ( .A1(n27), .A2(\REGISTERS[26][18] ), .B1(n22), .B2(
        \REGISTERS[21][18] ), .ZN(n576) );
  NAND4_X1 U677 ( .A1(n579), .A2(n578), .A3(n577), .A4(n576), .ZN(n585) );
  AOI22_X1 U678 ( .A1(n865), .A2(\REGISTERS[20][18] ), .B1(n19), .B2(
        \REGISTERS[4][18] ), .ZN(n583) );
  AOI22_X1 U679 ( .A1(n30), .A2(\REGISTERS[25][18] ), .B1(n8), .B2(
        \REGISTERS[1][18] ), .ZN(n582) );
  AOI22_X1 U680 ( .A1(n854), .A2(\REGISTERS[17][18] ), .B1(n869), .B2(
        \REGISTERS[18][18] ), .ZN(n581) );
  AOI22_X1 U681 ( .A1(n4), .A2(\REGISTERS[27][18] ), .B1(n3), .B2(
        \REGISTERS[2][18] ), .ZN(n580) );
  NAND4_X1 U682 ( .A1(n583), .A2(n582), .A3(n581), .A4(n580), .ZN(n584) );
  NOR4_X1 U683 ( .A1(n587), .A2(n586), .A3(n585), .A4(n584), .ZN(n588) );
  AOI22_X1 U684 ( .A1(n33), .A2(n100), .B1(n588), .B2(n36), .ZN(N265) );
  AOI22_X1 U685 ( .A1(n26), .A2(\REGISTERS[7][19] ), .B1(n4), .B2(
        \REGISTERS[27][19] ), .ZN(n592) );
  AOI22_X1 U686 ( .A1(n866), .A2(\REGISTERS[14][19] ), .B1(n21), .B2(
        \REGISTERS[18][19] ), .ZN(n591) );
  AOI22_X1 U687 ( .A1(n868), .A2(\REGISTERS[8][19] ), .B1(n7), .B2(
        \REGISTERS[19][19] ), .ZN(n590) );
  AOI22_X1 U688 ( .A1(n28), .A2(\REGISTERS[30][19] ), .B1(n29), .B2(
        \REGISTERS[11][19] ), .ZN(n589) );
  NAND4_X1 U689 ( .A1(n592), .A2(n591), .A3(n590), .A4(n589), .ZN(n608) );
  AOI22_X1 U690 ( .A1(n884), .A2(\REGISTERS[13][19] ), .B1(n8), .B2(
        \REGISTERS[1][19] ), .ZN(n596) );
  AOI22_X1 U691 ( .A1(n30), .A2(\REGISTERS[25][19] ), .B1(n15), .B2(
        \REGISTERS[22][19] ), .ZN(n595) );
  AOI22_X1 U692 ( .A1(n867), .A2(\REGISTERS[4][19] ), .B1(n9), .B2(
        \REGISTERS[9][19] ), .ZN(n594) );
  AOI22_X1 U693 ( .A1(n877), .A2(\REGISTERS[15][19] ), .B1(n5), .B2(
        \REGISTERS[31][19] ), .ZN(n593) );
  NAND4_X1 U694 ( .A1(n596), .A2(n595), .A3(n594), .A4(n593), .ZN(n607) );
  AOI22_X1 U695 ( .A1(n883), .A2(\REGISTERS[10][19] ), .B1(n1), .B2(
        \REGISTERS[0][19] ), .ZN(n600) );
  AOI22_X1 U696 ( .A1(n854), .A2(\REGISTERS[17][19] ), .B1(n2), .B2(
        \REGISTERS[23][19] ), .ZN(n599) );
  AOI22_X1 U697 ( .A1(n870), .A2(\REGISTERS[21][19] ), .B1(n17), .B2(
        \REGISTERS[20][19] ), .ZN(n598) );
  AOI22_X1 U698 ( .A1(n11), .A2(\REGISTERS[3][19] ), .B1(n13), .B2(
        \REGISTERS[12][19] ), .ZN(n597) );
  NAND4_X1 U699 ( .A1(n600), .A2(n599), .A3(n598), .A4(n597), .ZN(n606) );
  AOI22_X1 U700 ( .A1(n879), .A2(\REGISTERS[26][19] ), .B1(n23), .B2(
        \REGISTERS[16][19] ), .ZN(n604) );
  AOI22_X1 U701 ( .A1(n846), .A2(\REGISTERS[24][19] ), .B1(n3), .B2(
        \REGISTERS[2][19] ), .ZN(n603) );
  AOI22_X1 U702 ( .A1(n858), .A2(\REGISTERS[29][19] ), .B1(n24), .B2(
        \REGISTERS[5][19] ), .ZN(n602) );
  AOI22_X1 U703 ( .A1(n856), .A2(\REGISTERS[28][19] ), .B1(n16), .B2(
        \REGISTERS[6][19] ), .ZN(n601) );
  NAND4_X1 U704 ( .A1(n604), .A2(n603), .A3(n602), .A4(n601), .ZN(n605) );
  NOR4_X1 U705 ( .A1(n608), .A2(n607), .A3(n606), .A4(n605), .ZN(n609) );
  AOI22_X1 U706 ( .A1(n33), .A2(n2673), .B1(n609), .B2(n36), .ZN(N266) );
  AOI22_X1 U707 ( .A1(n879), .A2(\REGISTERS[26][20] ), .B1(n10), .B2(
        \REGISTERS[17][20] ), .ZN(n613) );
  AOI22_X1 U708 ( .A1(n870), .A2(\REGISTERS[21][20] ), .B1(n8), .B2(
        \REGISTERS[1][20] ), .ZN(n612) );
  AOI22_X1 U709 ( .A1(n26), .A2(\REGISTERS[7][20] ), .B1(n4), .B2(
        \REGISTERS[27][20] ), .ZN(n611) );
  AOI22_X1 U710 ( .A1(n880), .A2(\REGISTERS[30][20] ), .B1(n14), .B2(
        \REGISTERS[29][20] ), .ZN(n610) );
  NAND4_X1 U711 ( .A1(n613), .A2(n612), .A3(n611), .A4(n610), .ZN(n629) );
  AOI22_X1 U712 ( .A1(n883), .A2(\REGISTERS[10][20] ), .B1(n18), .B2(
        \REGISTERS[14][20] ), .ZN(n617) );
  AOI22_X1 U713 ( .A1(n855), .A2(\REGISTERS[3][20] ), .B1(n3), .B2(
        \REGISTERS[2][20] ), .ZN(n616) );
  AOI22_X1 U714 ( .A1(n842), .A2(\REGISTERS[23][20] ), .B1(n15), .B2(
        \REGISTERS[22][20] ), .ZN(n615) );
  AOI22_X1 U715 ( .A1(n847), .A2(\REGISTERS[19][20] ), .B1(n29), .B2(
        \REGISTERS[11][20] ), .ZN(n614) );
  NAND4_X1 U716 ( .A1(n617), .A2(n616), .A3(n615), .A4(n614), .ZN(n628) );
  AOI22_X1 U717 ( .A1(n882), .A2(\REGISTERS[25][20] ), .B1(n13), .B2(
        \REGISTERS[12][20] ), .ZN(n621) );
  AOI22_X1 U718 ( .A1(n25), .A2(\REGISTERS[15][20] ), .B1(n17), .B2(
        \REGISTERS[20][20] ), .ZN(n620) );
  AOI22_X1 U719 ( .A1(n860), .A2(\REGISTERS[6][20] ), .B1(n21), .B2(
        \REGISTERS[18][20] ), .ZN(n619) );
  AOI22_X1 U720 ( .A1(n884), .A2(\REGISTERS[13][20] ), .B1(n12), .B2(
        \REGISTERS[28][20] ), .ZN(n618) );
  NAND4_X1 U721 ( .A1(n621), .A2(n620), .A3(n619), .A4(n618), .ZN(n627) );
  AOI22_X1 U722 ( .A1(n868), .A2(\REGISTERS[8][20] ), .B1(n24), .B2(
        \REGISTERS[5][20] ), .ZN(n625) );
  AOI22_X1 U723 ( .A1(n867), .A2(\REGISTERS[4][20] ), .B1(n853), .B2(
        \REGISTERS[9][20] ), .ZN(n624) );
  AOI22_X1 U724 ( .A1(n1), .A2(\REGISTERS[0][20] ), .B1(n6), .B2(
        \REGISTERS[24][20] ), .ZN(n623) );
  AOI22_X1 U725 ( .A1(n871), .A2(\REGISTERS[16][20] ), .B1(n845), .B2(
        \REGISTERS[31][20] ), .ZN(n622) );
  NAND4_X1 U726 ( .A1(n625), .A2(n624), .A3(n623), .A4(n622), .ZN(n626) );
  NOR4_X1 U727 ( .A1(n629), .A2(n628), .A3(n627), .A4(n626), .ZN(n630) );
  AOI22_X1 U728 ( .A1(n33), .A2(n96), .B1(n630), .B2(n35), .ZN(N267) );
  AOI22_X1 U729 ( .A1(n855), .A2(\REGISTERS[3][21] ), .B1(n15), .B2(
        \REGISTERS[22][21] ), .ZN(n634) );
  AOI22_X1 U730 ( .A1(n857), .A2(\REGISTERS[12][21] ), .B1(n5), .B2(
        \REGISTERS[31][21] ), .ZN(n633) );
  AOI22_X1 U731 ( .A1(n858), .A2(\REGISTERS[29][21] ), .B1(n17), .B2(
        \REGISTERS[20][21] ), .ZN(n632) );
  AOI22_X1 U732 ( .A1(n856), .A2(\REGISTERS[28][21] ), .B1(n9), .B2(
        \REGISTERS[9][21] ), .ZN(n631) );
  NAND4_X1 U733 ( .A1(n634), .A2(n633), .A3(n632), .A4(n631), .ZN(n650) );
  AOI22_X1 U734 ( .A1(n20), .A2(\REGISTERS[8][21] ), .B1(n4), .B2(
        \REGISTERS[27][21] ), .ZN(n638) );
  AOI22_X1 U735 ( .A1(n870), .A2(\REGISTERS[21][21] ), .B1(n18), .B2(
        \REGISTERS[14][21] ), .ZN(n637) );
  AOI22_X1 U736 ( .A1(n847), .A2(\REGISTERS[19][21] ), .B1(n24), .B2(
        \REGISTERS[5][21] ), .ZN(n636) );
  AOI22_X1 U737 ( .A1(n26), .A2(\REGISTERS[7][21] ), .B1(n25), .B2(
        \REGISTERS[15][21] ), .ZN(n635) );
  NAND4_X1 U738 ( .A1(n638), .A2(n637), .A3(n636), .A4(n635), .ZN(n649) );
  AOI22_X1 U739 ( .A1(n882), .A2(\REGISTERS[25][21] ), .B1(n3), .B2(
        \REGISTERS[2][21] ), .ZN(n642) );
  AOI22_X1 U740 ( .A1(n880), .A2(\REGISTERS[30][21] ), .B1(n8), .B2(
        \REGISTERS[1][21] ), .ZN(n641) );
  AOI22_X1 U741 ( .A1(n884), .A2(\REGISTERS[13][21] ), .B1(n10), .B2(
        \REGISTERS[17][21] ), .ZN(n640) );
  AOI22_X1 U742 ( .A1(n841), .A2(\REGISTERS[0][21] ), .B1(n19), .B2(
        \REGISTERS[4][21] ), .ZN(n639) );
  NAND4_X1 U743 ( .A1(n642), .A2(n641), .A3(n640), .A4(n639), .ZN(n648) );
  AOI22_X1 U744 ( .A1(n883), .A2(\REGISTERS[10][21] ), .B1(n6), .B2(
        \REGISTERS[24][21] ), .ZN(n646) );
  AOI22_X1 U745 ( .A1(n16), .A2(\REGISTERS[6][21] ), .B1(n21), .B2(
        \REGISTERS[18][21] ), .ZN(n645) );
  AOI22_X1 U746 ( .A1(n879), .A2(\REGISTERS[26][21] ), .B1(n2), .B2(
        \REGISTERS[23][21] ), .ZN(n644) );
  AOI22_X1 U747 ( .A1(n881), .A2(\REGISTERS[11][21] ), .B1(n23), .B2(
        \REGISTERS[16][21] ), .ZN(n643) );
  NAND4_X1 U748 ( .A1(n646), .A2(n645), .A3(n644), .A4(n643), .ZN(n647) );
  NOR4_X1 U749 ( .A1(n650), .A2(n649), .A3(n648), .A4(n647), .ZN(n651) );
  AOI22_X1 U750 ( .A1(n33), .A2(n94), .B1(n651), .B2(n36), .ZN(N268) );
  AOI22_X1 U751 ( .A1(n878), .A2(\REGISTERS[7][22] ), .B1(n16), .B2(
        \REGISTERS[6][22] ), .ZN(n655) );
  AOI22_X1 U752 ( .A1(n854), .A2(\REGISTERS[17][22] ), .B1(n4), .B2(
        \REGISTERS[27][22] ), .ZN(n654) );
  AOI22_X1 U753 ( .A1(n6), .A2(\REGISTERS[24][22] ), .B1(n24), .B2(
        \REGISTERS[5][22] ), .ZN(n653) );
  AOI22_X1 U754 ( .A1(n857), .A2(\REGISTERS[12][22] ), .B1(n845), .B2(
        \REGISTERS[31][22] ), .ZN(n652) );
  NAND4_X1 U755 ( .A1(n655), .A2(n654), .A3(n653), .A4(n652), .ZN(n671) );
  AOI22_X1 U756 ( .A1(n879), .A2(\REGISTERS[26][22] ), .B1(n32), .B2(
        \REGISTERS[13][22] ), .ZN(n659) );
  AOI22_X1 U757 ( .A1(n866), .A2(\REGISTERS[14][22] ), .B1(n11), .B2(
        \REGISTERS[3][22] ), .ZN(n658) );
  AOI22_X1 U758 ( .A1(n22), .A2(\REGISTERS[21][22] ), .B1(n21), .B2(
        \REGISTERS[18][22] ), .ZN(n657) );
  AOI22_X1 U759 ( .A1(n842), .A2(\REGISTERS[23][22] ), .B1(n19), .B2(
        \REGISTERS[4][22] ), .ZN(n656) );
  NAND4_X1 U760 ( .A1(n659), .A2(n658), .A3(n657), .A4(n656), .ZN(n670) );
  AOI22_X1 U761 ( .A1(n843), .A2(\REGISTERS[2][22] ), .B1(n29), .B2(
        \REGISTERS[11][22] ), .ZN(n663) );
  AOI22_X1 U762 ( .A1(n882), .A2(\REGISTERS[25][22] ), .B1(n31), .B2(
        \REGISTERS[10][22] ), .ZN(n662) );
  AOI22_X1 U763 ( .A1(n880), .A2(\REGISTERS[30][22] ), .B1(n25), .B2(
        \REGISTERS[15][22] ), .ZN(n661) );
  AOI22_X1 U764 ( .A1(n868), .A2(\REGISTERS[8][22] ), .B1(n17), .B2(
        \REGISTERS[20][22] ), .ZN(n660) );
  NAND4_X1 U765 ( .A1(n663), .A2(n662), .A3(n661), .A4(n660), .ZN(n669) );
  AOI22_X1 U766 ( .A1(n858), .A2(\REGISTERS[29][22] ), .B1(n7), .B2(
        \REGISTERS[19][22] ), .ZN(n667) );
  AOI22_X1 U767 ( .A1(n871), .A2(\REGISTERS[16][22] ), .B1(n853), .B2(
        \REGISTERS[9][22] ), .ZN(n666) );
  AOI22_X1 U768 ( .A1(n841), .A2(\REGISTERS[0][22] ), .B1(n859), .B2(
        \REGISTERS[22][22] ), .ZN(n665) );
  AOI22_X1 U769 ( .A1(n856), .A2(\REGISTERS[28][22] ), .B1(n848), .B2(
        \REGISTERS[1][22] ), .ZN(n664) );
  NAND4_X1 U770 ( .A1(n667), .A2(n666), .A3(n665), .A4(n664), .ZN(n668) );
  NOR4_X1 U771 ( .A1(n671), .A2(n670), .A3(n669), .A4(n668), .ZN(n672) );
  AOI22_X1 U772 ( .A1(n33), .A2(n2672), .B1(n672), .B2(n36), .ZN(N269) );
  AOI22_X1 U773 ( .A1(n18), .A2(\REGISTERS[14][23] ), .B1(n24), .B2(
        \REGISTERS[5][23] ), .ZN(n676) );
  AOI22_X1 U774 ( .A1(n878), .A2(\REGISTERS[7][23] ), .B1(n27), .B2(
        \REGISTERS[26][23] ), .ZN(n675) );
  AOI22_X1 U775 ( .A1(n882), .A2(\REGISTERS[25][23] ), .B1(n7), .B2(
        \REGISTERS[19][23] ), .ZN(n674) );
  AOI22_X1 U776 ( .A1(n841), .A2(\REGISTERS[0][23] ), .B1(n17), .B2(
        \REGISTERS[20][23] ), .ZN(n673) );
  NAND4_X1 U777 ( .A1(n676), .A2(n675), .A3(n674), .A4(n673), .ZN(n692) );
  AOI22_X1 U778 ( .A1(n846), .A2(\REGISTERS[24][23] ), .B1(n853), .B2(
        \REGISTERS[9][23] ), .ZN(n680) );
  AOI22_X1 U779 ( .A1(n20), .A2(\REGISTERS[8][23] ), .B1(n845), .B2(
        \REGISTERS[31][23] ), .ZN(n679) );
  AOI22_X1 U780 ( .A1(n8), .A2(\REGISTERS[1][23] ), .B1(n21), .B2(
        \REGISTERS[18][23] ), .ZN(n678) );
  AOI22_X1 U781 ( .A1(n844), .A2(\REGISTERS[27][23] ), .B1(n11), .B2(
        \REGISTERS[3][23] ), .ZN(n677) );
  NAND4_X1 U782 ( .A1(n680), .A2(n679), .A3(n678), .A4(n677), .ZN(n691) );
  AOI22_X1 U783 ( .A1(n842), .A2(\REGISTERS[23][23] ), .B1(n871), .B2(
        \REGISTERS[16][23] ), .ZN(n684) );
  AOI22_X1 U784 ( .A1(n856), .A2(\REGISTERS[28][23] ), .B1(n25), .B2(
        \REGISTERS[15][23] ), .ZN(n683) );
  AOI22_X1 U785 ( .A1(n881), .A2(\REGISTERS[11][23] ), .B1(n859), .B2(
        \REGISTERS[22][23] ), .ZN(n682) );
  AOI22_X1 U786 ( .A1(n858), .A2(\REGISTERS[29][23] ), .B1(n19), .B2(
        \REGISTERS[4][23] ), .ZN(n681) );
  NAND4_X1 U787 ( .A1(n684), .A2(n683), .A3(n682), .A4(n681), .ZN(n690) );
  AOI22_X1 U788 ( .A1(n860), .A2(\REGISTERS[6][23] ), .B1(n13), .B2(
        \REGISTERS[12][23] ), .ZN(n688) );
  AOI22_X1 U789 ( .A1(n10), .A2(\REGISTERS[17][23] ), .B1(n3), .B2(
        \REGISTERS[2][23] ), .ZN(n687) );
  AOI22_X1 U790 ( .A1(n880), .A2(\REGISTERS[30][23] ), .B1(n31), .B2(
        \REGISTERS[10][23] ), .ZN(n686) );
  AOI22_X1 U791 ( .A1(n884), .A2(\REGISTERS[13][23] ), .B1(n22), .B2(
        \REGISTERS[21][23] ), .ZN(n685) );
  NAND4_X1 U792 ( .A1(n688), .A2(n687), .A3(n686), .A4(n685), .ZN(n689) );
  NOR4_X1 U793 ( .A1(n692), .A2(n691), .A3(n690), .A4(n689), .ZN(n693) );
  AOI22_X1 U794 ( .A1(n33), .A2(n90), .B1(n693), .B2(n36), .ZN(N270) );
  AOI22_X1 U795 ( .A1(n868), .A2(\REGISTERS[8][24] ), .B1(n3), .B2(
        \REGISTERS[2][24] ), .ZN(n697) );
  AOI22_X1 U796 ( .A1(n882), .A2(\REGISTERS[25][24] ), .B1(n18), .B2(
        \REGISTERS[14][24] ), .ZN(n696) );
  AOI22_X1 U797 ( .A1(n854), .A2(\REGISTERS[17][24] ), .B1(n4), .B2(
        \REGISTERS[27][24] ), .ZN(n695) );
  AOI22_X1 U798 ( .A1(n880), .A2(\REGISTERS[30][24] ), .B1(n27), .B2(
        \REGISTERS[26][24] ), .ZN(n694) );
  NAND4_X1 U799 ( .A1(n697), .A2(n696), .A3(n695), .A4(n694), .ZN(n713) );
  AOI22_X1 U800 ( .A1(n857), .A2(\REGISTERS[12][24] ), .B1(n5), .B2(
        \REGISTERS[31][24] ), .ZN(n701) );
  AOI22_X1 U801 ( .A1(n872), .A2(\REGISTERS[5][24] ), .B1(n871), .B2(
        \REGISTERS[16][24] ), .ZN(n700) );
  AOI22_X1 U802 ( .A1(n26), .A2(\REGISTERS[7][24] ), .B1(n859), .B2(
        \REGISTERS[22][24] ), .ZN(n699) );
  AOI22_X1 U803 ( .A1(n883), .A2(\REGISTERS[10][24] ), .B1(n8), .B2(
        \REGISTERS[1][24] ), .ZN(n698) );
  NAND4_X1 U804 ( .A1(n701), .A2(n700), .A3(n699), .A4(n698), .ZN(n712) );
  AOI22_X1 U805 ( .A1(n870), .A2(\REGISTERS[21][24] ), .B1(n11), .B2(
        \REGISTERS[3][24] ), .ZN(n705) );
  AOI22_X1 U806 ( .A1(n842), .A2(\REGISTERS[23][24] ), .B1(n7), .B2(
        \REGISTERS[19][24] ), .ZN(n704) );
  AOI22_X1 U807 ( .A1(n858), .A2(\REGISTERS[29][24] ), .B1(n21), .B2(
        \REGISTERS[18][24] ), .ZN(n703) );
  AOI22_X1 U808 ( .A1(n881), .A2(\REGISTERS[11][24] ), .B1(n9), .B2(
        \REGISTERS[9][24] ), .ZN(n702) );
  NAND4_X1 U809 ( .A1(n705), .A2(n704), .A3(n703), .A4(n702), .ZN(n711) );
  AOI22_X1 U810 ( .A1(n865), .A2(\REGISTERS[20][24] ), .B1(n6), .B2(
        \REGISTERS[24][24] ), .ZN(n709) );
  AOI22_X1 U811 ( .A1(n877), .A2(\REGISTERS[15][24] ), .B1(n1), .B2(
        \REGISTERS[0][24] ), .ZN(n708) );
  AOI22_X1 U812 ( .A1(n884), .A2(\REGISTERS[13][24] ), .B1(n19), .B2(
        \REGISTERS[4][24] ), .ZN(n707) );
  AOI22_X1 U813 ( .A1(n856), .A2(\REGISTERS[28][24] ), .B1(n16), .B2(
        \REGISTERS[6][24] ), .ZN(n706) );
  NAND4_X1 U814 ( .A1(n709), .A2(n708), .A3(n707), .A4(n706), .ZN(n710) );
  NOR4_X1 U815 ( .A1(n713), .A2(n712), .A3(n711), .A4(n710), .ZN(n714) );
  AOI22_X1 U816 ( .A1(n34), .A2(n88), .B1(n714), .B2(n36), .ZN(N271) );
  AOI22_X1 U817 ( .A1(n2), .A2(\REGISTERS[23][25] ), .B1(n24), .B2(
        \REGISTERS[5][25] ), .ZN(n718) );
  AOI22_X1 U818 ( .A1(n880), .A2(\REGISTERS[30][25] ), .B1(n29), .B2(
        \REGISTERS[11][25] ), .ZN(n717) );
  AOI22_X1 U819 ( .A1(n12), .A2(\REGISTERS[28][25] ), .B1(n20), .B2(
        \REGISTERS[8][25] ), .ZN(n716) );
  AOI22_X1 U820 ( .A1(n25), .A2(\REGISTERS[15][25] ), .B1(n7), .B2(
        \REGISTERS[19][25] ), .ZN(n715) );
  NAND4_X1 U821 ( .A1(n718), .A2(n717), .A3(n716), .A4(n715), .ZN(n734) );
  AOI22_X1 U822 ( .A1(n10), .A2(\REGISTERS[17][25] ), .B1(n21), .B2(
        \REGISTERS[18][25] ), .ZN(n722) );
  AOI22_X1 U823 ( .A1(n879), .A2(\REGISTERS[26][25] ), .B1(n6), .B2(
        \REGISTERS[24][25] ), .ZN(n721) );
  AOI22_X1 U824 ( .A1(n857), .A2(\REGISTERS[12][25] ), .B1(n9), .B2(
        \REGISTERS[9][25] ), .ZN(n720) );
  AOI22_X1 U825 ( .A1(n1), .A2(\REGISTERS[0][25] ), .B1(n5), .B2(
        \REGISTERS[31][25] ), .ZN(n719) );
  NAND4_X1 U826 ( .A1(n722), .A2(n721), .A3(n720), .A4(n719), .ZN(n733) );
  AOI22_X1 U827 ( .A1(n866), .A2(\REGISTERS[14][25] ), .B1(n4), .B2(
        \REGISTERS[27][25] ), .ZN(n726) );
  AOI22_X1 U828 ( .A1(n882), .A2(\REGISTERS[25][25] ), .B1(n11), .B2(
        \REGISTERS[3][25] ), .ZN(n725) );
  AOI22_X1 U829 ( .A1(n883), .A2(\REGISTERS[10][25] ), .B1(n19), .B2(
        \REGISTERS[4][25] ), .ZN(n724) );
  AOI22_X1 U830 ( .A1(n843), .A2(\REGISTERS[2][25] ), .B1(n859), .B2(
        \REGISTERS[22][25] ), .ZN(n723) );
  NAND4_X1 U831 ( .A1(n726), .A2(n725), .A3(n724), .A4(n723), .ZN(n732) );
  AOI22_X1 U832 ( .A1(n858), .A2(\REGISTERS[29][25] ), .B1(n17), .B2(
        \REGISTERS[20][25] ), .ZN(n730) );
  AOI22_X1 U833 ( .A1(n26), .A2(\REGISTERS[7][25] ), .B1(n22), .B2(
        \REGISTERS[21][25] ), .ZN(n729) );
  AOI22_X1 U834 ( .A1(n884), .A2(\REGISTERS[13][25] ), .B1(n16), .B2(
        \REGISTERS[6][25] ), .ZN(n728) );
  AOI22_X1 U835 ( .A1(n848), .A2(\REGISTERS[1][25] ), .B1(n871), .B2(
        \REGISTERS[16][25] ), .ZN(n727) );
  NAND4_X1 U836 ( .A1(n730), .A2(n729), .A3(n728), .A4(n727), .ZN(n731) );
  NOR4_X1 U837 ( .A1(n734), .A2(n733), .A3(n732), .A4(n731), .ZN(n735) );
  AOI22_X1 U838 ( .A1(n34), .A2(n86), .B1(n735), .B2(n35), .ZN(N272) );
  AOI22_X1 U839 ( .A1(n14), .A2(\REGISTERS[29][26] ), .B1(n871), .B2(
        \REGISTERS[16][26] ), .ZN(n739) );
  AOI22_X1 U840 ( .A1(n6), .A2(\REGISTERS[24][26] ), .B1(n859), .B2(
        \REGISTERS[22][26] ), .ZN(n738) );
  AOI22_X1 U841 ( .A1(n856), .A2(\REGISTERS[28][26] ), .B1(n29), .B2(
        \REGISTERS[11][26] ), .ZN(n737) );
  AOI22_X1 U842 ( .A1(n18), .A2(\REGISTERS[14][26] ), .B1(n5), .B2(
        \REGISTERS[31][26] ), .ZN(n736) );
  NAND4_X1 U843 ( .A1(n739), .A2(n738), .A3(n737), .A4(n736), .ZN(n755) );
  AOI22_X1 U844 ( .A1(n8), .A2(\REGISTERS[1][26] ), .B1(n13), .B2(
        \REGISTERS[12][26] ), .ZN(n743) );
  AOI22_X1 U845 ( .A1(n865), .A2(\REGISTERS[20][26] ), .B1(n9), .B2(
        \REGISTERS[9][26] ), .ZN(n742) );
  AOI22_X1 U846 ( .A1(n30), .A2(\REGISTERS[25][26] ), .B1(n3), .B2(
        \REGISTERS[2][26] ), .ZN(n741) );
  AOI22_X1 U847 ( .A1(n32), .A2(\REGISTERS[13][26] ), .B1(n847), .B2(
        \REGISTERS[19][26] ), .ZN(n740) );
  NAND4_X1 U848 ( .A1(n743), .A2(n742), .A3(n741), .A4(n740), .ZN(n754) );
  AOI22_X1 U849 ( .A1(n26), .A2(\REGISTERS[7][26] ), .B1(n11), .B2(
        \REGISTERS[3][26] ), .ZN(n747) );
  AOI22_X1 U850 ( .A1(n842), .A2(\REGISTERS[23][26] ), .B1(n24), .B2(
        \REGISTERS[5][26] ), .ZN(n746) );
  AOI22_X1 U851 ( .A1(n31), .A2(\REGISTERS[10][26] ), .B1(n19), .B2(
        \REGISTERS[4][26] ), .ZN(n745) );
  AOI22_X1 U852 ( .A1(n877), .A2(\REGISTERS[15][26] ), .B1(n4), .B2(
        \REGISTERS[27][26] ), .ZN(n744) );
  NAND4_X1 U853 ( .A1(n747), .A2(n746), .A3(n745), .A4(n744), .ZN(n753) );
  AOI22_X1 U854 ( .A1(n880), .A2(\REGISTERS[30][26] ), .B1(n1), .B2(
        \REGISTERS[0][26] ), .ZN(n751) );
  AOI22_X1 U855 ( .A1(n879), .A2(\REGISTERS[26][26] ), .B1(n16), .B2(
        \REGISTERS[6][26] ), .ZN(n750) );
  AOI22_X1 U856 ( .A1(n22), .A2(\REGISTERS[21][26] ), .B1(n20), .B2(
        \REGISTERS[8][26] ), .ZN(n749) );
  AOI22_X1 U857 ( .A1(n854), .A2(\REGISTERS[17][26] ), .B1(n21), .B2(
        \REGISTERS[18][26] ), .ZN(n748) );
  NAND4_X1 U858 ( .A1(n751), .A2(n750), .A3(n749), .A4(n748), .ZN(n752) );
  NOR4_X1 U859 ( .A1(n755), .A2(n754), .A3(n753), .A4(n752), .ZN(n756) );
  AOI22_X1 U860 ( .A1(n34), .A2(n84), .B1(n756), .B2(n35), .ZN(N273) );
  AOI22_X1 U861 ( .A1(n27), .A2(\REGISTERS[26][27] ), .B1(n8), .B2(
        \REGISTERS[1][27] ), .ZN(n760) );
  AOI22_X1 U862 ( .A1(n26), .A2(\REGISTERS[7][27] ), .B1(n10), .B2(
        \REGISTERS[17][27] ), .ZN(n759) );
  AOI22_X1 U863 ( .A1(n869), .A2(\REGISTERS[18][27] ), .B1(n872), .B2(
        \REGISTERS[5][27] ), .ZN(n758) );
  AOI22_X1 U864 ( .A1(n2), .A2(\REGISTERS[23][27] ), .B1(n843), .B2(
        \REGISTERS[2][27] ), .ZN(n757) );
  NAND4_X1 U865 ( .A1(n760), .A2(n759), .A3(n758), .A4(n757), .ZN(n776) );
  AOI22_X1 U866 ( .A1(n883), .A2(\REGISTERS[10][27] ), .B1(n15), .B2(
        \REGISTERS[22][27] ), .ZN(n764) );
  AOI22_X1 U867 ( .A1(n847), .A2(\REGISTERS[19][27] ), .B1(n857), .B2(
        \REGISTERS[12][27] ), .ZN(n763) );
  AOI22_X1 U868 ( .A1(n858), .A2(\REGISTERS[29][27] ), .B1(n881), .B2(
        \REGISTERS[11][27] ), .ZN(n762) );
  AOI22_X1 U869 ( .A1(n846), .A2(\REGISTERS[24][27] ), .B1(n9), .B2(
        \REGISTERS[9][27] ), .ZN(n761) );
  NAND4_X1 U870 ( .A1(n764), .A2(n763), .A3(n762), .A4(n761), .ZN(n775) );
  AOI22_X1 U871 ( .A1(n884), .A2(\REGISTERS[13][27] ), .B1(n17), .B2(
        \REGISTERS[20][27] ), .ZN(n768) );
  AOI22_X1 U872 ( .A1(n855), .A2(\REGISTERS[3][27] ), .B1(n5), .B2(
        \REGISTERS[31][27] ), .ZN(n767) );
  AOI22_X1 U873 ( .A1(n12), .A2(\REGISTERS[28][27] ), .B1(n25), .B2(
        \REGISTERS[15][27] ), .ZN(n766) );
  AOI22_X1 U874 ( .A1(n28), .A2(\REGISTERS[30][27] ), .B1(n18), .B2(
        \REGISTERS[14][27] ), .ZN(n765) );
  NAND4_X1 U875 ( .A1(n768), .A2(n767), .A3(n766), .A4(n765), .ZN(n774) );
  AOI22_X1 U876 ( .A1(n16), .A2(\REGISTERS[6][27] ), .B1(n4), .B2(
        \REGISTERS[27][27] ), .ZN(n772) );
  AOI22_X1 U877 ( .A1(n867), .A2(\REGISTERS[4][27] ), .B1(n23), .B2(
        \REGISTERS[16][27] ), .ZN(n771) );
  AOI22_X1 U878 ( .A1(n882), .A2(\REGISTERS[25][27] ), .B1(n1), .B2(
        \REGISTERS[0][27] ), .ZN(n770) );
  AOI22_X1 U879 ( .A1(n870), .A2(\REGISTERS[21][27] ), .B1(n20), .B2(
        \REGISTERS[8][27] ), .ZN(n769) );
  NAND4_X1 U880 ( .A1(n772), .A2(n771), .A3(n770), .A4(n769), .ZN(n773) );
  NOR4_X1 U881 ( .A1(n776), .A2(n775), .A3(n774), .A4(n773), .ZN(n777) );
  AOI22_X1 U882 ( .A1(n34), .A2(n2657), .B1(n777), .B2(n35), .ZN(N274) );
  AOI22_X1 U883 ( .A1(n32), .A2(\REGISTERS[13][28] ), .B1(n869), .B2(
        \REGISTERS[18][28] ), .ZN(n781) );
  AOI22_X1 U884 ( .A1(n841), .A2(\REGISTERS[0][28] ), .B1(n871), .B2(
        \REGISTERS[16][28] ), .ZN(n780) );
  AOI22_X1 U885 ( .A1(n6), .A2(\REGISTERS[24][28] ), .B1(n859), .B2(
        \REGISTERS[22][28] ), .ZN(n779) );
  AOI22_X1 U886 ( .A1(n4), .A2(\REGISTERS[27][28] ), .B1(n17), .B2(
        \REGISTERS[20][28] ), .ZN(n778) );
  NAND4_X1 U887 ( .A1(n781), .A2(n780), .A3(n779), .A4(n778), .ZN(n797) );
  AOI22_X1 U888 ( .A1(n22), .A2(\REGISTERS[21][28] ), .B1(n19), .B2(
        \REGISTERS[4][28] ), .ZN(n785) );
  AOI22_X1 U889 ( .A1(n860), .A2(\REGISTERS[6][28] ), .B1(n5), .B2(
        \REGISTERS[31][28] ), .ZN(n784) );
  AOI22_X1 U890 ( .A1(n31), .A2(\REGISTERS[10][28] ), .B1(n20), .B2(
        \REGISTERS[8][28] ), .ZN(n783) );
  AOI22_X1 U891 ( .A1(n25), .A2(\REGISTERS[15][28] ), .B1(n13), .B2(
        \REGISTERS[12][28] ), .ZN(n782) );
  NAND4_X1 U892 ( .A1(n785), .A2(n784), .A3(n783), .A4(n782), .ZN(n796) );
  AOI22_X1 U893 ( .A1(n26), .A2(\REGISTERS[7][28] ), .B1(n9), .B2(
        \REGISTERS[9][28] ), .ZN(n789) );
  AOI22_X1 U894 ( .A1(n848), .A2(\REGISTERS[1][28] ), .B1(n3), .B2(
        \REGISTERS[2][28] ), .ZN(n788) );
  AOI22_X1 U895 ( .A1(n866), .A2(\REGISTERS[14][28] ), .B1(n2), .B2(
        \REGISTERS[23][28] ), .ZN(n787) );
  AOI22_X1 U896 ( .A1(n14), .A2(\REGISTERS[29][28] ), .B1(n7), .B2(
        \REGISTERS[19][28] ), .ZN(n786) );
  NAND4_X1 U897 ( .A1(n789), .A2(n788), .A3(n787), .A4(n786), .ZN(n795) );
  AOI22_X1 U898 ( .A1(n880), .A2(\REGISTERS[30][28] ), .B1(n11), .B2(
        \REGISTERS[3][28] ), .ZN(n793) );
  AOI22_X1 U899 ( .A1(n856), .A2(\REGISTERS[28][28] ), .B1(n29), .B2(
        \REGISTERS[11][28] ), .ZN(n792) );
  AOI22_X1 U900 ( .A1(n10), .A2(\REGISTERS[17][28] ), .B1(n24), .B2(
        \REGISTERS[5][28] ), .ZN(n791) );
  AOI22_X1 U901 ( .A1(n879), .A2(\REGISTERS[26][28] ), .B1(n30), .B2(
        \REGISTERS[25][28] ), .ZN(n790) );
  NAND4_X1 U902 ( .A1(n793), .A2(n792), .A3(n791), .A4(n790), .ZN(n794) );
  NOR4_X1 U903 ( .A1(n797), .A2(n796), .A3(n795), .A4(n794), .ZN(n798) );
  AOI22_X1 U905 ( .A1(n846), .A2(\REGISTERS[24][29] ), .B1(n24), .B2(
        \REGISTERS[5][29] ), .ZN(n802) );
  AOI22_X1 U906 ( .A1(n30), .A2(\REGISTERS[25][29] ), .B1(n8), .B2(
        \REGISTERS[1][29] ), .ZN(n801) );
  AOI22_X1 U907 ( .A1(n854), .A2(\REGISTERS[17][29] ), .B1(n23), .B2(
        \REGISTERS[16][29] ), .ZN(n800) );
  AOI22_X1 U908 ( .A1(n20), .A2(\REGISTERS[8][29] ), .B1(n9), .B2(
        \REGISTERS[9][29] ), .ZN(n799) );
  NAND4_X1 U909 ( .A1(n802), .A2(n801), .A3(n800), .A4(n799), .ZN(n818) );
  AOI22_X1 U910 ( .A1(n877), .A2(\REGISTERS[15][29] ), .B1(n1), .B2(
        \REGISTERS[0][29] ), .ZN(n806) );
  AOI22_X1 U911 ( .A1(n12), .A2(\REGISTERS[28][29] ), .B1(n881), .B2(
        \REGISTERS[11][29] ), .ZN(n805) );
  AOI22_X1 U912 ( .A1(n16), .A2(\REGISTERS[6][29] ), .B1(n13), .B2(
        \REGISTERS[12][29] ), .ZN(n804) );
  AOI22_X1 U913 ( .A1(n847), .A2(\REGISTERS[19][29] ), .B1(n19), .B2(
        \REGISTERS[4][29] ), .ZN(n803) );
  NAND4_X1 U914 ( .A1(n806), .A2(n805), .A3(n804), .A4(n803), .ZN(n817) );
  AOI22_X1 U915 ( .A1(n883), .A2(\REGISTERS[10][29] ), .B1(n15), .B2(
        \REGISTERS[22][29] ), .ZN(n810) );
  AOI22_X1 U916 ( .A1(n26), .A2(\REGISTERS[7][29] ), .B1(n22), .B2(
        \REGISTERS[21][29] ), .ZN(n809) );
  AOI22_X1 U917 ( .A1(n884), .A2(\REGISTERS[13][29] ), .B1(n11), .B2(
        \REGISTERS[3][29] ), .ZN(n808) );
  AOI22_X1 U918 ( .A1(n28), .A2(\REGISTERS[30][29] ), .B1(n21), .B2(
        \REGISTERS[18][29] ), .ZN(n807) );
  NAND4_X1 U919 ( .A1(n810), .A2(n809), .A3(n808), .A4(n807), .ZN(n816) );
  AOI22_X1 U920 ( .A1(n27), .A2(\REGISTERS[26][29] ), .B1(n14), .B2(
        \REGISTERS[29][29] ), .ZN(n814) );
  AOI22_X1 U921 ( .A1(n18), .A2(\REGISTERS[14][29] ), .B1(n5), .B2(
        \REGISTERS[31][29] ), .ZN(n813) );
  AOI22_X1 U922 ( .A1(n844), .A2(\REGISTERS[27][29] ), .B1(n843), .B2(
        \REGISTERS[2][29] ), .ZN(n812) );
  AOI22_X1 U923 ( .A1(n842), .A2(\REGISTERS[23][29] ), .B1(n865), .B2(
        \REGISTERS[20][29] ), .ZN(n811) );
  NAND4_X1 U924 ( .A1(n814), .A2(n813), .A3(n812), .A4(n811), .ZN(n815) );
  NOR4_X1 U925 ( .A1(n818), .A2(n817), .A3(n816), .A4(n815), .ZN(n819) );
  AOI22_X1 U926 ( .A1(n34), .A2(n2665), .B1(n819), .B2(n35), .ZN(N276) );
  AOI22_X1 U927 ( .A1(n880), .A2(\REGISTERS[30][30] ), .B1(n857), .B2(
        \REGISTERS[12][30] ), .ZN(n823) );
  AOI22_X1 U928 ( .A1(n860), .A2(\REGISTERS[6][30] ), .B1(n872), .B2(
        \REGISTERS[5][30] ), .ZN(n822) );
  AOI22_X1 U929 ( .A1(n32), .A2(\REGISTERS[13][30] ), .B1(n8), .B2(
        \REGISTERS[1][30] ), .ZN(n821) );
  AOI22_X1 U930 ( .A1(n31), .A2(\REGISTERS[10][30] ), .B1(n859), .B2(
        \REGISTERS[22][30] ), .ZN(n820) );
  NAND4_X1 U931 ( .A1(n823), .A2(n822), .A3(n821), .A4(n820), .ZN(n839) );
  AOI22_X1 U932 ( .A1(n2), .A2(\REGISTERS[23][30] ), .B1(n5), .B2(
        \REGISTERS[31][30] ), .ZN(n827) );
  AOI22_X1 U933 ( .A1(n879), .A2(\REGISTERS[26][30] ), .B1(n871), .B2(
        \REGISTERS[16][30] ), .ZN(n826) );
  AOI22_X1 U934 ( .A1(n26), .A2(\REGISTERS[7][30] ), .B1(n19), .B2(
        \REGISTERS[4][30] ), .ZN(n825) );
  AOI22_X1 U935 ( .A1(n858), .A2(\REGISTERS[29][30] ), .B1(n7), .B2(
        \REGISTERS[19][30] ), .ZN(n824) );
  NAND4_X1 U936 ( .A1(n827), .A2(n826), .A3(n825), .A4(n824), .ZN(n838) );
  AOI22_X1 U937 ( .A1(n17), .A2(\REGISTERS[20][30] ), .B1(n6), .B2(
        \REGISTERS[24][30] ), .ZN(n831) );
  AOI22_X1 U938 ( .A1(n882), .A2(\REGISTERS[25][30] ), .B1(n25), .B2(
        \REGISTERS[15][30] ), .ZN(n830) );
  AOI22_X1 U939 ( .A1(n1), .A2(\REGISTERS[0][30] ), .B1(n869), .B2(
        \REGISTERS[18][30] ), .ZN(n829) );
  AOI22_X1 U940 ( .A1(n870), .A2(\REGISTERS[21][30] ), .B1(n11), .B2(
        \REGISTERS[3][30] ), .ZN(n828) );
  NAND4_X1 U941 ( .A1(n831), .A2(n830), .A3(n829), .A4(n828), .ZN(n837) );
  AOI22_X1 U942 ( .A1(n868), .A2(\REGISTERS[8][30] ), .B1(n29), .B2(
        \REGISTERS[11][30] ), .ZN(n835) );
  AOI22_X1 U943 ( .A1(n866), .A2(\REGISTERS[14][30] ), .B1(n4), .B2(
        \REGISTERS[27][30] ), .ZN(n834) );
  AOI22_X1 U944 ( .A1(n856), .A2(\REGISTERS[28][30] ), .B1(n10), .B2(
        \REGISTERS[17][30] ), .ZN(n833) );
  AOI22_X1 U945 ( .A1(n843), .A2(\REGISTERS[2][30] ), .B1(n9), .B2(
        \REGISTERS[9][30] ), .ZN(n832) );
  NAND4_X1 U946 ( .A1(n835), .A2(n834), .A3(n833), .A4(n832), .ZN(n836) );
  NOR4_X1 U947 ( .A1(n839), .A2(n838), .A3(n837), .A4(n836), .ZN(n840) );
  AOI22_X1 U948 ( .A1(n34), .A2(n2664), .B1(n840), .B2(n35), .ZN(N277) );
  AOI22_X1 U949 ( .A1(n2), .A2(\REGISTERS[23][31] ), .B1(n1), .B2(
        \REGISTERS[0][31] ), .ZN(n852) );
  AOI22_X1 U950 ( .A1(n844), .A2(\REGISTERS[27][31] ), .B1(n3), .B2(
        \REGISTERS[2][31] ), .ZN(n851) );
  AOI22_X1 U951 ( .A1(n846), .A2(\REGISTERS[24][31] ), .B1(n5), .B2(
        \REGISTERS[31][31] ), .ZN(n850) );
  AOI22_X1 U952 ( .A1(n848), .A2(\REGISTERS[1][31] ), .B1(n7), .B2(
        \REGISTERS[19][31] ), .ZN(n849) );
  NAND4_X1 U953 ( .A1(n852), .A2(n851), .A3(n850), .A4(n849), .ZN(n892) );
  AOI22_X1 U954 ( .A1(n10), .A2(\REGISTERS[17][31] ), .B1(n9), .B2(
        \REGISTERS[9][31] ), .ZN(n864) );
  AOI22_X1 U955 ( .A1(n12), .A2(\REGISTERS[28][31] ), .B1(n11), .B2(
        \REGISTERS[3][31] ), .ZN(n863) );
  AOI22_X1 U956 ( .A1(n14), .A2(\REGISTERS[29][31] ), .B1(n13), .B2(
        \REGISTERS[12][31] ), .ZN(n862) );
  AOI22_X1 U957 ( .A1(n16), .A2(\REGISTERS[6][31] ), .B1(n15), .B2(
        \REGISTERS[22][31] ), .ZN(n861) );
  NAND4_X1 U958 ( .A1(n864), .A2(n863), .A3(n862), .A4(n861), .ZN(n891) );
  AOI22_X1 U959 ( .A1(n866), .A2(\REGISTERS[14][31] ), .B1(n17), .B2(
        \REGISTERS[20][31] ), .ZN(n876) );
  AOI22_X1 U960 ( .A1(n20), .A2(\REGISTERS[8][31] ), .B1(n867), .B2(
        \REGISTERS[4][31] ), .ZN(n875) );
  AOI22_X1 U961 ( .A1(n870), .A2(\REGISTERS[21][31] ), .B1(n21), .B2(
        \REGISTERS[18][31] ), .ZN(n874) );
  AOI22_X1 U962 ( .A1(n872), .A2(\REGISTERS[5][31] ), .B1(n23), .B2(
        \REGISTERS[16][31] ), .ZN(n873) );
  NAND4_X1 U963 ( .A1(n876), .A2(n875), .A3(n874), .A4(n873), .ZN(n890) );
  AOI22_X1 U964 ( .A1(n26), .A2(\REGISTERS[7][31] ), .B1(n25), .B2(
        \REGISTERS[15][31] ), .ZN(n888) );
  AOI22_X1 U965 ( .A1(n28), .A2(\REGISTERS[30][31] ), .B1(n27), .B2(
        \REGISTERS[26][31] ), .ZN(n887) );
  AOI22_X1 U966 ( .A1(n30), .A2(\REGISTERS[25][31] ), .B1(n29), .B2(
        \REGISTERS[11][31] ), .ZN(n886) );
  AOI22_X1 U967 ( .A1(n32), .A2(\REGISTERS[13][31] ), .B1(n31), .B2(
        \REGISTERS[10][31] ), .ZN(n885) );
  NAND4_X1 U968 ( .A1(n888), .A2(n887), .A3(n886), .A4(n885), .ZN(n889) );
  NOR4_X1 U969 ( .A1(n892), .A2(n891), .A3(n890), .A4(n889), .ZN(n893) );
  AOI22_X1 U970 ( .A1(n34), .A2(n2671), .B1(n893), .B2(n35), .ZN(N278) );
  OAI221_X1 U971 ( .B1(ADD_WR[4]), .B2(n913), .C1(n895), .C2(ADD_RD2[4]), .A(
        WR), .ZN(n904) );
  AOI22_X1 U972 ( .A1(n898), .A2(ADD_RD2[3]), .B1(ADD_RD2[1]), .B2(n897), .ZN(
        n896) );
  OAI221_X1 U973 ( .B1(n898), .B2(ADD_RD2[3]), .C1(n897), .C2(ADD_RD2[1]), .A(
        n896), .ZN(n903) );
  AOI22_X1 U974 ( .A1(n901), .A2(ADD_RD2[2]), .B1(n900), .B2(ADD_RD2[0]), .ZN(
        n899) );
  OAI221_X1 U975 ( .B1(n901), .B2(ADD_RD2[2]), .C1(n900), .C2(ADD_RD2[0]), .A(
        n899), .ZN(n902) );
  INV_X1 U976 ( .A(ADD_RD2[2]), .ZN(n905) );
  NAND2_X1 U977 ( .A1(ADD_RD2[1]), .A2(n905), .ZN(n928) );
  INV_X1 U978 ( .A(ADD_RD2[3]), .ZN(n907) );
  NAND3_X1 U979 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[0]), .A3(n907), .ZN(n925) );
  NOR2_X1 U980 ( .A1(n928), .A2(n925), .ZN(n1604) );
  INV_X1 U981 ( .A(ADD_RD2[1]), .ZN(n906) );
  NAND2_X1 U982 ( .A1(n905), .A2(n906), .ZN(n931) );
  NAND3_X1 U983 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n913), .ZN(n920) );
  NOR2_X1 U984 ( .A1(n931), .A2(n920), .ZN(n1580) );
  AOI22_X1 U985 ( .A1(\REGISTERS[19][0] ), .A2(n58), .B1(\REGISTERS[9][0] ), 
        .B2(n42), .ZN(n912) );
  NAND2_X1 U986 ( .A1(ADD_RD2[2]), .A2(ADD_RD2[1]), .ZN(n926) );
  NOR2_X1 U987 ( .A1(n925), .A2(n926), .ZN(n1590) );
  NAND2_X1 U988 ( .A1(ADD_RD2[2]), .A2(n906), .ZN(n934) );
  NOR2_X1 U989 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .ZN(n908) );
  NAND2_X1 U990 ( .A1(ADD_RD2[4]), .A2(n908), .ZN(n930) );
  NOR2_X1 U991 ( .A1(n934), .A2(n930), .ZN(n1616) );
  AOI22_X1 U992 ( .A1(\REGISTERS[23][0] ), .A2(n48), .B1(\REGISTERS[20][0] ), 
        .B2(n66), .ZN(n911) );
  INV_X1 U993 ( .A(ADD_RD2[0]), .ZN(n914) );
  NAND3_X1 U994 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .A3(n914), .ZN(n932) );
  NOR2_X1 U995 ( .A1(n926), .A2(n932), .ZN(n1615) );
  NAND3_X1 U996 ( .A1(ADD_RD2[0]), .A2(n913), .A3(n907), .ZN(n933) );
  NOR2_X1 U997 ( .A1(n928), .A2(n933), .ZN(n1592) );
  AOI22_X1 U998 ( .A1(\REGISTERS[30][0] ), .A2(n65), .B1(\REGISTERS[3][0] ), 
        .B2(n50), .ZN(n910) );
  NAND2_X1 U999 ( .A1(n908), .A2(n913), .ZN(n929) );
  NOR2_X1 U1000 ( .A1(n931), .A2(n929), .ZN(n1614) );
  NAND3_X1 U1001 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(ADD_RD2[3]), .ZN(n919) );
  NOR2_X1 U1002 ( .A1(n926), .A2(n919), .ZN(n1600) );
  AOI22_X1 U1003 ( .A1(\REGISTERS[0][0] ), .A2(n64), .B1(\REGISTERS[31][0] ), 
        .B2(n54), .ZN(n909) );
  NAND4_X1 U1004 ( .A1(n912), .A2(n911), .A3(n910), .A4(n909), .ZN(n942) );
  NOR2_X1 U1005 ( .A1(n928), .A2(n932), .ZN(n1603) );
  NAND3_X1 U1006 ( .A1(ADD_RD2[3]), .A2(n914), .A3(n913), .ZN(n927) );
  NOR2_X1 U1007 ( .A1(n928), .A2(n927), .ZN(n1579) );
  AOI22_X1 U1008 ( .A1(\REGISTERS[26][0] ), .A2(n57), .B1(\REGISTERS[10][0] ), 
        .B2(n41), .ZN(n918) );
  NOR2_X1 U1009 ( .A1(n926), .A2(n929), .ZN(n1617) );
  NOR2_X1 U1010 ( .A1(n926), .A2(n927), .ZN(n1582) );
  AOI22_X1 U1011 ( .A1(\REGISTERS[6][0] ), .A2(n67), .B1(\REGISTERS[14][0] ), 
        .B2(n44), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(n920), .A2(n934), .ZN(n1587) );
  NOR2_X1 U1013 ( .A1(n934), .A2(n919), .ZN(n1618) );
  AOI22_X1 U1014 ( .A1(\REGISTERS[13][0] ), .A2(n1587), .B1(\REGISTERS[29][0] ), .B2(n68), .ZN(n916) );
  NOR2_X1 U1015 ( .A1(n931), .A2(n933), .ZN(n1577) );
  NOR2_X1 U1016 ( .A1(n920), .A2(n928), .ZN(n1591) );
  AOI22_X1 U1017 ( .A1(\REGISTERS[1][0] ), .A2(n39), .B1(\REGISTERS[11][0] ), 
        .B2(n49), .ZN(n915) );
  NAND4_X1 U1018 ( .A1(n918), .A2(n917), .A3(n916), .A4(n915), .ZN(n941) );
  NOR2_X1 U1019 ( .A1(n931), .A2(n919), .ZN(n1611) );
  NOR2_X1 U1020 ( .A1(n928), .A2(n919), .ZN(n1578) );
  AOI22_X1 U1021 ( .A1(\REGISTERS[25][0] ), .A2(n1611), .B1(\REGISTERS[27][0] ), .B2(n40), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n926), .ZN(n1601) );
  NOR2_X1 U1023 ( .A1(n931), .A2(n932), .ZN(n1589) );
  AOI22_X1 U1024 ( .A1(\REGISTERS[15][0] ), .A2(n55), .B1(\REGISTERS[24][0] ), 
        .B2(n47), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n933), .ZN(n1581) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n927), .ZN(n1576) );
  AOI22_X1 U1027 ( .A1(\REGISTERS[7][0] ), .A2(n1581), .B1(\REGISTERS[8][0] ), 
        .B2(n38), .ZN(n922) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n925), .ZN(n1594) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n930), .ZN(n1605) );
  AOI22_X1 U1030 ( .A1(\REGISTERS[17][0] ), .A2(n52), .B1(\REGISTERS[18][0] ), 
        .B2(n59), .ZN(n921) );
  NAND4_X1 U1031 ( .A1(n924), .A2(n923), .A3(n922), .A4(n921), .ZN(n940) );
  NOR2_X1 U1032 ( .A1(n925), .A2(n934), .ZN(n1599) );
  NOR2_X1 U1033 ( .A1(n926), .A2(n930), .ZN(n1593) );
  AOI22_X1 U1034 ( .A1(\REGISTERS[21][0] ), .A2(n53), .B1(\REGISTERS[22][0] ), 
        .B2(n51), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n927), .ZN(n1602) );
  NOR2_X1 U1036 ( .A1(n928), .A2(n929), .ZN(n1588) );
  AOI22_X1 U1037 ( .A1(\REGISTERS[12][0] ), .A2(n56), .B1(\REGISTERS[2][0] ), 
        .B2(n46), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(n934), .A2(n929), .ZN(n1575) );
  NOR2_X1 U1039 ( .A1(n931), .A2(n930), .ZN(n1613) );
  AOI22_X1 U1040 ( .A1(\REGISTERS[4][0] ), .A2(n1575), .B1(\REGISTERS[16][0] ), 
        .B2(n63), .ZN(n936) );
  NOR2_X1 U1041 ( .A1(n934), .A2(n932), .ZN(n1606) );
  NOR2_X1 U1042 ( .A1(n934), .A2(n933), .ZN(n1612) );
  AOI22_X1 U1043 ( .A1(\REGISTERS[28][0] ), .A2(n60), .B1(\REGISTERS[5][0] ), 
        .B2(n62), .ZN(n935) );
  NAND4_X1 U1044 ( .A1(n938), .A2(n937), .A3(n936), .A4(n935), .ZN(n939) );
  NOR4_X1 U1045 ( .A1(n942), .A2(n941), .A3(n940), .A4(n939), .ZN(n943) );
  AOI22_X1 U1046 ( .A1(n69), .A2(n2677), .B1(n943), .B2(n72), .ZN(N379) );
  AOI22_X1 U1047 ( .A1(\REGISTERS[3][1] ), .A2(n1592), .B1(\REGISTERS[28][1] ), 
        .B2(n60), .ZN(n947) );
  AOI22_X1 U1048 ( .A1(\REGISTERS[20][1] ), .A2(n1616), .B1(\REGISTERS[13][1] ), .B2(n45), .ZN(n946) );
  AOI22_X1 U1049 ( .A1(\REGISTERS[1][1] ), .A2(n1577), .B1(\REGISTERS[17][1] ), 
        .B2(n52), .ZN(n945) );
  AOI22_X1 U1050 ( .A1(\REGISTERS[18][1] ), .A2(n1605), .B1(\REGISTERS[6][1] ), 
        .B2(n67), .ZN(n944) );
  NAND4_X1 U1051 ( .A1(n947), .A2(n946), .A3(n945), .A4(n944), .ZN(n963) );
  AOI22_X1 U1052 ( .A1(\REGISTERS[12][1] ), .A2(n56), .B1(\REGISTERS[5][1] ), 
        .B2(n62), .ZN(n951) );
  AOI22_X1 U1053 ( .A1(\REGISTERS[24][1] ), .A2(n1589), .B1(\REGISTERS[30][1] ), .B2(n65), .ZN(n950) );
  AOI22_X1 U1054 ( .A1(\REGISTERS[4][1] ), .A2(n37), .B1(\REGISTERS[16][1] ), 
        .B2(n63), .ZN(n949) );
  AOI22_X1 U1055 ( .A1(\REGISTERS[27][1] ), .A2(n1578), .B1(\REGISTERS[0][1] ), 
        .B2(n64), .ZN(n948) );
  NAND4_X1 U1056 ( .A1(n951), .A2(n950), .A3(n949), .A4(n948), .ZN(n962) );
  AOI22_X1 U1057 ( .A1(\REGISTERS[26][1] ), .A2(n57), .B1(\REGISTERS[21][1] ), 
        .B2(n53), .ZN(n955) );
  AOI22_X1 U1058 ( .A1(\REGISTERS[14][1] ), .A2(n1582), .B1(\REGISTERS[11][1] ), .B2(n49), .ZN(n954) );
  AOI22_X1 U1059 ( .A1(\REGISTERS[8][1] ), .A2(n1576), .B1(\REGISTERS[15][1] ), 
        .B2(n55), .ZN(n953) );
  AOI22_X1 U1060 ( .A1(\REGISTERS[25][1] ), .A2(n1611), .B1(\REGISTERS[7][1] ), 
        .B2(n1581), .ZN(n952) );
  NAND4_X1 U1061 ( .A1(n955), .A2(n954), .A3(n953), .A4(n952), .ZN(n961) );
  AOI22_X1 U1062 ( .A1(\REGISTERS[23][1] ), .A2(n1590), .B1(\REGISTERS[19][1] ), .B2(n58), .ZN(n959) );
  AOI22_X1 U1063 ( .A1(\REGISTERS[22][1] ), .A2(n51), .B1(\REGISTERS[2][1] ), 
        .B2(n46), .ZN(n958) );
  AOI22_X1 U1064 ( .A1(\REGISTERS[10][1] ), .A2(n1579), .B1(\REGISTERS[29][1] ), .B2(n68), .ZN(n957) );
  AOI22_X1 U1065 ( .A1(\REGISTERS[9][1] ), .A2(n1580), .B1(\REGISTERS[31][1] ), 
        .B2(n54), .ZN(n956) );
  NAND4_X1 U1066 ( .A1(n959), .A2(n958), .A3(n957), .A4(n956), .ZN(n960) );
  NOR4_X1 U1067 ( .A1(n963), .A2(n962), .A3(n961), .A4(n960), .ZN(n964) );
  AOI22_X1 U1068 ( .A1(n70), .A2(n134), .B1(n964), .B2(n71), .ZN(N380) );
  AOI22_X1 U1069 ( .A1(\REGISTERS[9][2] ), .A2(n42), .B1(\REGISTERS[10][2] ), 
        .B2(n41), .ZN(n968) );
  AOI22_X1 U1070 ( .A1(\REGISTERS[30][2] ), .A2(n65), .B1(\REGISTERS[3][2] ), 
        .B2(n50), .ZN(n967) );
  AOI22_X1 U1071 ( .A1(\REGISTERS[12][2] ), .A2(n1602), .B1(\REGISTERS[6][2] ), 
        .B2(n67), .ZN(n966) );
  AOI22_X1 U1072 ( .A1(\REGISTERS[22][2] ), .A2(n1593), .B1(\REGISTERS[15][2] ), .B2(n55), .ZN(n965) );
  NAND4_X1 U1073 ( .A1(n968), .A2(n967), .A3(n966), .A4(n965), .ZN(n984) );
  AOI22_X1 U1074 ( .A1(\REGISTERS[19][2] ), .A2(n1604), .B1(\REGISTERS[18][2] ), .B2(n59), .ZN(n972) );
  AOI22_X1 U1075 ( .A1(\REGISTERS[21][2] ), .A2(n1599), .B1(\REGISTERS[26][2] ), .B2(n57), .ZN(n971) );
  AOI22_X1 U1076 ( .A1(\REGISTERS[5][2] ), .A2(n62), .B1(\REGISTERS[8][2] ), 
        .B2(n38), .ZN(n970) );
  AOI22_X1 U1077 ( .A1(\REGISTERS[17][2] ), .A2(n1594), .B1(\REGISTERS[14][2] ), .B2(n44), .ZN(n969) );
  NAND4_X1 U1078 ( .A1(n972), .A2(n971), .A3(n970), .A4(n969), .ZN(n983) );
  AOI22_X1 U1079 ( .A1(\REGISTERS[28][2] ), .A2(n1606), .B1(\REGISTERS[7][2] ), 
        .B2(n1581), .ZN(n976) );
  AOI22_X1 U1080 ( .A1(\REGISTERS[16][2] ), .A2(n1613), .B1(\REGISTERS[31][2] ), .B2(n54), .ZN(n975) );
  AOI22_X1 U1081 ( .A1(\REGISTERS[24][2] ), .A2(n47), .B1(\REGISTERS[11][2] ), 
        .B2(n49), .ZN(n974) );
  AOI22_X1 U1082 ( .A1(\REGISTERS[0][2] ), .A2(n1614), .B1(\REGISTERS[2][2] ), 
        .B2(n46), .ZN(n973) );
  NAND4_X1 U1083 ( .A1(n976), .A2(n975), .A3(n974), .A4(n973), .ZN(n982) );
  AOI22_X1 U1084 ( .A1(\REGISTERS[25][2] ), .A2(n1611), .B1(\REGISTERS[4][2] ), 
        .B2(n37), .ZN(n980) );
  AOI22_X1 U1085 ( .A1(\REGISTERS[20][2] ), .A2(n1616), .B1(\REGISTERS[29][2] ), .B2(n68), .ZN(n979) );
  AOI22_X1 U1086 ( .A1(\REGISTERS[1][2] ), .A2(n1577), .B1(\REGISTERS[27][2] ), 
        .B2(n40), .ZN(n978) );
  AOI22_X1 U1087 ( .A1(\REGISTERS[23][2] ), .A2(n48), .B1(\REGISTERS[13][2] ), 
        .B2(n45), .ZN(n977) );
  NAND4_X1 U1088 ( .A1(n980), .A2(n979), .A3(n978), .A4(n977), .ZN(n981) );
  NOR4_X1 U1089 ( .A1(n984), .A2(n983), .A3(n982), .A4(n981), .ZN(n985) );
  AOI22_X1 U1090 ( .A1(n70), .A2(n2669), .B1(n985), .B2(n72), .ZN(N381) );
  AOI22_X1 U1091 ( .A1(\REGISTERS[2][3] ), .A2(n46), .B1(\REGISTERS[12][3] ), 
        .B2(n56), .ZN(n989) );
  AOI22_X1 U1092 ( .A1(\REGISTERS[3][3] ), .A2(n50), .B1(\REGISTERS[8][3] ), 
        .B2(n38), .ZN(n988) );
  AOI22_X1 U1093 ( .A1(\REGISTERS[16][3] ), .A2(n63), .B1(\REGISTERS[31][3] ), 
        .B2(n54), .ZN(n987) );
  AOI22_X1 U1094 ( .A1(\REGISTERS[18][3] ), .A2(n1605), .B1(\REGISTERS[25][3] ), .B2(n61), .ZN(n986) );
  NAND4_X1 U1095 ( .A1(n989), .A2(n988), .A3(n987), .A4(n986), .ZN(n1005) );
  AOI22_X1 U1096 ( .A1(\REGISTERS[20][3] ), .A2(n66), .B1(\REGISTERS[26][3] ), 
        .B2(n57), .ZN(n993) );
  AOI22_X1 U1097 ( .A1(\REGISTERS[27][3] ), .A2(n1578), .B1(\REGISTERS[17][3] ), .B2(n52), .ZN(n992) );
  AOI22_X1 U1098 ( .A1(\REGISTERS[14][3] ), .A2(n44), .B1(\REGISTERS[23][3] ), 
        .B2(n48), .ZN(n991) );
  AOI22_X1 U1099 ( .A1(\REGISTERS[9][3] ), .A2(n1580), .B1(\REGISTERS[28][3] ), 
        .B2(n60), .ZN(n990) );
  NAND4_X1 U1100 ( .A1(n993), .A2(n992), .A3(n991), .A4(n990), .ZN(n1004) );
  AOI22_X1 U1101 ( .A1(\REGISTERS[30][3] ), .A2(n1615), .B1(\REGISTERS[5][3] ), 
        .B2(n62), .ZN(n997) );
  AOI22_X1 U1102 ( .A1(\REGISTERS[0][3] ), .A2(n1614), .B1(\REGISTERS[22][3] ), 
        .B2(n51), .ZN(n996) );
  AOI22_X1 U1103 ( .A1(\REGISTERS[15][3] ), .A2(n55), .B1(\REGISTERS[1][3] ), 
        .B2(n39), .ZN(n995) );
  AOI22_X1 U1104 ( .A1(\REGISTERS[21][3] ), .A2(n53), .B1(\REGISTERS[19][3] ), 
        .B2(n58), .ZN(n994) );
  NAND4_X1 U1105 ( .A1(n997), .A2(n996), .A3(n995), .A4(n994), .ZN(n1003) );
  AOI22_X1 U1106 ( .A1(\REGISTERS[4][3] ), .A2(n1575), .B1(\REGISTERS[7][3] ), 
        .B2(n43), .ZN(n1001) );
  AOI22_X1 U1107 ( .A1(\REGISTERS[10][3] ), .A2(n1579), .B1(\REGISTERS[24][3] ), .B2(n47), .ZN(n1000) );
  AOI22_X1 U1108 ( .A1(\REGISTERS[29][3] ), .A2(n1618), .B1(\REGISTERS[13][3] ), .B2(n45), .ZN(n999) );
  AOI22_X1 U1109 ( .A1(\REGISTERS[11][3] ), .A2(n49), .B1(\REGISTERS[6][3] ), 
        .B2(n67), .ZN(n998) );
  NAND4_X1 U1110 ( .A1(n1001), .A2(n1000), .A3(n999), .A4(n998), .ZN(n1002) );
  NOR4_X1 U1111 ( .A1(n1005), .A2(n1004), .A3(n1003), .A4(n1002), .ZN(n1006)
         );
  AOI22_X1 U1112 ( .A1(n70), .A2(n2670), .B1(n1006), .B2(n71), .ZN(N382) );
  AOI22_X1 U1113 ( .A1(\REGISTERS[0][4] ), .A2(n64), .B1(\REGISTERS[30][4] ), 
        .B2(n65), .ZN(n1010) );
  AOI22_X1 U1114 ( .A1(\REGISTERS[18][4] ), .A2(n1605), .B1(\REGISTERS[9][4] ), 
        .B2(n42), .ZN(n1009) );
  AOI22_X1 U1115 ( .A1(\REGISTERS[3][4] ), .A2(n1592), .B1(\REGISTERS[7][4] ), 
        .B2(n43), .ZN(n1008) );
  AOI22_X1 U1116 ( .A1(\REGISTERS[26][4] ), .A2(n1603), .B1(\REGISTERS[19][4] ), .B2(n58), .ZN(n1007) );
  NAND4_X1 U1117 ( .A1(n1010), .A2(n1009), .A3(n1008), .A4(n1007), .ZN(n1027)
         );
  AOI22_X1 U1118 ( .A1(\REGISTERS[27][4] ), .A2(n40), .B1(\REGISTERS[8][4] ), 
        .B2(n38), .ZN(n1014) );
  AOI22_X1 U1119 ( .A1(\REGISTERS[1][4] ), .A2(n1577), .B1(\REGISTERS[10][4] ), 
        .B2(n41), .ZN(n1013) );
  AOI22_X1 U1120 ( .A1(\REGISTERS[25][4] ), .A2(n61), .B1(\REGISTERS[22][4] ), 
        .B2(n51), .ZN(n1012) );
  AOI22_X1 U1121 ( .A1(\REGISTERS[4][4] ), .A2(n37), .B1(\REGISTERS[20][4] ), 
        .B2(n66), .ZN(n1011) );
  NAND4_X1 U1122 ( .A1(n1014), .A2(n1013), .A3(n1012), .A4(n1011), .ZN(n1026)
         );
  AOI22_X1 U1123 ( .A1(\REGISTERS[28][4] ), .A2(n60), .B1(\REGISTERS[23][4] ), 
        .B2(n48), .ZN(n1018) );
  AOI22_X1 U1124 ( .A1(\REGISTERS[14][4] ), .A2(n1582), .B1(\REGISTERS[5][4] ), 
        .B2(n62), .ZN(n1017) );
  AOI22_X1 U1125 ( .A1(\REGISTERS[16][4] ), .A2(n1613), .B1(\REGISTERS[2][4] ), 
        .B2(n46), .ZN(n1016) );
  AOI22_X1 U1126 ( .A1(\REGISTERS[21][4] ), .A2(n1599), .B1(\REGISTERS[31][4] ), .B2(n54), .ZN(n1015) );
  NAND4_X1 U1127 ( .A1(n1018), .A2(n1017), .A3(n1016), .A4(n1015), .ZN(n1025)
         );
  AOI22_X1 U1128 ( .A1(\REGISTERS[29][4] ), .A2(n1618), .B1(\REGISTERS[24][4] ), .B2(n47), .ZN(n1022) );
  AOI22_X1 U1129 ( .A1(\REGISTERS[13][4] ), .A2(n1587), .B1(\REGISTERS[6][4] ), 
        .B2(n67), .ZN(n1021) );
  AOI22_X1 U1130 ( .A1(\REGISTERS[15][4] ), .A2(n1601), .B1(\REGISTERS[12][4] ), .B2(n56), .ZN(n1020) );
  AOI22_X1 U1131 ( .A1(\REGISTERS[11][4] ), .A2(n49), .B1(\REGISTERS[17][4] ), 
        .B2(n52), .ZN(n1019) );
  NAND4_X1 U1132 ( .A1(n1022), .A2(n1021), .A3(n1020), .A4(n1019), .ZN(n1023)
         );
  NOR4_X1 U1133 ( .A1(n1027), .A2(n1026), .A3(n1025), .A4(n1023), .ZN(n1028)
         );
  AOI22_X1 U1134 ( .A1(n70), .A2(n2676), .B1(n1028), .B2(n72), .ZN(N383) );
  AOI22_X1 U1135 ( .A1(\REGISTERS[25][5] ), .A2(n61), .B1(\REGISTERS[16][5] ), 
        .B2(n63), .ZN(n1032) );
  AOI22_X1 U1136 ( .A1(\REGISTERS[14][5] ), .A2(n1582), .B1(\REGISTERS[12][5] ), .B2(n56), .ZN(n1031) );
  AOI22_X1 U1137 ( .A1(\REGISTERS[30][5] ), .A2(n1615), .B1(\REGISTERS[8][5] ), 
        .B2(n38), .ZN(n1030) );
  AOI22_X1 U1138 ( .A1(\REGISTERS[3][5] ), .A2(n50), .B1(\REGISTERS[0][5] ), 
        .B2(n64), .ZN(n1029) );
  NAND4_X1 U1139 ( .A1(n1032), .A2(n1031), .A3(n1030), .A4(n1029), .ZN(n1048)
         );
  AOI22_X1 U1140 ( .A1(\REGISTERS[20][5] ), .A2(n66), .B1(\REGISTERS[10][5] ), 
        .B2(n41), .ZN(n1036) );
  AOI22_X1 U1141 ( .A1(\REGISTERS[28][5] ), .A2(n1606), .B1(\REGISTERS[18][5] ), .B2(n59), .ZN(n1035) );
  AOI22_X1 U1142 ( .A1(\REGISTERS[17][5] ), .A2(n1594), .B1(\REGISTERS[5][5] ), 
        .B2(n62), .ZN(n1034) );
  AOI22_X1 U1143 ( .A1(\REGISTERS[13][5] ), .A2(n45), .B1(\REGISTERS[31][5] ), 
        .B2(n54), .ZN(n1033) );
  NAND4_X1 U1144 ( .A1(n1036), .A2(n1035), .A3(n1034), .A4(n1033), .ZN(n1047)
         );
  AOI22_X1 U1145 ( .A1(\REGISTERS[26][5] ), .A2(n1603), .B1(\REGISTERS[15][5] ), .B2(n55), .ZN(n1040) );
  AOI22_X1 U1146 ( .A1(\REGISTERS[11][5] ), .A2(n49), .B1(\REGISTERS[19][5] ), 
        .B2(n58), .ZN(n1039) );
  AOI22_X1 U1147 ( .A1(\REGISTERS[21][5] ), .A2(n53), .B1(\REGISTERS[6][5] ), 
        .B2(n67), .ZN(n1038) );
  AOI22_X1 U1148 ( .A1(\REGISTERS[22][5] ), .A2(n51), .B1(\REGISTERS[4][5] ), 
        .B2(n37), .ZN(n1037) );
  NAND4_X1 U1149 ( .A1(n1040), .A2(n1039), .A3(n1038), .A4(n1037), .ZN(n1046)
         );
  AOI22_X1 U1150 ( .A1(\REGISTERS[29][5] ), .A2(n68), .B1(\REGISTERS[7][5] ), 
        .B2(n43), .ZN(n1044) );
  AOI22_X1 U1151 ( .A1(\REGISTERS[1][5] ), .A2(n1577), .B1(\REGISTERS[2][5] ), 
        .B2(n46), .ZN(n1043) );
  AOI22_X1 U1152 ( .A1(\REGISTERS[23][5] ), .A2(n48), .B1(\REGISTERS[27][5] ), 
        .B2(n40), .ZN(n1042) );
  AOI22_X1 U1153 ( .A1(\REGISTERS[24][5] ), .A2(n47), .B1(\REGISTERS[9][5] ), 
        .B2(n42), .ZN(n1041) );
  NAND4_X1 U1154 ( .A1(n1044), .A2(n1043), .A3(n1042), .A4(n1041), .ZN(n1045)
         );
  NOR4_X1 U1155 ( .A1(n1048), .A2(n1047), .A3(n1046), .A4(n1045), .ZN(n1049)
         );
  AOI22_X1 U1156 ( .A1(n70), .A2(n2662), .B1(n1049), .B2(n71), .ZN(N384) );
  AOI22_X1 U1157 ( .A1(\REGISTERS[21][6] ), .A2(n1599), .B1(\REGISTERS[28][6] ), .B2(n60), .ZN(n1053) );
  AOI22_X1 U1158 ( .A1(\REGISTERS[18][6] ), .A2(n59), .B1(\REGISTERS[22][6] ), 
        .B2(n51), .ZN(n1052) );
  AOI22_X1 U1159 ( .A1(\REGISTERS[11][6] ), .A2(n1591), .B1(\REGISTERS[9][6] ), 
        .B2(n42), .ZN(n1051) );
  AOI22_X1 U1160 ( .A1(\REGISTERS[16][6] ), .A2(n1613), .B1(\REGISTERS[20][6] ), .B2(n66), .ZN(n1050) );
  NAND4_X1 U1161 ( .A1(n1053), .A2(n1052), .A3(n1051), .A4(n1050), .ZN(n1069)
         );
  AOI22_X1 U1162 ( .A1(\REGISTERS[6][6] ), .A2(n1617), .B1(\REGISTERS[26][6] ), 
        .B2(n57), .ZN(n1057) );
  AOI22_X1 U1163 ( .A1(\REGISTERS[25][6] ), .A2(n61), .B1(\REGISTERS[10][6] ), 
        .B2(n41), .ZN(n1056) );
  AOI22_X1 U1164 ( .A1(\REGISTERS[5][6] ), .A2(n1612), .B1(\REGISTERS[30][6] ), 
        .B2(n65), .ZN(n1055) );
  AOI22_X1 U1165 ( .A1(\REGISTERS[3][6] ), .A2(n50), .B1(\REGISTERS[12][6] ), 
        .B2(n56), .ZN(n1054) );
  NAND4_X1 U1166 ( .A1(n1057), .A2(n1056), .A3(n1055), .A4(n1054), .ZN(n1068)
         );
  AOI22_X1 U1167 ( .A1(\REGISTERS[13][6] ), .A2(n1587), .B1(\REGISTERS[8][6] ), 
        .B2(n38), .ZN(n1061) );
  AOI22_X1 U1168 ( .A1(\REGISTERS[15][6] ), .A2(n1601), .B1(\REGISTERS[29][6] ), .B2(n68), .ZN(n1060) );
  AOI22_X1 U1169 ( .A1(\REGISTERS[27][6] ), .A2(n40), .B1(\REGISTERS[24][6] ), 
        .B2(n47), .ZN(n1059) );
  AOI22_X1 U1170 ( .A1(\REGISTERS[14][6] ), .A2(n44), .B1(\REGISTERS[2][6] ), 
        .B2(n46), .ZN(n1058) );
  NAND4_X1 U1171 ( .A1(n1061), .A2(n1060), .A3(n1059), .A4(n1058), .ZN(n1067)
         );
  AOI22_X1 U1172 ( .A1(\REGISTERS[31][6] ), .A2(n1600), .B1(\REGISTERS[1][6] ), 
        .B2(n39), .ZN(n1065) );
  AOI22_X1 U1173 ( .A1(\REGISTERS[7][6] ), .A2(n1581), .B1(\REGISTERS[4][6] ), 
        .B2(n37), .ZN(n1064) );
  AOI22_X1 U1174 ( .A1(\REGISTERS[19][6] ), .A2(n1604), .B1(\REGISTERS[17][6] ), .B2(n52), .ZN(n1063) );
  AOI22_X1 U1175 ( .A1(\REGISTERS[0][6] ), .A2(n64), .B1(\REGISTERS[23][6] ), 
        .B2(n48), .ZN(n1062) );
  NAND4_X1 U1176 ( .A1(n1065), .A2(n1064), .A3(n1063), .A4(n1062), .ZN(n1066)
         );
  NOR4_X1 U1177 ( .A1(n1069), .A2(n1068), .A3(n1067), .A4(n1066), .ZN(n1070)
         );
  AOI22_X1 U1178 ( .A1(n1628), .A2(n2659), .B1(n1070), .B2(n71), .ZN(N385) );
  AOI22_X1 U1179 ( .A1(\REGISTERS[27][7] ), .A2(n40), .B1(\REGISTERS[1][7] ), 
        .B2(n39), .ZN(n1074) );
  AOI22_X1 U1180 ( .A1(\REGISTERS[29][7] ), .A2(n68), .B1(\REGISTERS[15][7] ), 
        .B2(n55), .ZN(n1073) );
  AOI22_X1 U1181 ( .A1(\REGISTERS[5][7] ), .A2(n62), .B1(\REGISTERS[30][7] ), 
        .B2(n65), .ZN(n1072) );
  AOI22_X1 U1182 ( .A1(\REGISTERS[28][7] ), .A2(n1606), .B1(\REGISTERS[17][7] ), .B2(n52), .ZN(n1071) );
  NAND4_X1 U1183 ( .A1(n1074), .A2(n1073), .A3(n1072), .A4(n1071), .ZN(n1090)
         );
  AOI22_X1 U1184 ( .A1(\REGISTERS[2][7] ), .A2(n1588), .B1(\REGISTERS[20][7] ), 
        .B2(n66), .ZN(n1078) );
  AOI22_X1 U1185 ( .A1(\REGISTERS[25][7] ), .A2(n1611), .B1(\REGISTERS[21][7] ), .B2(n53), .ZN(n1077) );
  AOI22_X1 U1186 ( .A1(\REGISTERS[12][7] ), .A2(n1602), .B1(\REGISTERS[26][7] ), .B2(n57), .ZN(n1076) );
  AOI22_X1 U1187 ( .A1(\REGISTERS[24][7] ), .A2(n1589), .B1(\REGISTERS[4][7] ), 
        .B2(n37), .ZN(n1075) );
  NAND4_X1 U1188 ( .A1(n1078), .A2(n1077), .A3(n1076), .A4(n1075), .ZN(n1089)
         );
  AOI22_X1 U1189 ( .A1(\REGISTERS[10][7] ), .A2(n1579), .B1(\REGISTERS[11][7] ), .B2(n49), .ZN(n1082) );
  AOI22_X1 U1190 ( .A1(\REGISTERS[16][7] ), .A2(n1613), .B1(\REGISTERS[18][7] ), .B2(n59), .ZN(n1081) );
  AOI22_X1 U1191 ( .A1(\REGISTERS[31][7] ), .A2(n1600), .B1(\REGISTERS[14][7] ), .B2(n44), .ZN(n1080) );
  AOI22_X1 U1192 ( .A1(\REGISTERS[9][7] ), .A2(n42), .B1(\REGISTERS[22][7] ), 
        .B2(n51), .ZN(n1079) );
  NAND4_X1 U1193 ( .A1(n1082), .A2(n1081), .A3(n1080), .A4(n1079), .ZN(n1088)
         );
  AOI22_X1 U1194 ( .A1(\REGISTERS[6][7] ), .A2(n67), .B1(\REGISTERS[13][7] ), 
        .B2(n45), .ZN(n1086) );
  AOI22_X1 U1195 ( .A1(\REGISTERS[7][7] ), .A2(n1581), .B1(\REGISTERS[3][7] ), 
        .B2(n50), .ZN(n1085) );
  AOI22_X1 U1196 ( .A1(\REGISTERS[19][7] ), .A2(n58), .B1(\REGISTERS[8][7] ), 
        .B2(n38), .ZN(n1084) );
  AOI22_X1 U1197 ( .A1(\REGISTERS[23][7] ), .A2(n1590), .B1(\REGISTERS[0][7] ), 
        .B2(n64), .ZN(n1083) );
  NAND4_X1 U1198 ( .A1(n1086), .A2(n1085), .A3(n1084), .A4(n1083), .ZN(n1087)
         );
  NOR4_X1 U1199 ( .A1(n1090), .A2(n1089), .A3(n1088), .A4(n1087), .ZN(n1091)
         );
  AOI22_X1 U1200 ( .A1(n1628), .A2(n122), .B1(n1091), .B2(n72), .ZN(N386) );
  AOI22_X1 U1201 ( .A1(\REGISTERS[30][8] ), .A2(n1615), .B1(\REGISTERS[24][8] ), .B2(n47), .ZN(n1095) );
  AOI22_X1 U1202 ( .A1(\REGISTERS[0][8] ), .A2(n1614), .B1(\REGISTERS[16][8] ), 
        .B2(n63), .ZN(n1094) );
  AOI22_X1 U1203 ( .A1(\REGISTERS[13][8] ), .A2(n1587), .B1(\REGISTERS[20][8] ), .B2(n66), .ZN(n1093) );
  AOI22_X1 U1204 ( .A1(\REGISTERS[14][8] ), .A2(n44), .B1(\REGISTERS[2][8] ), 
        .B2(n46), .ZN(n1092) );
  NAND4_X1 U1205 ( .A1(n1095), .A2(n1094), .A3(n1093), .A4(n1092), .ZN(n1111)
         );
  AOI22_X1 U1206 ( .A1(\REGISTERS[31][8] ), .A2(n54), .B1(\REGISTERS[15][8] ), 
        .B2(n55), .ZN(n1099) );
  AOI22_X1 U1207 ( .A1(\REGISTERS[27][8] ), .A2(n40), .B1(\REGISTERS[12][8] ), 
        .B2(n56), .ZN(n1098) );
  AOI22_X1 U1208 ( .A1(\REGISTERS[7][8] ), .A2(n1581), .B1(\REGISTERS[22][8] ), 
        .B2(n51), .ZN(n1097) );
  AOI22_X1 U1209 ( .A1(\REGISTERS[21][8] ), .A2(n1599), .B1(\REGISTERS[9][8] ), 
        .B2(n42), .ZN(n1096) );
  NAND4_X1 U1210 ( .A1(n1099), .A2(n1098), .A3(n1097), .A4(n1096), .ZN(n1110)
         );
  AOI22_X1 U1211 ( .A1(\REGISTERS[29][8] ), .A2(n1618), .B1(\REGISTERS[6][8] ), 
        .B2(n67), .ZN(n1103) );
  AOI22_X1 U1212 ( .A1(\REGISTERS[25][8] ), .A2(n1611), .B1(\REGISTERS[5][8] ), 
        .B2(n62), .ZN(n1102) );
  AOI22_X1 U1213 ( .A1(\REGISTERS[26][8] ), .A2(n57), .B1(\REGISTERS[17][8] ), 
        .B2(n52), .ZN(n1101) );
  AOI22_X1 U1214 ( .A1(\REGISTERS[8][8] ), .A2(n1576), .B1(\REGISTERS[11][8] ), 
        .B2(n49), .ZN(n1100) );
  NAND4_X1 U1215 ( .A1(n1103), .A2(n1102), .A3(n1101), .A4(n1100), .ZN(n1109)
         );
  AOI22_X1 U1216 ( .A1(\REGISTERS[19][8] ), .A2(n58), .B1(\REGISTERS[1][8] ), 
        .B2(n39), .ZN(n1107) );
  AOI22_X1 U1217 ( .A1(\REGISTERS[3][8] ), .A2(n50), .B1(\REGISTERS[18][8] ), 
        .B2(n59), .ZN(n1106) );
  AOI22_X1 U1218 ( .A1(\REGISTERS[28][8] ), .A2(n1606), .B1(\REGISTERS[10][8] ), .B2(n41), .ZN(n1105) );
  AOI22_X1 U1219 ( .A1(\REGISTERS[4][8] ), .A2(n1575), .B1(\REGISTERS[23][8] ), 
        .B2(n48), .ZN(n1104) );
  NAND4_X1 U1220 ( .A1(n1107), .A2(n1106), .A3(n1105), .A4(n1104), .ZN(n1108)
         );
  NOR4_X1 U1221 ( .A1(n1111), .A2(n1110), .A3(n1109), .A4(n1108), .ZN(n1112)
         );
  AOI22_X1 U1222 ( .A1(n1628), .A2(n2675), .B1(n1112), .B2(n72), .ZN(N387) );
  AOI22_X1 U1223 ( .A1(\REGISTERS[15][9] ), .A2(n1601), .B1(\REGISTERS[26][9] ), .B2(n57), .ZN(n1116) );
  AOI22_X1 U1224 ( .A1(\REGISTERS[2][9] ), .A2(n1588), .B1(\REGISTERS[25][9] ), 
        .B2(n61), .ZN(n1115) );
  AOI22_X1 U1225 ( .A1(\REGISTERS[19][9] ), .A2(n58), .B1(\REGISTERS[24][9] ), 
        .B2(n47), .ZN(n1114) );
  AOI22_X1 U1226 ( .A1(\REGISTERS[3][9] ), .A2(n50), .B1(\REGISTERS[16][9] ), 
        .B2(n63), .ZN(n1113) );
  NAND4_X1 U1227 ( .A1(n1116), .A2(n1115), .A3(n1114), .A4(n1113), .ZN(n1132)
         );
  AOI22_X1 U1228 ( .A1(\REGISTERS[21][9] ), .A2(n1599), .B1(\REGISTERS[6][9] ), 
        .B2(n67), .ZN(n1120) );
  AOI22_X1 U1229 ( .A1(\REGISTERS[5][9] ), .A2(n1612), .B1(\REGISTERS[9][9] ), 
        .B2(n42), .ZN(n1119) );
  AOI22_X1 U1230 ( .A1(\REGISTERS[31][9] ), .A2(n54), .B1(\REGISTERS[11][9] ), 
        .B2(n49), .ZN(n1118) );
  AOI22_X1 U1231 ( .A1(\REGISTERS[27][9] ), .A2(n40), .B1(\REGISTERS[13][9] ), 
        .B2(n45), .ZN(n1117) );
  NAND4_X1 U1232 ( .A1(n1120), .A2(n1119), .A3(n1118), .A4(n1117), .ZN(n1131)
         );
  AOI22_X1 U1233 ( .A1(\REGISTERS[22][9] ), .A2(n1593), .B1(\REGISTERS[7][9] ), 
        .B2(n43), .ZN(n1124) );
  AOI22_X1 U1234 ( .A1(\REGISTERS[8][9] ), .A2(n1576), .B1(\REGISTERS[20][9] ), 
        .B2(n66), .ZN(n1123) );
  AOI22_X1 U1235 ( .A1(\REGISTERS[14][9] ), .A2(n44), .B1(\REGISTERS[1][9] ), 
        .B2(n39), .ZN(n1122) );
  AOI22_X1 U1236 ( .A1(\REGISTERS[17][9] ), .A2(n52), .B1(\REGISTERS[28][9] ), 
        .B2(n60), .ZN(n1121) );
  NAND4_X1 U1237 ( .A1(n1124), .A2(n1123), .A3(n1122), .A4(n1121), .ZN(n1130)
         );
  AOI22_X1 U1238 ( .A1(\REGISTERS[30][9] ), .A2(n1615), .B1(\REGISTERS[12][9] ), .B2(n56), .ZN(n1128) );
  AOI22_X1 U1239 ( .A1(\REGISTERS[29][9] ), .A2(n1618), .B1(\REGISTERS[4][9] ), 
        .B2(n37), .ZN(n1127) );
  AOI22_X1 U1240 ( .A1(\REGISTERS[10][9] ), .A2(n1579), .B1(\REGISTERS[0][9] ), 
        .B2(n64), .ZN(n1126) );
  AOI22_X1 U1241 ( .A1(\REGISTERS[18][9] ), .A2(n59), .B1(\REGISTERS[23][9] ), 
        .B2(n48), .ZN(n1125) );
  NAND4_X1 U1242 ( .A1(n1128), .A2(n1127), .A3(n1126), .A4(n1125), .ZN(n1129)
         );
  NOR4_X1 U1243 ( .A1(n1132), .A2(n1131), .A3(n1130), .A4(n1129), .ZN(n1133)
         );
  AOI22_X1 U1244 ( .A1(n1628), .A2(n2674), .B1(n1133), .B2(n71), .ZN(N388) );
  AOI22_X1 U1245 ( .A1(\REGISTERS[3][10] ), .A2(n50), .B1(\REGISTERS[9][10] ), 
        .B2(n42), .ZN(n1137) );
  AOI22_X1 U1246 ( .A1(\REGISTERS[27][10] ), .A2(n1578), .B1(
        \REGISTERS[17][10] ), .B2(n52), .ZN(n1136) );
  AOI22_X1 U1247 ( .A1(\REGISTERS[2][10] ), .A2(n1588), .B1(
        \REGISTERS[18][10] ), .B2(n59), .ZN(n1135) );
  AOI22_X1 U1248 ( .A1(\REGISTERS[4][10] ), .A2(n1575), .B1(
        \REGISTERS[19][10] ), .B2(n58), .ZN(n1134) );
  NAND4_X1 U1249 ( .A1(n1137), .A2(n1136), .A3(n1135), .A4(n1134), .ZN(n1153)
         );
  AOI22_X1 U1250 ( .A1(\REGISTERS[23][10] ), .A2(n1590), .B1(
        \REGISTERS[8][10] ), .B2(n38), .ZN(n1141) );
  AOI22_X1 U1251 ( .A1(\REGISTERS[1][10] ), .A2(n1577), .B1(
        \REGISTERS[16][10] ), .B2(n63), .ZN(n1140) );
  AOI22_X1 U1252 ( .A1(\REGISTERS[24][10] ), .A2(n1589), .B1(
        \REGISTERS[26][10] ), .B2(n57), .ZN(n1139) );
  AOI22_X1 U1253 ( .A1(\REGISTERS[31][10] ), .A2(n54), .B1(\REGISTERS[11][10] ), .B2(n49), .ZN(n1138) );
  NAND4_X1 U1254 ( .A1(n1141), .A2(n1140), .A3(n1139), .A4(n1138), .ZN(n1152)
         );
  AOI22_X1 U1255 ( .A1(\REGISTERS[22][10] ), .A2(n1593), .B1(
        \REGISTERS[29][10] ), .B2(n68), .ZN(n1145) );
  AOI22_X1 U1256 ( .A1(\REGISTERS[15][10] ), .A2(n1601), .B1(
        \REGISTERS[0][10] ), .B2(n64), .ZN(n1144) );
  AOI22_X1 U1257 ( .A1(\REGISTERS[10][10] ), .A2(n1579), .B1(
        \REGISTERS[25][10] ), .B2(n61), .ZN(n1143) );
  AOI22_X1 U1258 ( .A1(\REGISTERS[14][10] ), .A2(n1582), .B1(
        \REGISTERS[6][10] ), .B2(n67), .ZN(n1142) );
  NAND4_X1 U1259 ( .A1(n1145), .A2(n1144), .A3(n1143), .A4(n1142), .ZN(n1151)
         );
  AOI22_X1 U1260 ( .A1(\REGISTERS[20][10] ), .A2(n66), .B1(\REGISTERS[7][10] ), 
        .B2(n43), .ZN(n1149) );
  AOI22_X1 U1261 ( .A1(\REGISTERS[12][10] ), .A2(n56), .B1(\REGISTERS[28][10] ), .B2(n60), .ZN(n1148) );
  AOI22_X1 U1262 ( .A1(\REGISTERS[21][10] ), .A2(n1599), .B1(
        \REGISTERS[30][10] ), .B2(n65), .ZN(n1147) );
  AOI22_X1 U1263 ( .A1(\REGISTERS[5][10] ), .A2(n1612), .B1(
        \REGISTERS[13][10] ), .B2(n45), .ZN(n1146) );
  NAND4_X1 U1264 ( .A1(n1149), .A2(n1148), .A3(n1147), .A4(n1146), .ZN(n1150)
         );
  NOR4_X1 U1265 ( .A1(n1153), .A2(n1152), .A3(n1151), .A4(n1150), .ZN(n1154)
         );
  AOI22_X1 U1266 ( .A1(n1628), .A2(n2661), .B1(n1154), .B2(n72), .ZN(N389) );
  AOI22_X1 U1267 ( .A1(\REGISTERS[23][11] ), .A2(n1590), .B1(
        \REGISTERS[21][11] ), .B2(n53), .ZN(n1158) );
  AOI22_X1 U1268 ( .A1(\REGISTERS[10][11] ), .A2(n1579), .B1(
        \REGISTERS[6][11] ), .B2(n67), .ZN(n1157) );
  AOI22_X1 U1269 ( .A1(\REGISTERS[2][11] ), .A2(n1588), .B1(
        \REGISTERS[14][11] ), .B2(n44), .ZN(n1156) );
  AOI22_X1 U1270 ( .A1(\REGISTERS[9][11] ), .A2(n42), .B1(\REGISTERS[7][11] ), 
        .B2(n43), .ZN(n1155) );
  NAND4_X1 U1271 ( .A1(n1158), .A2(n1157), .A3(n1156), .A4(n1155), .ZN(n1174)
         );
  AOI22_X1 U1272 ( .A1(\REGISTERS[1][11] ), .A2(n1577), .B1(
        \REGISTERS[27][11] ), .B2(n40), .ZN(n1162) );
  AOI22_X1 U1273 ( .A1(\REGISTERS[13][11] ), .A2(n1587), .B1(
        \REGISTERS[11][11] ), .B2(n49), .ZN(n1161) );
  AOI22_X1 U1274 ( .A1(\REGISTERS[18][11] ), .A2(n1605), .B1(
        \REGISTERS[24][11] ), .B2(n47), .ZN(n1160) );
  AOI22_X1 U1275 ( .A1(\REGISTERS[3][11] ), .A2(n1592), .B1(
        \REGISTERS[20][11] ), .B2(n66), .ZN(n1159) );
  NAND4_X1 U1276 ( .A1(n1162), .A2(n1161), .A3(n1160), .A4(n1159), .ZN(n1173)
         );
  AOI22_X1 U1277 ( .A1(\REGISTERS[29][11] ), .A2(n1618), .B1(
        \REGISTERS[4][11] ), .B2(n37), .ZN(n1166) );
  AOI22_X1 U1278 ( .A1(\REGISTERS[25][11] ), .A2(n1611), .B1(
        \REGISTERS[30][11] ), .B2(n65), .ZN(n1165) );
  AOI22_X1 U1279 ( .A1(\REGISTERS[8][11] ), .A2(n1576), .B1(
        \REGISTERS[22][11] ), .B2(n51), .ZN(n1164) );
  AOI22_X1 U1280 ( .A1(\REGISTERS[19][11] ), .A2(n58), .B1(\REGISTERS[5][11] ), 
        .B2(n62), .ZN(n1163) );
  NAND4_X1 U1281 ( .A1(n1166), .A2(n1165), .A3(n1164), .A4(n1163), .ZN(n1172)
         );
  AOI22_X1 U1282 ( .A1(\REGISTERS[26][11] ), .A2(n1603), .B1(
        \REGISTERS[15][11] ), .B2(n55), .ZN(n1170) );
  AOI22_X1 U1283 ( .A1(\REGISTERS[31][11] ), .A2(n1600), .B1(
        \REGISTERS[0][11] ), .B2(n64), .ZN(n1169) );
  AOI22_X1 U1284 ( .A1(\REGISTERS[17][11] ), .A2(n52), .B1(\REGISTERS[28][11] ), .B2(n60), .ZN(n1168) );
  AOI22_X1 U1285 ( .A1(\REGISTERS[12][11] ), .A2(n56), .B1(\REGISTERS[16][11] ), .B2(n63), .ZN(n1167) );
  NAND4_X1 U1286 ( .A1(n1170), .A2(n1169), .A3(n1168), .A4(n1167), .ZN(n1171)
         );
  NOR4_X1 U1287 ( .A1(n1174), .A2(n1173), .A3(n1172), .A4(n1171), .ZN(n1175)
         );
  AOI22_X1 U1288 ( .A1(n1628), .A2(n114), .B1(n1175), .B2(n71), .ZN(N390) );
  AOI22_X1 U1289 ( .A1(\REGISTERS[25][12] ), .A2(n1611), .B1(
        \REGISTERS[8][12] ), .B2(n38), .ZN(n1179) );
  AOI22_X1 U1290 ( .A1(\REGISTERS[21][12] ), .A2(n1599), .B1(
        \REGISTERS[30][12] ), .B2(n65), .ZN(n1178) );
  AOI22_X1 U1291 ( .A1(\REGISTERS[26][12] ), .A2(n1603), .B1(
        \REGISTERS[18][12] ), .B2(n59), .ZN(n1177) );
  AOI22_X1 U1292 ( .A1(\REGISTERS[19][12] ), .A2(n58), .B1(\REGISTERS[22][12] ), .B2(n51), .ZN(n1176) );
  NAND4_X1 U1293 ( .A1(n1179), .A2(n1178), .A3(n1177), .A4(n1176), .ZN(n1195)
         );
  AOI22_X1 U1294 ( .A1(\REGISTERS[3][12] ), .A2(n1592), .B1(
        \REGISTERS[10][12] ), .B2(n41), .ZN(n1183) );
  AOI22_X1 U1295 ( .A1(\REGISTERS[11][12] ), .A2(n1591), .B1(
        \REGISTERS[5][12] ), .B2(n62), .ZN(n1182) );
  AOI22_X1 U1296 ( .A1(\REGISTERS[4][12] ), .A2(n1575), .B1(
        \REGISTERS[23][12] ), .B2(n48), .ZN(n1181) );
  AOI22_X1 U1297 ( .A1(\REGISTERS[20][12] ), .A2(n1616), .B1(
        \REGISTERS[0][12] ), .B2(n64), .ZN(n1180) );
  NAND4_X1 U1298 ( .A1(n1183), .A2(n1182), .A3(n1181), .A4(n1180), .ZN(n1194)
         );
  AOI22_X1 U1299 ( .A1(\REGISTERS[6][12] ), .A2(n1617), .B1(
        \REGISTERS[28][12] ), .B2(n60), .ZN(n1187) );
  AOI22_X1 U1300 ( .A1(\REGISTERS[9][12] ), .A2(n1580), .B1(
        \REGISTERS[15][12] ), .B2(n55), .ZN(n1186) );
  AOI22_X1 U1301 ( .A1(\REGISTERS[2][12] ), .A2(n1588), .B1(
        \REGISTERS[27][12] ), .B2(n40), .ZN(n1185) );
  AOI22_X1 U1302 ( .A1(\REGISTERS[31][12] ), .A2(n1600), .B1(
        \REGISTERS[1][12] ), .B2(n39), .ZN(n1184) );
  NAND4_X1 U1303 ( .A1(n1187), .A2(n1186), .A3(n1185), .A4(n1184), .ZN(n1193)
         );
  AOI22_X1 U1304 ( .A1(\REGISTERS[17][12] ), .A2(n52), .B1(\REGISTERS[13][12] ), .B2(n45), .ZN(n1191) );
  AOI22_X1 U1305 ( .A1(\REGISTERS[16][12] ), .A2(n1613), .B1(
        \REGISTERS[12][12] ), .B2(n56), .ZN(n1190) );
  AOI22_X1 U1306 ( .A1(\REGISTERS[14][12] ), .A2(n1582), .B1(
        \REGISTERS[7][12] ), .B2(n43), .ZN(n1189) );
  AOI22_X1 U1307 ( .A1(\REGISTERS[24][12] ), .A2(n1589), .B1(
        \REGISTERS[29][12] ), .B2(n68), .ZN(n1188) );
  NAND4_X1 U1308 ( .A1(n1191), .A2(n1190), .A3(n1189), .A4(n1188), .ZN(n1192)
         );
  NOR4_X1 U1309 ( .A1(n1195), .A2(n1194), .A3(n1193), .A4(n1192), .ZN(n1196)
         );
  AOI22_X1 U1310 ( .A1(n69), .A2(n2666), .B1(n1196), .B2(n72), .ZN(N391) );
  AOI22_X1 U1311 ( .A1(\REGISTERS[31][13] ), .A2(n1600), .B1(
        \REGISTERS[27][13] ), .B2(n40), .ZN(n1200) );
  AOI22_X1 U1312 ( .A1(\REGISTERS[22][13] ), .A2(n1593), .B1(
        \REGISTERS[8][13] ), .B2(n38), .ZN(n1199) );
  AOI22_X1 U1313 ( .A1(\REGISTERS[14][13] ), .A2(n1582), .B1(
        \REGISTERS[21][13] ), .B2(n53), .ZN(n1198) );
  AOI22_X1 U1314 ( .A1(\REGISTERS[5][13] ), .A2(n1612), .B1(\REGISTERS[6][13] ), .B2(n1617), .ZN(n1197) );
  NAND4_X1 U1315 ( .A1(n1200), .A2(n1199), .A3(n1198), .A4(n1197), .ZN(n1216)
         );
  AOI22_X1 U1316 ( .A1(\REGISTERS[12][13] ), .A2(n56), .B1(\REGISTERS[4][13] ), 
        .B2(n37), .ZN(n1204) );
  AOI22_X1 U1317 ( .A1(\REGISTERS[13][13] ), .A2(n1587), .B1(
        \REGISTERS[30][13] ), .B2(n65), .ZN(n1203) );
  AOI22_X1 U1318 ( .A1(\REGISTERS[17][13] ), .A2(n1594), .B1(
        \REGISTERS[3][13] ), .B2(n50), .ZN(n1202) );
  AOI22_X1 U1319 ( .A1(\REGISTERS[11][13] ), .A2(n1591), .B1(
        \REGISTERS[20][13] ), .B2(n66), .ZN(n1201) );
  NAND4_X1 U1320 ( .A1(n1204), .A2(n1203), .A3(n1202), .A4(n1201), .ZN(n1215)
         );
  AOI22_X1 U1321 ( .A1(\REGISTERS[23][13] ), .A2(n1590), .B1(
        \REGISTERS[18][13] ), .B2(n59), .ZN(n1208) );
  AOI22_X1 U1322 ( .A1(\REGISTERS[0][13] ), .A2(n1614), .B1(
        \REGISTERS[29][13] ), .B2(n68), .ZN(n1207) );
  AOI22_X1 U1323 ( .A1(\REGISTERS[9][13] ), .A2(n1580), .B1(
        \REGISTERS[26][13] ), .B2(n57), .ZN(n1206) );
  AOI22_X1 U1324 ( .A1(\REGISTERS[28][13] ), .A2(n1606), .B1(
        \REGISTERS[7][13] ), .B2(n43), .ZN(n1205) );
  NAND4_X1 U1325 ( .A1(n1208), .A2(n1207), .A3(n1206), .A4(n1205), .ZN(n1214)
         );
  AOI22_X1 U1326 ( .A1(\REGISTERS[24][13] ), .A2(n1589), .B1(
        \REGISTERS[16][13] ), .B2(n63), .ZN(n1212) );
  AOI22_X1 U1327 ( .A1(\REGISTERS[19][13] ), .A2(n58), .B1(\REGISTERS[1][13] ), 
        .B2(n39), .ZN(n1211) );
  AOI22_X1 U1328 ( .A1(\REGISTERS[10][13] ), .A2(n1579), .B1(
        \REGISTERS[25][13] ), .B2(n61), .ZN(n1210) );
  AOI22_X1 U1329 ( .A1(\REGISTERS[2][13] ), .A2(n1588), .B1(
        \REGISTERS[15][13] ), .B2(n55), .ZN(n1209) );
  NAND4_X1 U1330 ( .A1(n1212), .A2(n1211), .A3(n1210), .A4(n1209), .ZN(n1213)
         );
  NOR4_X1 U1331 ( .A1(n1216), .A2(n1215), .A3(n1214), .A4(n1213), .ZN(n1217)
         );
  AOI22_X1 U1332 ( .A1(n69), .A2(n110), .B1(n1217), .B2(n71), .ZN(N392) );
  AOI22_X1 U1333 ( .A1(\REGISTERS[22][14] ), .A2(n1593), .B1(
        \REGISTERS[13][14] ), .B2(n45), .ZN(n1221) );
  AOI22_X1 U1334 ( .A1(\REGISTERS[7][14] ), .A2(n1581), .B1(\REGISTERS[5][14] ), .B2(n62), .ZN(n1220) );
  AOI22_X1 U1335 ( .A1(\REGISTERS[26][14] ), .A2(n1603), .B1(
        \REGISTERS[27][14] ), .B2(n40), .ZN(n1219) );
  AOI22_X1 U1336 ( .A1(\REGISTERS[20][14] ), .A2(n1616), .B1(
        \REGISTERS[25][14] ), .B2(n61), .ZN(n1218) );
  NAND4_X1 U1337 ( .A1(n1221), .A2(n1220), .A3(n1219), .A4(n1218), .ZN(n1237)
         );
  AOI22_X1 U1338 ( .A1(\REGISTERS[4][14] ), .A2(n1575), .B1(
        \REGISTERS[18][14] ), .B2(n59), .ZN(n1225) );
  AOI22_X1 U1339 ( .A1(\REGISTERS[12][14] ), .A2(n1602), .B1(
        \REGISTERS[1][14] ), .B2(n39), .ZN(n1224) );
  AOI22_X1 U1340 ( .A1(\REGISTERS[24][14] ), .A2(n47), .B1(\REGISTERS[14][14] ), .B2(n44), .ZN(n1223) );
  AOI22_X1 U1341 ( .A1(\REGISTERS[19][14] ), .A2(n58), .B1(\REGISTERS[9][14] ), 
        .B2(n42), .ZN(n1222) );
  NAND4_X1 U1342 ( .A1(n1225), .A2(n1224), .A3(n1223), .A4(n1222), .ZN(n1236)
         );
  AOI22_X1 U1343 ( .A1(\REGISTERS[17][14] ), .A2(n1594), .B1(
        \REGISTERS[11][14] ), .B2(n49), .ZN(n1229) );
  AOI22_X1 U1344 ( .A1(\REGISTERS[31][14] ), .A2(n1600), .B1(
        \REGISTERS[30][14] ), .B2(n65), .ZN(n1228) );
  AOI22_X1 U1345 ( .A1(\REGISTERS[28][14] ), .A2(n1606), .B1(
        \REGISTERS[10][14] ), .B2(n41), .ZN(n1227) );
  AOI22_X1 U1346 ( .A1(\REGISTERS[2][14] ), .A2(n1588), .B1(
        \REGISTERS[21][14] ), .B2(n53), .ZN(n1226) );
  NAND4_X1 U1347 ( .A1(n1229), .A2(n1228), .A3(n1227), .A4(n1226), .ZN(n1235)
         );
  AOI22_X1 U1348 ( .A1(\REGISTERS[29][14] ), .A2(n1618), .B1(
        \REGISTERS[23][14] ), .B2(n48), .ZN(n1233) );
  AOI22_X1 U1349 ( .A1(\REGISTERS[0][14] ), .A2(n1614), .B1(
        \REGISTERS[15][14] ), .B2(n55), .ZN(n1232) );
  AOI22_X1 U1350 ( .A1(\REGISTERS[16][14] ), .A2(n1613), .B1(
        \REGISTERS[6][14] ), .B2(n67), .ZN(n1231) );
  AOI22_X1 U1351 ( .A1(\REGISTERS[8][14] ), .A2(n1576), .B1(\REGISTERS[3][14] ), .B2(n50), .ZN(n1230) );
  NAND4_X1 U1352 ( .A1(n1233), .A2(n1232), .A3(n1231), .A4(n1230), .ZN(n1234)
         );
  NOR4_X1 U1353 ( .A1(n1237), .A2(n1236), .A3(n1235), .A4(n1234), .ZN(n1238)
         );
  AOI22_X1 U1354 ( .A1(n69), .A2(n2660), .B1(n1238), .B2(n72), .ZN(N393) );
  AOI22_X1 U1355 ( .A1(\REGISTERS[16][15] ), .A2(n63), .B1(\REGISTERS[30][15] ), .B2(n1615), .ZN(n1242) );
  AOI22_X1 U1356 ( .A1(\REGISTERS[29][15] ), .A2(n1618), .B1(
        \REGISTERS[12][15] ), .B2(n56), .ZN(n1241) );
  AOI22_X1 U1357 ( .A1(\REGISTERS[24][15] ), .A2(n47), .B1(\REGISTERS[10][15] ), .B2(n41), .ZN(n1240) );
  AOI22_X1 U1358 ( .A1(\REGISTERS[18][15] ), .A2(n1605), .B1(
        \REGISTERS[14][15] ), .B2(n44), .ZN(n1239) );
  NAND4_X1 U1359 ( .A1(n1242), .A2(n1241), .A3(n1240), .A4(n1239), .ZN(n1258)
         );
  AOI22_X1 U1360 ( .A1(\REGISTERS[20][15] ), .A2(n66), .B1(\REGISTERS[26][15] ), .B2(n57), .ZN(n1246) );
  AOI22_X1 U1361 ( .A1(\REGISTERS[6][15] ), .A2(n1617), .B1(\REGISTERS[4][15] ), .B2(n37), .ZN(n1245) );
  AOI22_X1 U1362 ( .A1(\REGISTERS[7][15] ), .A2(n1581), .B1(\REGISTERS[8][15] ), .B2(n38), .ZN(n1244) );
  AOI22_X1 U1363 ( .A1(\REGISTERS[19][15] ), .A2(n58), .B1(\REGISTERS[2][15] ), 
        .B2(n46), .ZN(n1243) );
  NAND4_X1 U1364 ( .A1(n1246), .A2(n1245), .A3(n1244), .A4(n1243), .ZN(n1257)
         );
  AOI22_X1 U1365 ( .A1(\REGISTERS[17][15] ), .A2(n1594), .B1(
        \REGISTERS[23][15] ), .B2(n48), .ZN(n1250) );
  AOI22_X1 U1366 ( .A1(\REGISTERS[27][15] ), .A2(n1578), .B1(
        \REGISTERS[28][15] ), .B2(n60), .ZN(n1249) );
  AOI22_X1 U1367 ( .A1(\REGISTERS[25][15] ), .A2(n1611), .B1(
        \REGISTERS[15][15] ), .B2(n1601), .ZN(n1248) );
  AOI22_X1 U1368 ( .A1(\REGISTERS[3][15] ), .A2(n1592), .B1(\REGISTERS[9][15] ), .B2(n42), .ZN(n1247) );
  NAND4_X1 U1369 ( .A1(n1250), .A2(n1249), .A3(n1248), .A4(n1247), .ZN(n1256)
         );
  AOI22_X1 U1370 ( .A1(\REGISTERS[22][15] ), .A2(n51), .B1(\REGISTERS[5][15] ), 
        .B2(n62), .ZN(n1254) );
  AOI22_X1 U1371 ( .A1(\REGISTERS[0][15] ), .A2(n1614), .B1(\REGISTERS[1][15] ), .B2(n39), .ZN(n1253) );
  AOI22_X1 U1372 ( .A1(\REGISTERS[31][15] ), .A2(n1600), .B1(
        \REGISTERS[11][15] ), .B2(n1591), .ZN(n1252) );
  AOI22_X1 U1373 ( .A1(\REGISTERS[13][15] ), .A2(n1587), .B1(
        \REGISTERS[21][15] ), .B2(n53), .ZN(n1251) );
  NAND4_X1 U1374 ( .A1(n1254), .A2(n1253), .A3(n1252), .A4(n1251), .ZN(n1255)
         );
  NOR4_X1 U1375 ( .A1(n1258), .A2(n1257), .A3(n1256), .A4(n1255), .ZN(n1259)
         );
  AOI22_X1 U1376 ( .A1(n69), .A2(n2658), .B1(n1259), .B2(n71), .ZN(N394) );
  AOI22_X1 U1377 ( .A1(\REGISTERS[11][16] ), .A2(n1591), .B1(
        \REGISTERS[3][16] ), .B2(n50), .ZN(n1263) );
  AOI22_X1 U1378 ( .A1(\REGISTERS[12][16] ), .A2(n1602), .B1(
        \REGISTERS[20][16] ), .B2(n66), .ZN(n1262) );
  AOI22_X1 U1379 ( .A1(\REGISTERS[29][16] ), .A2(n1618), .B1(
        \REGISTERS[23][16] ), .B2(n48), .ZN(n1261) );
  AOI22_X1 U1380 ( .A1(\REGISTERS[6][16] ), .A2(n1617), .B1(\REGISTERS[0][16] ), .B2(n64), .ZN(n1260) );
  NAND4_X1 U1381 ( .A1(n1263), .A2(n1262), .A3(n1261), .A4(n1260), .ZN(n1279)
         );
  AOI22_X1 U1382 ( .A1(\REGISTERS[17][16] ), .A2(n1594), .B1(
        \REGISTERS[2][16] ), .B2(n46), .ZN(n1267) );
  AOI22_X1 U1383 ( .A1(\REGISTERS[18][16] ), .A2(n1605), .B1(
        \REGISTERS[24][16] ), .B2(n47), .ZN(n1266) );
  AOI22_X1 U1384 ( .A1(\REGISTERS[22][16] ), .A2(n51), .B1(\REGISTERS[5][16] ), 
        .B2(n62), .ZN(n1265) );
  AOI22_X1 U1385 ( .A1(\REGISTERS[4][16] ), .A2(n1575), .B1(
        \REGISTERS[28][16] ), .B2(n60), .ZN(n1264) );
  NAND4_X1 U1386 ( .A1(n1267), .A2(n1266), .A3(n1265), .A4(n1264), .ZN(n1278)
         );
  AOI22_X1 U1387 ( .A1(\REGISTERS[27][16] ), .A2(n1578), .B1(
        \REGISTERS[26][16] ), .B2(n57), .ZN(n1271) );
  AOI22_X1 U1388 ( .A1(\REGISTERS[9][16] ), .A2(n1580), .B1(
        \REGISTERS[14][16] ), .B2(n44), .ZN(n1270) );
  AOI22_X1 U1389 ( .A1(\REGISTERS[16][16] ), .A2(n1613), .B1(
        \REGISTERS[1][16] ), .B2(n39), .ZN(n1269) );
  AOI22_X1 U1390 ( .A1(\REGISTERS[19][16] ), .A2(n58), .B1(\REGISTERS[30][16] ), .B2(n1615), .ZN(n1268) );
  NAND4_X1 U1391 ( .A1(n1271), .A2(n1270), .A3(n1269), .A4(n1268), .ZN(n1277)
         );
  AOI22_X1 U1392 ( .A1(\REGISTERS[25][16] ), .A2(n1611), .B1(
        \REGISTERS[15][16] ), .B2(n1601), .ZN(n1275) );
  AOI22_X1 U1393 ( .A1(\REGISTERS[7][16] ), .A2(n1581), .B1(
        \REGISTERS[31][16] ), .B2(n54), .ZN(n1274) );
  AOI22_X1 U1394 ( .A1(\REGISTERS[13][16] ), .A2(n1587), .B1(
        \REGISTERS[21][16] ), .B2(n53), .ZN(n1273) );
  AOI22_X1 U1395 ( .A1(\REGISTERS[10][16] ), .A2(n41), .B1(\REGISTERS[8][16] ), 
        .B2(n38), .ZN(n1272) );
  NAND4_X1 U1396 ( .A1(n1275), .A2(n1274), .A3(n1273), .A4(n1272), .ZN(n1276)
         );
  NOR4_X1 U1397 ( .A1(n1279), .A2(n1278), .A3(n1277), .A4(n1276), .ZN(n1280)
         );
  AOI22_X1 U1398 ( .A1(n69), .A2(n2668), .B1(n1280), .B2(n72), .ZN(N395) );
  AOI22_X1 U1399 ( .A1(\REGISTERS[24][17] ), .A2(n1589), .B1(
        \REGISTERS[0][17] ), .B2(n64), .ZN(n1284) );
  AOI22_X1 U1400 ( .A1(\REGISTERS[6][17] ), .A2(n1617), .B1(
        \REGISTERS[29][17] ), .B2(n68), .ZN(n1283) );
  AOI22_X1 U1401 ( .A1(\REGISTERS[5][17] ), .A2(n1612), .B1(
        \REGISTERS[21][17] ), .B2(n53), .ZN(n1282) );
  AOI22_X1 U1402 ( .A1(\REGISTERS[28][17] ), .A2(n1606), .B1(
        \REGISTERS[1][17] ), .B2(n39), .ZN(n1281) );
  NAND4_X1 U1403 ( .A1(n1284), .A2(n1283), .A3(n1282), .A4(n1281), .ZN(n1300)
         );
  AOI22_X1 U1404 ( .A1(\REGISTERS[14][17] ), .A2(n1582), .B1(
        \REGISTERS[16][17] ), .B2(n63), .ZN(n1288) );
  AOI22_X1 U1405 ( .A1(\REGISTERS[27][17] ), .A2(n1578), .B1(
        \REGISTERS[25][17] ), .B2(n61), .ZN(n1287) );
  AOI22_X1 U1406 ( .A1(\REGISTERS[3][17] ), .A2(n1592), .B1(
        \REGISTERS[10][17] ), .B2(n41), .ZN(n1286) );
  AOI22_X1 U1407 ( .A1(\REGISTERS[19][17] ), .A2(n1604), .B1(
        \REGISTERS[8][17] ), .B2(n38), .ZN(n1285) );
  NAND4_X1 U1408 ( .A1(n1288), .A2(n1287), .A3(n1286), .A4(n1285), .ZN(n1299)
         );
  AOI22_X1 U1409 ( .A1(\REGISTERS[17][17] ), .A2(n1594), .B1(
        \REGISTERS[9][17] ), .B2(n42), .ZN(n1292) );
  AOI22_X1 U1410 ( .A1(\REGISTERS[2][17] ), .A2(n1588), .B1(
        \REGISTERS[23][17] ), .B2(n48), .ZN(n1291) );
  AOI22_X1 U1411 ( .A1(\REGISTERS[18][17] ), .A2(n1605), .B1(
        \REGISTERS[7][17] ), .B2(n43), .ZN(n1290) );
  AOI22_X1 U1412 ( .A1(\REGISTERS[15][17] ), .A2(n1601), .B1(
        \REGISTERS[13][17] ), .B2(n45), .ZN(n1289) );
  NAND4_X1 U1413 ( .A1(n1292), .A2(n1291), .A3(n1290), .A4(n1289), .ZN(n1298)
         );
  AOI22_X1 U1414 ( .A1(\REGISTERS[26][17] ), .A2(n1603), .B1(
        \REGISTERS[11][17] ), .B2(n49), .ZN(n1296) );
  AOI22_X1 U1415 ( .A1(\REGISTERS[22][17] ), .A2(n51), .B1(\REGISTERS[4][17] ), 
        .B2(n37), .ZN(n1295) );
  AOI22_X1 U1416 ( .A1(\REGISTERS[20][17] ), .A2(n1616), .B1(
        \REGISTERS[12][17] ), .B2(n56), .ZN(n1294) );
  AOI22_X1 U1417 ( .A1(\REGISTERS[31][17] ), .A2(n1600), .B1(
        \REGISTERS[30][17] ), .B2(n65), .ZN(n1293) );
  NAND4_X1 U1418 ( .A1(n1296), .A2(n1295), .A3(n1294), .A4(n1293), .ZN(n1297)
         );
  NOR4_X1 U1419 ( .A1(n1300), .A2(n1299), .A3(n1298), .A4(n1297), .ZN(n1301)
         );
  AOI22_X1 U1420 ( .A1(n69), .A2(n2667), .B1(n1301), .B2(n71), .ZN(N396) );
  AOI22_X1 U1421 ( .A1(\REGISTERS[30][18] ), .A2(n1615), .B1(
        \REGISTERS[20][18] ), .B2(n66), .ZN(n1305) );
  AOI22_X1 U1422 ( .A1(\REGISTERS[21][18] ), .A2(n1599), .B1(
        \REGISTERS[4][18] ), .B2(n1575), .ZN(n1304) );
  AOI22_X1 U1423 ( .A1(\REGISTERS[17][18] ), .A2(n1594), .B1(
        \REGISTERS[18][18] ), .B2(n59), .ZN(n1303) );
  AOI22_X1 U1424 ( .A1(\REGISTERS[11][18] ), .A2(n1591), .B1(
        \REGISTERS[3][18] ), .B2(n50), .ZN(n1302) );
  NAND4_X1 U1425 ( .A1(n1305), .A2(n1304), .A3(n1303), .A4(n1302), .ZN(n1321)
         );
  AOI22_X1 U1426 ( .A1(\REGISTERS[14][18] ), .A2(n1582), .B1(
        \REGISTERS[16][18] ), .B2(n63), .ZN(n1309) );
  AOI22_X1 U1427 ( .A1(\REGISTERS[12][18] ), .A2(n1602), .B1(
        \REGISTERS[15][18] ), .B2(n55), .ZN(n1308) );
  AOI22_X1 U1428 ( .A1(\REGISTERS[24][18] ), .A2(n1589), .B1(
        \REGISTERS[25][18] ), .B2(n61), .ZN(n1307) );
  AOI22_X1 U1429 ( .A1(\REGISTERS[22][18] ), .A2(n51), .B1(\REGISTERS[23][18] ), .B2(n48), .ZN(n1306) );
  NAND4_X1 U1430 ( .A1(n1309), .A2(n1308), .A3(n1307), .A4(n1306), .ZN(n1320)
         );
  AOI22_X1 U1431 ( .A1(\REGISTERS[9][18] ), .A2(n1580), .B1(\REGISTERS[7][18] ), .B2(n43), .ZN(n1313) );
  AOI22_X1 U1432 ( .A1(\REGISTERS[0][18] ), .A2(n1614), .B1(
        \REGISTERS[27][18] ), .B2(n40), .ZN(n1312) );
  AOI22_X1 U1433 ( .A1(\REGISTERS[13][18] ), .A2(n1587), .B1(
        \REGISTERS[31][18] ), .B2(n54), .ZN(n1311) );
  AOI22_X1 U1434 ( .A1(\REGISTERS[28][18] ), .A2(n1606), .B1(
        \REGISTERS[2][18] ), .B2(n46), .ZN(n1310) );
  NAND4_X1 U1435 ( .A1(n1313), .A2(n1312), .A3(n1311), .A4(n1310), .ZN(n1319)
         );
  AOI22_X1 U1436 ( .A1(\REGISTERS[19][18] ), .A2(n1604), .B1(
        \REGISTERS[26][18] ), .B2(n57), .ZN(n1317) );
  AOI22_X1 U1437 ( .A1(\REGISTERS[29][18] ), .A2(n68), .B1(\REGISTERS[8][18] ), 
        .B2(n38), .ZN(n1316) );
  AOI22_X1 U1438 ( .A1(\REGISTERS[6][18] ), .A2(n1617), .B1(\REGISTERS[5][18] ), .B2(n62), .ZN(n1315) );
  AOI22_X1 U1439 ( .A1(\REGISTERS[10][18] ), .A2(n1579), .B1(
        \REGISTERS[1][18] ), .B2(n39), .ZN(n1314) );
  NAND4_X1 U1440 ( .A1(n1317), .A2(n1316), .A3(n1315), .A4(n1314), .ZN(n1318)
         );
  NOR4_X1 U1441 ( .A1(n1321), .A2(n1320), .A3(n1319), .A4(n1318), .ZN(n1322)
         );
  AOI22_X1 U1442 ( .A1(n69), .A2(n100), .B1(n1322), .B2(n72), .ZN(N397) );
  AOI22_X1 U1443 ( .A1(\REGISTERS[25][19] ), .A2(n61), .B1(\REGISTERS[10][19] ), .B2(n41), .ZN(n1326) );
  AOI22_X1 U1444 ( .A1(\REGISTERS[8][19] ), .A2(n1576), .B1(
        \REGISTERS[29][19] ), .B2(n68), .ZN(n1325) );
  AOI22_X1 U1445 ( .A1(\REGISTERS[20][19] ), .A2(n1616), .B1(
        \REGISTERS[2][19] ), .B2(n46), .ZN(n1324) );
  AOI22_X1 U1446 ( .A1(\REGISTERS[19][19] ), .A2(n1604), .B1(
        \REGISTERS[17][19] ), .B2(n52), .ZN(n1323) );
  NAND4_X1 U1447 ( .A1(n1326), .A2(n1325), .A3(n1324), .A4(n1323), .ZN(n1342)
         );
  AOI22_X1 U1448 ( .A1(\REGISTERS[9][19] ), .A2(n1580), .B1(\REGISTERS[0][19] ), .B2(n64), .ZN(n1330) );
  AOI22_X1 U1449 ( .A1(\REGISTERS[5][19] ), .A2(n1612), .B1(
        \REGISTERS[28][19] ), .B2(n60), .ZN(n1329) );
  AOI22_X1 U1450 ( .A1(\REGISTERS[21][19] ), .A2(n53), .B1(\REGISTERS[6][19] ), 
        .B2(n67), .ZN(n1328) );
  AOI22_X1 U1451 ( .A1(\REGISTERS[12][19] ), .A2(n56), .B1(\REGISTERS[16][19] ), .B2(n63), .ZN(n1327) );
  NAND4_X1 U1452 ( .A1(n1330), .A2(n1329), .A3(n1328), .A4(n1327), .ZN(n1341)
         );
  AOI22_X1 U1453 ( .A1(\REGISTERS[7][19] ), .A2(n43), .B1(\REGISTERS[24][19] ), 
        .B2(n47), .ZN(n1334) );
  AOI22_X1 U1454 ( .A1(\REGISTERS[14][19] ), .A2(n44), .B1(\REGISTERS[15][19] ), .B2(n55), .ZN(n1333) );
  AOI22_X1 U1455 ( .A1(\REGISTERS[18][19] ), .A2(n1605), .B1(
        \REGISTERS[3][19] ), .B2(n50), .ZN(n1332) );
  AOI22_X1 U1456 ( .A1(\REGISTERS[1][19] ), .A2(n1577), .B1(
        \REGISTERS[13][19] ), .B2(n45), .ZN(n1331) );
  NAND4_X1 U1457 ( .A1(n1334), .A2(n1333), .A3(n1332), .A4(n1331), .ZN(n1340)
         );
  AOI22_X1 U1458 ( .A1(\REGISTERS[30][19] ), .A2(n1615), .B1(
        \REGISTERS[4][19] ), .B2(n1575), .ZN(n1338) );
  AOI22_X1 U1459 ( .A1(\REGISTERS[22][19] ), .A2(n51), .B1(\REGISTERS[23][19] ), .B2(n48), .ZN(n1337) );
  AOI22_X1 U1460 ( .A1(\REGISTERS[11][19] ), .A2(n1591), .B1(
        \REGISTERS[31][19] ), .B2(n54), .ZN(n1336) );
  AOI22_X1 U1461 ( .A1(\REGISTERS[27][19] ), .A2(n1578), .B1(
        \REGISTERS[26][19] ), .B2(n57), .ZN(n1335) );
  NAND4_X1 U1462 ( .A1(n1338), .A2(n1337), .A3(n1336), .A4(n1335), .ZN(n1339)
         );
  NOR4_X1 U1463 ( .A1(n1342), .A2(n1341), .A3(n1340), .A4(n1339), .ZN(n1343)
         );
  AOI22_X1 U1464 ( .A1(n69), .A2(n2673), .B1(n1343), .B2(n72), .ZN(N398) );
  AOI22_X1 U1465 ( .A1(\REGISTERS[29][20] ), .A2(n1618), .B1(
        \REGISTERS[3][20] ), .B2(n50), .ZN(n1347) );
  AOI22_X1 U1466 ( .A1(\REGISTERS[20][20] ), .A2(n1616), .B1(
        \REGISTERS[31][20] ), .B2(n54), .ZN(n1346) );
  AOI22_X1 U1467 ( .A1(\REGISTERS[6][20] ), .A2(n1617), .B1(\REGISTERS[4][20] ), .B2(n37), .ZN(n1345) );
  AOI22_X1 U1468 ( .A1(\REGISTERS[2][20] ), .A2(n1588), .B1(
        \REGISTERS[16][20] ), .B2(n63), .ZN(n1344) );
  NAND4_X1 U1469 ( .A1(n1347), .A2(n1346), .A3(n1345), .A4(n1344), .ZN(n1363)
         );
  AOI22_X1 U1470 ( .A1(\REGISTERS[21][20] ), .A2(n1599), .B1(
        \REGISTERS[28][20] ), .B2(n60), .ZN(n1351) );
  AOI22_X1 U1471 ( .A1(\REGISTERS[10][20] ), .A2(n1579), .B1(
        \REGISTERS[8][20] ), .B2(n38), .ZN(n1350) );
  AOI22_X1 U1472 ( .A1(\REGISTERS[23][20] ), .A2(n1590), .B1(
        \REGISTERS[13][20] ), .B2(n45), .ZN(n1349) );
  AOI22_X1 U1473 ( .A1(\REGISTERS[26][20] ), .A2(n1603), .B1(
        \REGISTERS[25][20] ), .B2(n61), .ZN(n1348) );
  NAND4_X1 U1474 ( .A1(n1351), .A2(n1350), .A3(n1349), .A4(n1348), .ZN(n1362)
         );
  AOI22_X1 U1475 ( .A1(\REGISTERS[27][20] ), .A2(n1578), .B1(
        \REGISTERS[7][20] ), .B2(n43), .ZN(n1355) );
  AOI22_X1 U1476 ( .A1(\REGISTERS[19][20] ), .A2(n1604), .B1(
        \REGISTERS[9][20] ), .B2(n42), .ZN(n1354) );
  AOI22_X1 U1477 ( .A1(\REGISTERS[18][20] ), .A2(n1605), .B1(
        \REGISTERS[24][20] ), .B2(n47), .ZN(n1353) );
  AOI22_X1 U1478 ( .A1(\REGISTERS[30][20] ), .A2(n1615), .B1(
        \REGISTERS[12][20] ), .B2(n56), .ZN(n1352) );
  NAND4_X1 U1479 ( .A1(n1355), .A2(n1354), .A3(n1353), .A4(n1352), .ZN(n1361)
         );
  AOI22_X1 U1480 ( .A1(\REGISTERS[11][20] ), .A2(n1591), .B1(
        \REGISTERS[15][20] ), .B2(n55), .ZN(n1359) );
  AOI22_X1 U1481 ( .A1(\REGISTERS[17][20] ), .A2(n1594), .B1(
        \REGISTERS[5][20] ), .B2(n62), .ZN(n1358) );
  AOI22_X1 U1482 ( .A1(\REGISTERS[1][20] ), .A2(n1577), .B1(
        \REGISTERS[14][20] ), .B2(n44), .ZN(n1357) );
  AOI22_X1 U1483 ( .A1(\REGISTERS[22][20] ), .A2(n51), .B1(\REGISTERS[0][20] ), 
        .B2(n64), .ZN(n1356) );
  NAND4_X1 U1484 ( .A1(n1359), .A2(n1358), .A3(n1357), .A4(n1356), .ZN(n1360)
         );
  NOR4_X1 U1485 ( .A1(n1363), .A2(n1362), .A3(n1361), .A4(n1360), .ZN(n1364)
         );
  AOI22_X1 U1486 ( .A1(n69), .A2(n96), .B1(n1364), .B2(n71), .ZN(N399) );
  AOI22_X1 U1487 ( .A1(\REGISTERS[12][21] ), .A2(n1602), .B1(
        \REGISTERS[26][21] ), .B2(n57), .ZN(n1368) );
  AOI22_X1 U1488 ( .A1(\REGISTERS[22][21] ), .A2(n1593), .B1(
        \REGISTERS[20][21] ), .B2(n66), .ZN(n1367) );
  AOI22_X1 U1489 ( .A1(\REGISTERS[5][21] ), .A2(n1612), .B1(
        \REGISTERS[16][21] ), .B2(n63), .ZN(n1366) );
  AOI22_X1 U1490 ( .A1(\REGISTERS[28][21] ), .A2(n60), .B1(\REGISTERS[27][21] ), .B2(n40), .ZN(n1365) );
  NAND4_X1 U1491 ( .A1(n1368), .A2(n1367), .A3(n1366), .A4(n1365), .ZN(n1384)
         );
  AOI22_X1 U1492 ( .A1(\REGISTERS[0][21] ), .A2(n1614), .B1(\REGISTERS[6][21] ), .B2(n67), .ZN(n1372) );
  AOI22_X1 U1493 ( .A1(\REGISTERS[9][21] ), .A2(n1580), .B1(\REGISTERS[8][21] ), .B2(n1576), .ZN(n1371) );
  AOI22_X1 U1494 ( .A1(\REGISTERS[3][21] ), .A2(n1592), .B1(
        \REGISTERS[30][21] ), .B2(n65), .ZN(n1370) );
  AOI22_X1 U1495 ( .A1(\REGISTERS[2][21] ), .A2(n46), .B1(\REGISTERS[24][21] ), 
        .B2(n47), .ZN(n1369) );
  NAND4_X1 U1496 ( .A1(n1372), .A2(n1371), .A3(n1370), .A4(n1369), .ZN(n1383)
         );
  AOI22_X1 U1497 ( .A1(\REGISTERS[29][21] ), .A2(n68), .B1(\REGISTERS[15][21] ), .B2(n55), .ZN(n1376) );
  AOI22_X1 U1498 ( .A1(\REGISTERS[19][21] ), .A2(n1604), .B1(
        \REGISTERS[11][21] ), .B2(n49), .ZN(n1375) );
  AOI22_X1 U1499 ( .A1(\REGISTERS[1][21] ), .A2(n1577), .B1(
        \REGISTERS[13][21] ), .B2(n45), .ZN(n1374) );
  AOI22_X1 U1500 ( .A1(\REGISTERS[10][21] ), .A2(n1579), .B1(
        \REGISTERS[18][21] ), .B2(n59), .ZN(n1373) );
  NAND4_X1 U1501 ( .A1(n1376), .A2(n1375), .A3(n1374), .A4(n1373), .ZN(n1382)
         );
  AOI22_X1 U1502 ( .A1(\REGISTERS[21][21] ), .A2(n1599), .B1(
        \REGISTERS[4][21] ), .B2(n37), .ZN(n1380) );
  AOI22_X1 U1503 ( .A1(\REGISTERS[14][21] ), .A2(n1582), .B1(
        \REGISTERS[17][21] ), .B2(n52), .ZN(n1379) );
  AOI22_X1 U1504 ( .A1(\REGISTERS[7][21] ), .A2(n1581), .B1(
        \REGISTERS[25][21] ), .B2(n61), .ZN(n1378) );
  AOI22_X1 U1505 ( .A1(\REGISTERS[31][21] ), .A2(n54), .B1(\REGISTERS[23][21] ), .B2(n48), .ZN(n1377) );
  NAND4_X1 U1506 ( .A1(n1380), .A2(n1379), .A3(n1378), .A4(n1377), .ZN(n1381)
         );
  NOR4_X1 U1507 ( .A1(n1384), .A2(n1383), .A3(n1382), .A4(n1381), .ZN(n1385)
         );
  AOI22_X1 U1508 ( .A1(n69), .A2(n94), .B1(n1385), .B2(n72), .ZN(N400) );
  AOI22_X1 U1509 ( .A1(\REGISTERS[13][22] ), .A2(n45), .B1(\REGISTERS[22][22] ), .B2(n51), .ZN(n1389) );
  AOI22_X1 U1510 ( .A1(\REGISTERS[9][22] ), .A2(n42), .B1(\REGISTERS[1][22] ), 
        .B2(n39), .ZN(n1388) );
  AOI22_X1 U1511 ( .A1(\REGISTERS[31][22] ), .A2(n1600), .B1(
        \REGISTERS[4][22] ), .B2(n37), .ZN(n1387) );
  AOI22_X1 U1512 ( .A1(\REGISTERS[27][22] ), .A2(n40), .B1(\REGISTERS[20][22] ), .B2(n66), .ZN(n1386) );
  NAND4_X1 U1513 ( .A1(n1389), .A2(n1388), .A3(n1387), .A4(n1386), .ZN(n1405)
         );
  AOI22_X1 U1514 ( .A1(\REGISTERS[23][22] ), .A2(n1590), .B1(
        \REGISTERS[25][22] ), .B2(n61), .ZN(n1393) );
  AOI22_X1 U1515 ( .A1(\REGISTERS[21][22] ), .A2(n53), .B1(\REGISTERS[11][22] ), .B2(n49), .ZN(n1392) );
  AOI22_X1 U1516 ( .A1(\REGISTERS[3][22] ), .A2(n1592), .B1(
        \REGISTERS[28][22] ), .B2(n60), .ZN(n1391) );
  AOI22_X1 U1517 ( .A1(\REGISTERS[12][22] ), .A2(n1602), .B1(
        \REGISTERS[29][22] ), .B2(n68), .ZN(n1390) );
  NAND4_X1 U1518 ( .A1(n1393), .A2(n1392), .A3(n1391), .A4(n1390), .ZN(n1404)
         );
  AOI22_X1 U1519 ( .A1(\REGISTERS[24][22] ), .A2(n1589), .B1(
        \REGISTERS[14][22] ), .B2(n44), .ZN(n1397) );
  AOI22_X1 U1520 ( .A1(\REGISTERS[18][22] ), .A2(n59), .B1(\REGISTERS[8][22] ), 
        .B2(n1576), .ZN(n1396) );
  AOI22_X1 U1521 ( .A1(\REGISTERS[6][22] ), .A2(n1617), .B1(
        \REGISTERS[19][22] ), .B2(n58), .ZN(n1395) );
  AOI22_X1 U1522 ( .A1(\REGISTERS[5][22] ), .A2(n62), .B1(\REGISTERS[16][22] ), 
        .B2(n63), .ZN(n1394) );
  NAND4_X1 U1523 ( .A1(n1397), .A2(n1396), .A3(n1395), .A4(n1394), .ZN(n1403)
         );
  AOI22_X1 U1524 ( .A1(\REGISTERS[2][22] ), .A2(n1588), .B1(
        \REGISTERS[15][22] ), .B2(n55), .ZN(n1401) );
  AOI22_X1 U1525 ( .A1(\REGISTERS[10][22] ), .A2(n41), .B1(\REGISTERS[30][22] ), .B2(n65), .ZN(n1400) );
  AOI22_X1 U1526 ( .A1(\REGISTERS[7][22] ), .A2(n43), .B1(\REGISTERS[17][22] ), 
        .B2(n52), .ZN(n1399) );
  AOI22_X1 U1527 ( .A1(\REGISTERS[26][22] ), .A2(n1603), .B1(
        \REGISTERS[0][22] ), .B2(n64), .ZN(n1398) );
  NAND4_X1 U1528 ( .A1(n1401), .A2(n1400), .A3(n1399), .A4(n1398), .ZN(n1402)
         );
  NOR4_X1 U1529 ( .A1(n1405), .A2(n1404), .A3(n1403), .A4(n1402), .ZN(n1406)
         );
  AOI22_X1 U1530 ( .A1(n69), .A2(n2672), .B1(n1406), .B2(n72), .ZN(N401) );
  AOI22_X1 U1531 ( .A1(\REGISTERS[14][23] ), .A2(n44), .B1(\REGISTERS[4][23] ), 
        .B2(n37), .ZN(n1410) );
  AOI22_X1 U1532 ( .A1(\REGISTERS[2][23] ), .A2(n46), .B1(\REGISTERS[10][23] ), 
        .B2(n41), .ZN(n1409) );
  AOI22_X1 U1533 ( .A1(\REGISTERS[20][23] ), .A2(n1616), .B1(
        \REGISTERS[1][23] ), .B2(n39), .ZN(n1408) );
  AOI22_X1 U1534 ( .A1(\REGISTERS[6][23] ), .A2(n1617), .B1(
        \REGISTERS[17][23] ), .B2(n52), .ZN(n1407) );
  NAND4_X1 U1535 ( .A1(n1410), .A2(n1409), .A3(n1408), .A4(n1407), .ZN(n1426)
         );
  AOI22_X1 U1536 ( .A1(\REGISTERS[18][23] ), .A2(n1605), .B1(
        \REGISTERS[3][23] ), .B2(n50), .ZN(n1414) );
  AOI22_X1 U1537 ( .A1(\REGISTERS[19][23] ), .A2(n1604), .B1(
        \REGISTERS[29][23] ), .B2(n68), .ZN(n1413) );
  AOI22_X1 U1538 ( .A1(\REGISTERS[16][23] ), .A2(n1613), .B1(
        \REGISTERS[30][23] ), .B2(n65), .ZN(n1412) );
  AOI22_X1 U1539 ( .A1(\REGISTERS[27][23] ), .A2(n1578), .B1(
        \REGISTERS[21][23] ), .B2(n53), .ZN(n1411) );
  NAND4_X1 U1540 ( .A1(n1414), .A2(n1413), .A3(n1412), .A4(n1411), .ZN(n1425)
         );
  AOI22_X1 U1541 ( .A1(\REGISTERS[9][23] ), .A2(n1580), .B1(
        \REGISTERS[31][23] ), .B2(n54), .ZN(n1418) );
  AOI22_X1 U1542 ( .A1(\REGISTERS[22][23] ), .A2(n1593), .B1(
        \REGISTERS[12][23] ), .B2(n56), .ZN(n1417) );
  AOI22_X1 U1543 ( .A1(\REGISTERS[0][23] ), .A2(n64), .B1(\REGISTERS[24][23] ), 
        .B2(n47), .ZN(n1416) );
  AOI22_X1 U1544 ( .A1(\REGISTERS[5][23] ), .A2(n62), .B1(\REGISTERS[11][23] ), 
        .B2(n49), .ZN(n1415) );
  NAND4_X1 U1545 ( .A1(n1418), .A2(n1417), .A3(n1416), .A4(n1415), .ZN(n1424)
         );
  AOI22_X1 U1546 ( .A1(\REGISTERS[28][23] ), .A2(n1606), .B1(
        \REGISTERS[15][23] ), .B2(n55), .ZN(n1422) );
  AOI22_X1 U1547 ( .A1(\REGISTERS[8][23] ), .A2(n38), .B1(\REGISTERS[23][23] ), 
        .B2(n48), .ZN(n1421) );
  AOI22_X1 U1548 ( .A1(\REGISTERS[26][23] ), .A2(n1603), .B1(
        \REGISTERS[13][23] ), .B2(n45), .ZN(n1420) );
  AOI22_X1 U1549 ( .A1(\REGISTERS[7][23] ), .A2(n1581), .B1(
        \REGISTERS[25][23] ), .B2(n61), .ZN(n1419) );
  NAND4_X1 U1550 ( .A1(n1422), .A2(n1421), .A3(n1420), .A4(n1419), .ZN(n1423)
         );
  NOR4_X1 U1551 ( .A1(n1426), .A2(n1425), .A3(n1424), .A4(n1423), .ZN(n1427)
         );
  AOI22_X1 U1552 ( .A1(n69), .A2(n90), .B1(n1427), .B2(n72), .ZN(N402) );
  AOI22_X1 U1553 ( .A1(\REGISTERS[8][24] ), .A2(n1576), .B1(\REGISTERS[4][24] ), .B2(n37), .ZN(n1431) );
  AOI22_X1 U1554 ( .A1(\REGISTERS[5][24] ), .A2(n62), .B1(\REGISTERS[1][24] ), 
        .B2(n39), .ZN(n1430) );
  AOI22_X1 U1555 ( .A1(\REGISTERS[25][24] ), .A2(n1611), .B1(
        \REGISTERS[20][24] ), .B2(n66), .ZN(n1429) );
  AOI22_X1 U1556 ( .A1(\REGISTERS[22][24] ), .A2(n1593), .B1(
        \REGISTERS[24][24] ), .B2(n47), .ZN(n1428) );
  NAND4_X1 U1557 ( .A1(n1431), .A2(n1430), .A3(n1429), .A4(n1428), .ZN(n1447)
         );
  AOI22_X1 U1558 ( .A1(\REGISTERS[0][24] ), .A2(n1614), .B1(
        \REGISTERS[28][24] ), .B2(n60), .ZN(n1435) );
  AOI22_X1 U1559 ( .A1(\REGISTERS[19][24] ), .A2(n1604), .B1(
        \REGISTERS[11][24] ), .B2(n49), .ZN(n1434) );
  AOI22_X1 U1560 ( .A1(\REGISTERS[12][24] ), .A2(n1602), .B1(
        \REGISTERS[9][24] ), .B2(n42), .ZN(n1433) );
  AOI22_X1 U1561 ( .A1(\REGISTERS[17][24] ), .A2(n52), .B1(\REGISTERS[21][24] ), .B2(n53), .ZN(n1432) );
  NAND4_X1 U1562 ( .A1(n1435), .A2(n1434), .A3(n1433), .A4(n1432), .ZN(n1446)
         );
  AOI22_X1 U1563 ( .A1(\REGISTERS[27][24] ), .A2(n40), .B1(\REGISTERS[3][24] ), 
        .B2(n50), .ZN(n1439) );
  AOI22_X1 U1564 ( .A1(\REGISTERS[16][24] ), .A2(n1613), .B1(
        \REGISTERS[15][24] ), .B2(n55), .ZN(n1438) );
  AOI22_X1 U1565 ( .A1(\REGISTERS[29][24] ), .A2(n1618), .B1(
        \REGISTERS[6][24] ), .B2(n67), .ZN(n1437) );
  AOI22_X1 U1566 ( .A1(\REGISTERS[30][24] ), .A2(n65), .B1(\REGISTERS[18][24] ), .B2(n59), .ZN(n1436) );
  NAND4_X1 U1567 ( .A1(n1439), .A2(n1438), .A3(n1437), .A4(n1436), .ZN(n1445)
         );
  AOI22_X1 U1568 ( .A1(\REGISTERS[14][24] ), .A2(n1582), .B1(
        \REGISTERS[7][24] ), .B2(n43), .ZN(n1443) );
  AOI22_X1 U1569 ( .A1(\REGISTERS[26][24] ), .A2(n57), .B1(\REGISTERS[13][24] ), .B2(n45), .ZN(n1442) );
  AOI22_X1 U1570 ( .A1(\REGISTERS[2][24] ), .A2(n46), .B1(\REGISTERS[31][24] ), 
        .B2(n54), .ZN(n1441) );
  AOI22_X1 U1571 ( .A1(\REGISTERS[10][24] ), .A2(n41), .B1(\REGISTERS[23][24] ), .B2(n48), .ZN(n1440) );
  NAND4_X1 U1572 ( .A1(n1443), .A2(n1442), .A3(n1441), .A4(n1440), .ZN(n1444)
         );
  NOR4_X1 U1573 ( .A1(n1447), .A2(n1446), .A3(n1445), .A4(n1444), .ZN(n1448)
         );
  AOI22_X1 U1574 ( .A1(n70), .A2(n88), .B1(n1448), .B2(n72), .ZN(N403) );
  AOI22_X1 U1575 ( .A1(\REGISTERS[14][25] ), .A2(n44), .B1(\REGISTERS[22][25] ), .B2(n51), .ZN(n1452) );
  AOI22_X1 U1576 ( .A1(\REGISTERS[23][25] ), .A2(n1590), .B1(
        \REGISTERS[29][25] ), .B2(n68), .ZN(n1451) );
  AOI22_X1 U1577 ( .A1(\REGISTERS[27][25] ), .A2(n1578), .B1(
        \REGISTERS[4][25] ), .B2(n37), .ZN(n1450) );
  AOI22_X1 U1578 ( .A1(\REGISTERS[24][25] ), .A2(n1589), .B1(
        \REGISTERS[10][25] ), .B2(n41), .ZN(n1449) );
  NAND4_X1 U1579 ( .A1(n1452), .A2(n1451), .A3(n1450), .A4(n1449), .ZN(n1468)
         );
  AOI22_X1 U1580 ( .A1(\REGISTERS[25][25] ), .A2(n61), .B1(\REGISTERS[1][25] ), 
        .B2(n39), .ZN(n1456) );
  AOI22_X1 U1581 ( .A1(\REGISTERS[26][25] ), .A2(n1603), .B1(
        \REGISTERS[0][25] ), .B2(n64), .ZN(n1455) );
  AOI22_X1 U1582 ( .A1(\REGISTERS[18][25] ), .A2(n59), .B1(\REGISTERS[9][25] ), 
        .B2(n42), .ZN(n1454) );
  AOI22_X1 U1583 ( .A1(\REGISTERS[3][25] ), .A2(n50), .B1(\REGISTERS[6][25] ), 
        .B2(n67), .ZN(n1453) );
  NAND4_X1 U1584 ( .A1(n1456), .A2(n1455), .A3(n1454), .A4(n1453), .ZN(n1467)
         );
  AOI22_X1 U1585 ( .A1(\REGISTERS[8][25] ), .A2(n38), .B1(\REGISTERS[12][25] ), 
        .B2(n56), .ZN(n1460) );
  AOI22_X1 U1586 ( .A1(\REGISTERS[17][25] ), .A2(n1594), .B1(
        \REGISTERS[16][25] ), .B2(n63), .ZN(n1459) );
  AOI22_X1 U1587 ( .A1(\REGISTERS[11][25] ), .A2(n1591), .B1(
        \REGISTERS[31][25] ), .B2(n54), .ZN(n1458) );
  AOI22_X1 U1588 ( .A1(\REGISTERS[2][25] ), .A2(n46), .B1(\REGISTERS[13][25] ), 
        .B2(n45), .ZN(n1457) );
  NAND4_X1 U1589 ( .A1(n1460), .A2(n1459), .A3(n1458), .A4(n1457), .ZN(n1466)
         );
  AOI22_X1 U1590 ( .A1(\REGISTERS[19][25] ), .A2(n58), .B1(\REGISTERS[7][25] ), 
        .B2(n43), .ZN(n1464) );
  AOI22_X1 U1591 ( .A1(\REGISTERS[5][25] ), .A2(n1612), .B1(
        \REGISTERS[28][25] ), .B2(n60), .ZN(n1463) );
  AOI22_X1 U1592 ( .A1(\REGISTERS[30][25] ), .A2(n1615), .B1(
        \REGISTERS[15][25] ), .B2(n55), .ZN(n1462) );
  AOI22_X1 U1593 ( .A1(\REGISTERS[20][25] ), .A2(n66), .B1(\REGISTERS[21][25] ), .B2(n53), .ZN(n1461) );
  NAND4_X1 U1594 ( .A1(n1464), .A2(n1463), .A3(n1462), .A4(n1461), .ZN(n1465)
         );
  NOR4_X1 U1595 ( .A1(n1468), .A2(n1467), .A3(n1466), .A4(n1465), .ZN(n1469)
         );
  AOI22_X1 U1596 ( .A1(n70), .A2(n86), .B1(n1469), .B2(n71), .ZN(N404) );
  AOI22_X1 U1597 ( .A1(\REGISTERS[12][26] ), .A2(n56), .B1(\REGISTERS[10][26] ), .B2(n41), .ZN(n1473) );
  AOI22_X1 U1598 ( .A1(\REGISTERS[15][26] ), .A2(n1601), .B1(
        \REGISTERS[0][26] ), .B2(n64), .ZN(n1472) );
  AOI22_X1 U1599 ( .A1(\REGISTERS[1][26] ), .A2(n39), .B1(\REGISTERS[4][26] ), 
        .B2(n37), .ZN(n1471) );
  AOI22_X1 U1600 ( .A1(\REGISTERS[28][26] ), .A2(n60), .B1(\REGISTERS[23][26] ), .B2(n48), .ZN(n1470) );
  NAND4_X1 U1601 ( .A1(n1473), .A2(n1472), .A3(n1471), .A4(n1470), .ZN(n1489)
         );
  AOI22_X1 U1602 ( .A1(\REGISTERS[22][26] ), .A2(n1593), .B1(
        \REGISTERS[6][26] ), .B2(n67), .ZN(n1477) );
  AOI22_X1 U1603 ( .A1(\REGISTERS[25][26] ), .A2(n1611), .B1(
        \REGISTERS[27][26] ), .B2(n40), .ZN(n1476) );
  AOI22_X1 U1604 ( .A1(\REGISTERS[19][26] ), .A2(n1604), .B1(
        \REGISTERS[17][26] ), .B2(n52), .ZN(n1475) );
  AOI22_X1 U1605 ( .A1(\REGISTERS[24][26] ), .A2(n1589), .B1(
        \REGISTERS[30][26] ), .B2(n65), .ZN(n1474) );
  NAND4_X1 U1606 ( .A1(n1477), .A2(n1476), .A3(n1475), .A4(n1474), .ZN(n1488)
         );
  AOI22_X1 U1607 ( .A1(\REGISTERS[16][26] ), .A2(n1613), .B1(
        \REGISTERS[11][26] ), .B2(n49), .ZN(n1481) );
  AOI22_X1 U1608 ( .A1(\REGISTERS[3][26] ), .A2(n1592), .B1(
        \REGISTERS[18][26] ), .B2(n59), .ZN(n1480) );
  AOI22_X1 U1609 ( .A1(\REGISTERS[9][26] ), .A2(n42), .B1(\REGISTERS[7][26] ), 
        .B2(n43), .ZN(n1479) );
  AOI22_X1 U1610 ( .A1(\REGISTERS[31][26] ), .A2(n54), .B1(\REGISTERS[14][26] ), .B2(n44), .ZN(n1478) );
  NAND4_X1 U1611 ( .A1(n1481), .A2(n1480), .A3(n1479), .A4(n1478), .ZN(n1487)
         );
  AOI22_X1 U1612 ( .A1(\REGISTERS[21][26] ), .A2(n53), .B1(\REGISTERS[8][26] ), 
        .B2(n38), .ZN(n1485) );
  AOI22_X1 U1613 ( .A1(\REGISTERS[20][26] ), .A2(n1616), .B1(
        \REGISTERS[2][26] ), .B2(n46), .ZN(n1484) );
  AOI22_X1 U1614 ( .A1(\REGISTERS[13][26] ), .A2(n1587), .B1(
        \REGISTERS[5][26] ), .B2(n62), .ZN(n1483) );
  AOI22_X1 U1615 ( .A1(\REGISTERS[29][26] ), .A2(n68), .B1(\REGISTERS[26][26] ), .B2(n57), .ZN(n1482) );
  NAND4_X1 U1616 ( .A1(n1485), .A2(n1484), .A3(n1483), .A4(n1482), .ZN(n1486)
         );
  NOR4_X1 U1617 ( .A1(n1489), .A2(n1488), .A3(n1487), .A4(n1486), .ZN(n1490)
         );
  AOI22_X1 U1618 ( .A1(n70), .A2(n84), .B1(n1490), .B2(n71), .ZN(N405) );
  AOI22_X1 U1619 ( .A1(\REGISTERS[26][27] ), .A2(n57), .B1(\REGISTERS[7][27] ), 
        .B2(n43), .ZN(n1494) );
  AOI22_X1 U1620 ( .A1(\REGISTERS[9][27] ), .A2(n1580), .B1(
        \REGISTERS[20][27] ), .B2(n66), .ZN(n1493) );
  AOI22_X1 U1621 ( .A1(\REGISTERS[18][27] ), .A2(n1605), .B1(
        \REGISTERS[27][27] ), .B2(n40), .ZN(n1492) );
  AOI22_X1 U1622 ( .A1(\REGISTERS[31][27] ), .A2(n1600), .B1(
        \REGISTERS[0][27] ), .B2(n64), .ZN(n1491) );
  NAND4_X1 U1623 ( .A1(n1494), .A2(n1493), .A3(n1492), .A4(n1491), .ZN(n1510)
         );
  AOI22_X1 U1624 ( .A1(\REGISTERS[2][27] ), .A2(n46), .B1(\REGISTERS[29][27] ), 
        .B2(n68), .ZN(n1498) );
  AOI22_X1 U1625 ( .A1(\REGISTERS[1][27] ), .A2(n1577), .B1(
        \REGISTERS[19][27] ), .B2(n58), .ZN(n1497) );
  AOI22_X1 U1626 ( .A1(\REGISTERS[5][27] ), .A2(n1612), .B1(
        \REGISTERS[22][27] ), .B2(n51), .ZN(n1496) );
  AOI22_X1 U1627 ( .A1(\REGISTERS[15][27] ), .A2(n1601), .B1(
        \REGISTERS[14][27] ), .B2(n44), .ZN(n1495) );
  NAND4_X1 U1628 ( .A1(n1498), .A2(n1497), .A3(n1496), .A4(n1495), .ZN(n1509)
         );
  AOI22_X1 U1629 ( .A1(\REGISTERS[10][27] ), .A2(n1579), .B1(
        \REGISTERS[6][27] ), .B2(n67), .ZN(n1502) );
  AOI22_X1 U1630 ( .A1(\REGISTERS[11][27] ), .A2(n1591), .B1(
        \REGISTERS[30][27] ), .B2(n65), .ZN(n1501) );
  AOI22_X1 U1631 ( .A1(\REGISTERS[3][27] ), .A2(n1592), .B1(
        \REGISTERS[25][27] ), .B2(n61), .ZN(n1500) );
  AOI22_X1 U1632 ( .A1(\REGISTERS[16][27] ), .A2(n1613), .B1(
        \REGISTERS[8][27] ), .B2(n38), .ZN(n1499) );
  NAND4_X1 U1633 ( .A1(n1502), .A2(n1501), .A3(n1500), .A4(n1499), .ZN(n1508)
         );
  AOI22_X1 U1634 ( .A1(\REGISTERS[17][27] ), .A2(n52), .B1(\REGISTERS[28][27] ), .B2(n60), .ZN(n1506) );
  AOI22_X1 U1635 ( .A1(\REGISTERS[12][27] ), .A2(n1602), .B1(
        \REGISTERS[24][27] ), .B2(n47), .ZN(n1505) );
  AOI22_X1 U1636 ( .A1(\REGISTERS[13][27] ), .A2(n45), .B1(\REGISTERS[4][27] ), 
        .B2(n37), .ZN(n1504) );
  AOI22_X1 U1637 ( .A1(\REGISTERS[23][27] ), .A2(n1590), .B1(
        \REGISTERS[21][27] ), .B2(n53), .ZN(n1503) );
  NAND4_X1 U1638 ( .A1(n1506), .A2(n1505), .A3(n1504), .A4(n1503), .ZN(n1507)
         );
  NOR4_X1 U1639 ( .A1(n1510), .A2(n1509), .A3(n1508), .A4(n1507), .ZN(n1511)
         );
  AOI22_X1 U1640 ( .A1(n70), .A2(n2657), .B1(n1511), .B2(n71), .ZN(N406) );
  AOI22_X1 U1641 ( .A1(\REGISTERS[20][28] ), .A2(n66), .B1(\REGISTERS[19][28] ), .B2(n58), .ZN(n1515) );
  AOI22_X1 U1642 ( .A1(\REGISTERS[4][28] ), .A2(n1575), .B1(
        \REGISTERS[28][28] ), .B2(n60), .ZN(n1514) );
  AOI22_X1 U1643 ( .A1(\REGISTERS[6][28] ), .A2(n1617), .B1(
        \REGISTERS[29][28] ), .B2(n68), .ZN(n1513) );
  AOI22_X1 U1644 ( .A1(\REGISTERS[21][28] ), .A2(n1599), .B1(
        \REGISTERS[30][28] ), .B2(n65), .ZN(n1512) );
  NAND4_X1 U1645 ( .A1(n1515), .A2(n1514), .A3(n1513), .A4(n1512), .ZN(n1531)
         );
  AOI22_X1 U1646 ( .A1(\REGISTERS[13][28] ), .A2(n1587), .B1(
        \REGISTERS[16][28] ), .B2(n63), .ZN(n1519) );
  AOI22_X1 U1647 ( .A1(\REGISTERS[24][28] ), .A2(n1589), .B1(
        \REGISTERS[14][28] ), .B2(n44), .ZN(n1518) );
  AOI22_X1 U1648 ( .A1(\REGISTERS[12][28] ), .A2(n56), .B1(\REGISTERS[23][28] ), .B2(n48), .ZN(n1517) );
  AOI22_X1 U1649 ( .A1(\REGISTERS[9][28] ), .A2(n42), .B1(\REGISTERS[7][28] ), 
        .B2(n43), .ZN(n1516) );
  NAND4_X1 U1650 ( .A1(n1519), .A2(n1518), .A3(n1517), .A4(n1516), .ZN(n1530)
         );
  AOI22_X1 U1651 ( .A1(\REGISTERS[18][28] ), .A2(n59), .B1(\REGISTERS[17][28] ), .B2(n52), .ZN(n1523) );
  AOI22_X1 U1652 ( .A1(\REGISTERS[8][28] ), .A2(n1576), .B1(\REGISTERS[5][28] ), .B2(n62), .ZN(n1522) );
  AOI22_X1 U1653 ( .A1(\REGISTERS[11][28] ), .A2(n1591), .B1(
        \REGISTERS[26][28] ), .B2(n57), .ZN(n1521) );
  AOI22_X1 U1654 ( .A1(\REGISTERS[15][28] ), .A2(n1601), .B1(
        \REGISTERS[3][28] ), .B2(n50), .ZN(n1520) );
  NAND4_X1 U1655 ( .A1(n1523), .A2(n1522), .A3(n1521), .A4(n1520), .ZN(n1529)
         );
  AOI22_X1 U1656 ( .A1(\REGISTERS[0][28] ), .A2(n64), .B1(\REGISTERS[10][28] ), 
        .B2(n41), .ZN(n1527) );
  AOI22_X1 U1657 ( .A1(\REGISTERS[2][28] ), .A2(n1588), .B1(\REGISTERS[1][28] ), .B2(n39), .ZN(n1526) );
  AOI22_X1 U1658 ( .A1(\REGISTERS[22][28] ), .A2(n1593), .B1(
        \REGISTERS[25][28] ), .B2(n61), .ZN(n1525) );
  AOI22_X1 U1659 ( .A1(\REGISTERS[27][28] ), .A2(n40), .B1(\REGISTERS[31][28] ), .B2(n54), .ZN(n1524) );
  NAND4_X1 U1660 ( .A1(n1527), .A2(n1526), .A3(n1525), .A4(n1524), .ZN(n1528)
         );
  NOR4_X1 U1661 ( .A1(n1531), .A2(n1530), .A3(n1529), .A4(n1528), .ZN(n1532)
         );
  AOI22_X1 U1663 ( .A1(\REGISTERS[24][29] ), .A2(n47), .B1(\REGISTERS[9][29] ), 
        .B2(n42), .ZN(n1536) );
  AOI22_X1 U1664 ( .A1(\REGISTERS[10][29] ), .A2(n41), .B1(\REGISTERS[26][29] ), .B2(n57), .ZN(n1535) );
  AOI22_X1 U1665 ( .A1(\REGISTERS[20][29] ), .A2(n1616), .B1(
        \REGISTERS[23][29] ), .B2(n48), .ZN(n1534) );
  AOI22_X1 U1666 ( .A1(\REGISTERS[8][29] ), .A2(n38), .B1(\REGISTERS[12][29] ), 
        .B2(n56), .ZN(n1533) );
  NAND4_X1 U1667 ( .A1(n1536), .A2(n1535), .A3(n1534), .A4(n1533), .ZN(n1552)
         );
  AOI22_X1 U1668 ( .A1(\REGISTERS[17][29] ), .A2(n1594), .B1(
        \REGISTERS[30][29] ), .B2(n65), .ZN(n1540) );
  AOI22_X1 U1669 ( .A1(\REGISTERS[19][29] ), .A2(n58), .B1(\REGISTERS[2][29] ), 
        .B2(n46), .ZN(n1539) );
  AOI22_X1 U1670 ( .A1(\REGISTERS[16][29] ), .A2(n63), .B1(\REGISTERS[6][29] ), 
        .B2(n67), .ZN(n1538) );
  AOI22_X1 U1671 ( .A1(\REGISTERS[3][29] ), .A2(n1592), .B1(
        \REGISTERS[14][29] ), .B2(n44), .ZN(n1537) );
  NAND4_X1 U1672 ( .A1(n1540), .A2(n1539), .A3(n1538), .A4(n1537), .ZN(n1551)
         );
  AOI22_X1 U1673 ( .A1(\REGISTERS[0][29] ), .A2(n1614), .B1(
        \REGISTERS[31][29] ), .B2(n54), .ZN(n1544) );
  AOI22_X1 U1674 ( .A1(\REGISTERS[28][29] ), .A2(n1606), .B1(
        \REGISTERS[13][29] ), .B2(n45), .ZN(n1543) );
  AOI22_X1 U1675 ( .A1(\REGISTERS[15][29] ), .A2(n55), .B1(\REGISTERS[11][29] ), .B2(n49), .ZN(n1542) );
  AOI22_X1 U1676 ( .A1(\REGISTERS[4][29] ), .A2(n1575), .B1(
        \REGISTERS[27][29] ), .B2(n40), .ZN(n1541) );
  NAND4_X1 U1677 ( .A1(n1544), .A2(n1543), .A3(n1542), .A4(n1541), .ZN(n1550)
         );
  AOI22_X1 U1678 ( .A1(\REGISTERS[25][29] ), .A2(n61), .B1(\REGISTERS[18][29] ), .B2(n59), .ZN(n1548) );
  AOI22_X1 U1679 ( .A1(\REGISTERS[22][29] ), .A2(n1593), .B1(
        \REGISTERS[29][29] ), .B2(n68), .ZN(n1547) );
  AOI22_X1 U1680 ( .A1(\REGISTERS[5][29] ), .A2(n1612), .B1(\REGISTERS[7][29] ), .B2(n43), .ZN(n1546) );
  AOI22_X1 U1681 ( .A1(\REGISTERS[1][29] ), .A2(n39), .B1(\REGISTERS[21][29] ), 
        .B2(n53), .ZN(n1545) );
  NAND4_X1 U1682 ( .A1(n1548), .A2(n1547), .A3(n1546), .A4(n1545), .ZN(n1549)
         );
  NOR4_X1 U1683 ( .A1(n1552), .A2(n1551), .A3(n1550), .A4(n1549), .ZN(n1553)
         );
  AOI22_X1 U1684 ( .A1(n70), .A2(n2665), .B1(n1553), .B2(n71), .ZN(N408) );
  AOI22_X1 U1685 ( .A1(\REGISTERS[16][30] ), .A2(n63), .B1(\REGISTERS[17][30] ), .B2(n52), .ZN(n1557) );
  AOI22_X1 U1686 ( .A1(\REGISTERS[30][30] ), .A2(n1615), .B1(
        \REGISTERS[4][30] ), .B2(n37), .ZN(n1556) );
  AOI22_X1 U1687 ( .A1(\REGISTERS[22][30] ), .A2(n51), .B1(\REGISTERS[27][30] ), .B2(n40), .ZN(n1555) );
  AOI22_X1 U1688 ( .A1(\REGISTERS[23][30] ), .A2(n1590), .B1(
        \REGISTERS[8][30] ), .B2(n38), .ZN(n1554) );
  NAND4_X1 U1689 ( .A1(n1557), .A2(n1556), .A3(n1555), .A4(n1554), .ZN(n1573)
         );
  AOI22_X1 U1690 ( .A1(\REGISTERS[3][30] ), .A2(n50), .B1(\REGISTERS[28][30] ), 
        .B2(n60), .ZN(n1561) );
  AOI22_X1 U1691 ( .A1(\REGISTERS[20][30] ), .A2(n66), .B1(\REGISTERS[14][30] ), .B2(n44), .ZN(n1560) );
  AOI22_X1 U1692 ( .A1(\REGISTERS[6][30] ), .A2(n67), .B1(\REGISTERS[11][30] ), 
        .B2(n49), .ZN(n1559) );
  AOI22_X1 U1693 ( .A1(\REGISTERS[13][30] ), .A2(n45), .B1(\REGISTERS[18][30] ), .B2(n59), .ZN(n1558) );
  NAND4_X1 U1694 ( .A1(n1561), .A2(n1560), .A3(n1559), .A4(n1558), .ZN(n1572)
         );
  AOI22_X1 U1695 ( .A1(\REGISTERS[15][30] ), .A2(n1601), .B1(
        \REGISTERS[21][30] ), .B2(n53), .ZN(n1565) );
  AOI22_X1 U1696 ( .A1(\REGISTERS[5][30] ), .A2(n1612), .B1(\REGISTERS[9][30] ), .B2(n42), .ZN(n1564) );
  AOI22_X1 U1697 ( .A1(\REGISTERS[31][30] ), .A2(n54), .B1(\REGISTERS[25][30] ), .B2(n61), .ZN(n1563) );
  AOI22_X1 U1698 ( .A1(\REGISTERS[12][30] ), .A2(n1602), .B1(
        \REGISTERS[0][30] ), .B2(n64), .ZN(n1562) );
  NAND4_X1 U1699 ( .A1(n1565), .A2(n1564), .A3(n1563), .A4(n1562), .ZN(n1571)
         );
  AOI22_X1 U1700 ( .A1(\REGISTERS[1][30] ), .A2(n1577), .B1(
        \REGISTERS[24][30] ), .B2(n47), .ZN(n1569) );
  AOI22_X1 U1701 ( .A1(\REGISTERS[26][30] ), .A2(n1603), .B1(
        \REGISTERS[2][30] ), .B2(n46), .ZN(n1568) );
  AOI22_X1 U1702 ( .A1(\REGISTERS[19][30] ), .A2(n1604), .B1(
        \REGISTERS[29][30] ), .B2(n68), .ZN(n1567) );
  AOI22_X1 U1703 ( .A1(\REGISTERS[10][30] ), .A2(n41), .B1(\REGISTERS[7][30] ), 
        .B2(n43), .ZN(n1566) );
  NAND4_X1 U1704 ( .A1(n1569), .A2(n1568), .A3(n1567), .A4(n1566), .ZN(n1570)
         );
  NOR4_X1 U1705 ( .A1(n1573), .A2(n1572), .A3(n1571), .A4(n1570), .ZN(n1574)
         );
  AOI22_X1 U1706 ( .A1(n70), .A2(n2664), .B1(n1574), .B2(n71), .ZN(N409) );
  AOI22_X1 U1707 ( .A1(\REGISTERS[8][31] ), .A2(n1576), .B1(\REGISTERS[4][31] ), .B2(n37), .ZN(n1586) );
  AOI22_X1 U1708 ( .A1(\REGISTERS[27][31] ), .A2(n1578), .B1(
        \REGISTERS[1][31] ), .B2(n39), .ZN(n1585) );
  AOI22_X1 U1709 ( .A1(\REGISTERS[9][31] ), .A2(n1580), .B1(
        \REGISTERS[10][31] ), .B2(n41), .ZN(n1584) );
  AOI22_X1 U1710 ( .A1(\REGISTERS[14][31] ), .A2(n1582), .B1(
        \REGISTERS[7][31] ), .B2(n43), .ZN(n1583) );
  NAND4_X1 U1711 ( .A1(n1586), .A2(n1585), .A3(n1584), .A4(n1583), .ZN(n1626)
         );
  AOI22_X1 U1712 ( .A1(\REGISTERS[2][31] ), .A2(n46), .B1(\REGISTERS[13][31] ), 
        .B2(n45), .ZN(n1598) );
  AOI22_X1 U1713 ( .A1(\REGISTERS[23][31] ), .A2(n1590), .B1(
        \REGISTERS[24][31] ), .B2(n47), .ZN(n1597) );
  AOI22_X1 U1714 ( .A1(\REGISTERS[3][31] ), .A2(n50), .B1(\REGISTERS[11][31] ), 
        .B2(n49), .ZN(n1596) );
  AOI22_X1 U1715 ( .A1(\REGISTERS[17][31] ), .A2(n52), .B1(\REGISTERS[22][31] ), .B2(n51), .ZN(n1595) );
  NAND4_X1 U1716 ( .A1(n1598), .A2(n1597), .A3(n1596), .A4(n1595), .ZN(n1625)
         );
  AOI22_X1 U1717 ( .A1(\REGISTERS[31][31] ), .A2(n1600), .B1(
        \REGISTERS[21][31] ), .B2(n53), .ZN(n1610) );
  AOI22_X1 U1718 ( .A1(\REGISTERS[12][31] ), .A2(n1602), .B1(
        \REGISTERS[15][31] ), .B2(n55), .ZN(n1609) );
  AOI22_X1 U1719 ( .A1(\REGISTERS[19][31] ), .A2(n58), .B1(\REGISTERS[26][31] ), .B2(n57), .ZN(n1608) );
  AOI22_X1 U1720 ( .A1(\REGISTERS[28][31] ), .A2(n1606), .B1(
        \REGISTERS[18][31] ), .B2(n59), .ZN(n1607) );
  NAND4_X1 U1721 ( .A1(n1610), .A2(n1609), .A3(n1608), .A4(n1607), .ZN(n1624)
         );
  AOI22_X1 U1722 ( .A1(\REGISTERS[5][31] ), .A2(n62), .B1(\REGISTERS[25][31] ), 
        .B2(n61), .ZN(n1622) );
  AOI22_X1 U1723 ( .A1(\REGISTERS[0][31] ), .A2(n1614), .B1(
        \REGISTERS[16][31] ), .B2(n63), .ZN(n1621) );
  AOI22_X1 U1724 ( .A1(\REGISTERS[20][31] ), .A2(n1616), .B1(
        \REGISTERS[30][31] ), .B2(n65), .ZN(n1620) );
  AOI22_X1 U1725 ( .A1(\REGISTERS[29][31] ), .A2(n1618), .B1(
        \REGISTERS[6][31] ), .B2(n67), .ZN(n1619) );
  NAND4_X1 U1726 ( .A1(n1622), .A2(n1621), .A3(n1620), .A4(n1619), .ZN(n1623)
         );
  NOR4_X1 U1727 ( .A1(n1626), .A2(n1625), .A3(n1624), .A4(n1623), .ZN(n1627)
         );
  AOI22_X1 U1728 ( .A1(n70), .A2(n2671), .B1(n1627), .B2(n71), .ZN(N410) );
  OAI21_X1 U1729 ( .B1(n1630), .B2(n1629), .A(RST), .ZN(N81) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_0 \clk_gate_REGISTERS_reg[0]  ( 
        .CLK(CLK), .EN(N144), .ENCLK(net2402), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_31 \clk_gate_REGISTERS_reg[1]  ( 
        .CLK(CLK), .EN(N143), .ENCLK(net2408), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_30 \clk_gate_REGISTERS_reg[2]  ( 
        .CLK(CLK), .EN(N142), .ENCLK(net2413), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_29 \clk_gate_REGISTERS_reg[3]  ( 
        .CLK(CLK), .EN(N141), .ENCLK(net2418), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_28 \clk_gate_REGISTERS_reg[4]  ( 
        .CLK(CLK), .EN(N140), .ENCLK(net2423), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_27 \clk_gate_REGISTERS_reg[5]  ( 
        .CLK(CLK), .EN(N139), .ENCLK(net2428), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_26 \clk_gate_REGISTERS_reg[6]  ( 
        .CLK(CLK), .EN(N138), .ENCLK(net2433), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_25 \clk_gate_REGISTERS_reg[7]  ( 
        .CLK(CLK), .EN(N137), .ENCLK(net2438), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_24 \clk_gate_REGISTERS_reg[8]  ( 
        .CLK(CLK), .EN(N136), .ENCLK(net2443), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_23 \clk_gate_REGISTERS_reg[9]  ( 
        .CLK(CLK), .EN(N135), .ENCLK(net2448), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_22 \clk_gate_REGISTERS_reg[10]  ( 
        .CLK(CLK), .EN(N134), .ENCLK(net2453), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_21 \clk_gate_REGISTERS_reg[11]  ( 
        .CLK(CLK), .EN(N133), .ENCLK(net2458), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_20 \clk_gate_REGISTERS_reg[12]  ( 
        .CLK(CLK), .EN(N132), .ENCLK(net2463), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_19 \clk_gate_REGISTERS_reg[13]  ( 
        .CLK(CLK), .EN(N131), .ENCLK(net2468), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_18 \clk_gate_REGISTERS_reg[14]  ( 
        .CLK(CLK), .EN(N130), .ENCLK(net2473), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_17 \clk_gate_REGISTERS_reg[15]  ( 
        .CLK(CLK), .EN(N129), .ENCLK(net2478), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_16 \clk_gate_REGISTERS_reg[16]  ( 
        .CLK(CLK), .EN(N128), .ENCLK(net2483), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_15 \clk_gate_REGISTERS_reg[17]  ( 
        .CLK(CLK), .EN(N127), .ENCLK(net2488), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_14 \clk_gate_REGISTERS_reg[18]  ( 
        .CLK(CLK), .EN(N126), .ENCLK(net2493), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_13 \clk_gate_REGISTERS_reg[19]  ( 
        .CLK(CLK), .EN(N125), .ENCLK(net2498), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_12 \clk_gate_REGISTERS_reg[20]  ( 
        .CLK(CLK), .EN(N124), .ENCLK(net2503), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_11 \clk_gate_REGISTERS_reg[21]  ( 
        .CLK(CLK), .EN(N123), .ENCLK(net2508), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_10 \clk_gate_REGISTERS_reg[22]  ( 
        .CLK(CLK), .EN(N122), .ENCLK(net2513), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_9 \clk_gate_REGISTERS_reg[23]  ( 
        .CLK(CLK), .EN(N121), .ENCLK(net2518), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_8 \clk_gate_REGISTERS_reg[24]  ( 
        .CLK(CLK), .EN(N120), .ENCLK(net2523), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_7 \clk_gate_REGISTERS_reg[25]  ( 
        .CLK(CLK), .EN(N119), .ENCLK(net2528), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_6 \clk_gate_REGISTERS_reg[26]  ( 
        .CLK(CLK), .EN(N118), .ENCLK(net2533), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_5 \clk_gate_REGISTERS_reg[27]  ( 
        .CLK(CLK), .EN(N117), .ENCLK(net2538), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_4 \clk_gate_REGISTERS_reg[28]  ( 
        .CLK(CLK), .EN(N116), .ENCLK(net2543), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_3 \clk_gate_REGISTERS_reg[29]  ( 
        .CLK(CLK), .EN(N115), .ENCLK(net2548), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_2 \clk_gate_REGISTERS_reg[30]  ( 
        .CLK(CLK), .EN(N114), .ENCLK(net2553), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_FILE_WIDTH32_LENGTH5_1 \clk_gate_REGISTERS_reg[31]  ( 
        .CLK(CLK), .EN(N81), .ENCLK(net2558), .TE(1'b0) );
  INV_X2 U34 ( .A(n100), .ZN(n99) );
  INV_X2 U50 ( .A(n122), .ZN(n121) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n2656), .CK(net2558), .Q(
        \REGISTERS[31][23] ) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n2655), .CK(net2548), .Q(
        \REGISTERS[29][23] ) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n2654), .CK(net2538), .Q(
        \REGISTERS[27][23] ) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n2653), .CK(net2528), .Q(
        \REGISTERS[25][23] ) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n2652), .CK(net2518), .Q(
        \REGISTERS[23][23] ) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n2651), .CK(net2508), .Q(
        \REGISTERS[21][23] ) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n2650), .CK(net2503), .Q(
        \REGISTERS[20][23] ) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n2649), .CK(net2493), .Q(
        \REGISTERS[18][23] ) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n2648), .CK(net2483), .Q(
        \REGISTERS[16][23] ) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n2647), .CK(net2473), .Q(
        \REGISTERS[14][23] ) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n2646), .CK(net2468), .Q(
        \REGISTERS[13][23] ) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n2645), .CK(net2463), .Q(
        \REGISTERS[12][23] ) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n2644), .CK(net2458), .Q(
        \REGISTERS[11][23] ) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n2643), .CK(net2453), .Q(
        \REGISTERS[10][23] ) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n2642), .CK(net2448), .Q(
        \REGISTERS[9][23] ) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n2641), .CK(net2443), .Q(
        \REGISTERS[8][23] ) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n2640), .CK(net2558), .Q(
        \REGISTERS[31][24] ) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n2639), .CK(net2548), .Q(
        \REGISTERS[29][24] ) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n2638), .CK(net2538), .Q(
        \REGISTERS[27][24] ) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n2637), .CK(net2528), .Q(
        \REGISTERS[25][24] ) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n2636), .CK(net2518), .Q(
        \REGISTERS[23][24] ) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n2635), .CK(net2508), .Q(
        \REGISTERS[21][24] ) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n2634), .CK(net2503), .Q(
        \REGISTERS[20][24] ) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n2633), .CK(net2493), .Q(
        \REGISTERS[18][24] ) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n2632), .CK(net2483), .Q(
        \REGISTERS[16][24] ) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n2631), .CK(net2473), .Q(
        \REGISTERS[14][24] ) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n2630), .CK(net2468), .Q(
        \REGISTERS[13][24] ) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n2629), .CK(net2463), .Q(
        \REGISTERS[12][24] ) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n2628), .CK(net2458), .Q(
        \REGISTERS[11][24] ) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n2627), .CK(net2453), .Q(
        \REGISTERS[10][24] ) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n2626), .CK(net2448), .Q(
        \REGISTERS[9][24] ) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n2625), .CK(net2443), .Q(
        \REGISTERS[8][24] ) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n2624), .CK(net2503), .Q(
        \REGISTERS[20][20] ) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n2623), .CK(net2493), .Q(
        \REGISTERS[18][20] ) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n2622), .CK(net2483), .Q(
        \REGISTERS[16][20] ) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n2621), .CK(net2473), .Q(
        \REGISTERS[14][20] ) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n2620), .CK(net2468), .Q(
        \REGISTERS[13][20] ) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n2619), .CK(net2463), .Q(
        \REGISTERS[12][20] ) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n2618), .CK(net2458), .Q(
        \REGISTERS[11][20] ) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n2617), .CK(net2453), .Q(
        \REGISTERS[10][20] ) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n2616), .CK(net2448), .Q(
        \REGISTERS[9][20] ) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n2615), .CK(net2443), .Q(
        \REGISTERS[8][20] ) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n2614), .CK(net2503), .Q(
        \REGISTERS[20][26] ) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n2613), .CK(net2493), .Q(
        \REGISTERS[18][26] ) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n2612), .CK(net2483), .Q(
        \REGISTERS[16][26] ) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n2611), .CK(net2473), .Q(
        \REGISTERS[14][26] ) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n2610), .CK(net2468), .Q(
        \REGISTERS[13][26] ) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n2609), .CK(net2463), .Q(
        \REGISTERS[12][26] ) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n2608), .CK(net2458), .Q(
        \REGISTERS[11][26] ) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n2607), .CK(net2453), .Q(
        \REGISTERS[10][26] ) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n2606), .CK(net2448), .Q(
        \REGISTERS[9][26] ) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n2605), .CK(net2443), .Q(
        \REGISTERS[8][26] ) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n2604), .CK(net2503), .Q(
        \REGISTERS[20][6] ) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n2603), .CK(net2493), .Q(
        \REGISTERS[18][6] ) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n2602), .CK(net2483), .Q(
        \REGISTERS[16][6] ) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n2601), .CK(net2473), .Q(
        \REGISTERS[14][6] ) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n2600), .CK(net2468), .Q(
        \REGISTERS[13][6] ) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n2599), .CK(net2463), .Q(
        \REGISTERS[12][6] ) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n2598), .CK(net2458), .Q(
        \REGISTERS[11][6] ) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n2597), .CK(net2453), .Q(
        \REGISTERS[10][6] ) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n2596), .CK(net2448), .Q(\REGISTERS[9][6] ) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n2595), .CK(net2443), .Q(\REGISTERS[8][6] ) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n2594), .CK(net2503), .Q(
        \REGISTERS[20][22] ) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n2593), .CK(net2503), .Q(
        \REGISTERS[20][3] ) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n2592), .CK(net2493), .Q(
        \REGISTERS[18][22] ) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n2591), .CK(net2493), .Q(
        \REGISTERS[18][3] ) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n2590), .CK(net2483), .Q(
        \REGISTERS[16][22] ) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n2589), .CK(net2483), .Q(
        \REGISTERS[16][3] ) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n2588), .CK(net2473), .Q(
        \REGISTERS[14][22] ) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n2587), .CK(net2473), .Q(
        \REGISTERS[14][3] ) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n2586), .CK(net2468), .Q(
        \REGISTERS[13][22] ) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n2585), .CK(net2468), .Q(
        \REGISTERS[13][3] ) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n2584), .CK(net2463), .Q(
        \REGISTERS[12][22] ) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n2583), .CK(net2463), .Q(
        \REGISTERS[12][3] ) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n2582), .CK(net2458), .Q(
        \REGISTERS[11][22] ) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n2581), .CK(net2458), .Q(
        \REGISTERS[11][3] ) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n2580), .CK(net2453), .Q(
        \REGISTERS[10][22] ) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n2579), .CK(net2453), .Q(
        \REGISTERS[10][3] ) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n2578), .CK(net2448), .Q(
        \REGISTERS[9][22] ) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n2577), .CK(net2448), .Q(\REGISTERS[9][3] ) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n2576), .CK(net2443), .Q(
        \REGISTERS[8][22] ) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n2575), .CK(net2443), .Q(\REGISTERS[8][3] ) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n2574), .CK(net2503), .Q(
        \REGISTERS[20][1] ) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n2573), .CK(net2493), .Q(
        \REGISTERS[18][1] ) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n2572), .CK(net2483), .Q(
        \REGISTERS[16][1] ) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n2571), .CK(net2473), .Q(
        \REGISTERS[14][1] ) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n2570), .CK(net2468), .Q(
        \REGISTERS[13][1] ) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n2569), .CK(net2463), .Q(
        \REGISTERS[12][1] ) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n2568), .CK(net2458), .Q(
        \REGISTERS[11][1] ) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n2567), .CK(net2453), .Q(
        \REGISTERS[10][1] ) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n2566), .CK(net2448), .Q(\REGISTERS[9][1] ) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n2565), .CK(net2443), .Q(\REGISTERS[8][1] ) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n2564), .CK(net2523), .Q(
        \REGISTERS[24][5] ) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n2563), .CK(net2503), .Q(
        \REGISTERS[20][5] ) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n2562), .CK(net2483), .Q(
        \REGISTERS[16][5] ) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n2561), .CK(net2473), .Q(
        \REGISTERS[14][5] ) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n2560), .CK(net2468), .Q(
        \REGISTERS[13][5] ) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n2559), .CK(net2463), .Q(
        \REGISTERS[12][5] ) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n2558), .CK(net2458), .Q(
        \REGISTERS[11][5] ) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n2557), .CK(net2453), .Q(
        \REGISTERS[10][5] ) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n2556), .CK(net2448), .Q(\REGISTERS[9][5] ) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n2555), .CK(net2443), .Q(\REGISTERS[8][5] ) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n2554), .CK(net2503), .Q(
        \REGISTERS[20][18] ) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n2553), .CK(net2493), .Q(
        \REGISTERS[18][18] ) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n2552), .CK(net2483), .Q(
        \REGISTERS[16][18] ) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n2551), .CK(net2473), .Q(
        \REGISTERS[14][18] ) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n2550), .CK(net2468), .Q(
        \REGISTERS[13][18] ) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n2549), .CK(net2463), .Q(
        \REGISTERS[12][18] ) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n2548), .CK(net2458), .Q(
        \REGISTERS[11][18] ) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n2547), .CK(net2453), .Q(
        \REGISTERS[10][18] ) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n2546), .CK(net2448), .Q(
        \REGISTERS[9][18] ) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n2545), .CK(net2443), .Q(
        \REGISTERS[8][18] ) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n2544), .CK(net2503), .Q(
        \REGISTERS[20][31] ) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n2543), .CK(net2503), .Q(
        \REGISTERS[20][8] ) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n2542), .CK(net2493), .Q(
        \REGISTERS[18][31] ) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n2541), .CK(net2493), .Q(
        \REGISTERS[18][8] ) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n2540), .CK(net2483), .Q(
        \REGISTERS[16][31] ) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n2539), .CK(net2483), .Q(
        \REGISTERS[16][8] ) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n2538), .CK(net2473), .Q(
        \REGISTERS[14][31] ) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n2537), .CK(net2473), .Q(
        \REGISTERS[14][8] ) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n2536), .CK(net2468), .Q(
        \REGISTERS[13][31] ) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n2535), .CK(net2468), .Q(
        \REGISTERS[13][8] ) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n2534), .CK(net2463), .Q(
        \REGISTERS[12][31] ) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n2533), .CK(net2463), .Q(
        \REGISTERS[12][8] ) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n2532), .CK(net2458), .Q(
        \REGISTERS[11][31] ) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n2531), .CK(net2458), .Q(
        \REGISTERS[11][8] ) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n2530), .CK(net2453), .Q(
        \REGISTERS[10][31] ) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n2529), .CK(net2453), .Q(
        \REGISTERS[10][8] ) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n2528), .CK(net2448), .Q(
        \REGISTERS[9][31] ) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n2527), .CK(net2448), .Q(\REGISTERS[9][8] ) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n2526), .CK(net2443), .Q(
        \REGISTERS[8][31] ) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n2525), .CK(net2443), .Q(\REGISTERS[8][8] ) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n2524), .CK(net2503), .Q(
        \REGISTERS[20][13] ) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n2523), .CK(net2493), .Q(
        \REGISTERS[18][13] ) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n2522), .CK(net2483), .Q(
        \REGISTERS[16][13] ) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n2521), .CK(net2473), .Q(
        \REGISTERS[14][13] ) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n2520), .CK(net2468), .Q(
        \REGISTERS[13][13] ) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n2519), .CK(net2463), .Q(
        \REGISTERS[12][13] ) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n2518), .CK(net2458), .Q(
        \REGISTERS[11][13] ) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n2517), .CK(net2453), .Q(
        \REGISTERS[10][13] ) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n2516), .CK(net2448), .Q(
        \REGISTERS[9][13] ) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n2515), .CK(net2443), .Q(
        \REGISTERS[8][13] ) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n2514), .CK(net2503), .Q(
        \REGISTERS[20][9] ) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n2513), .CK(net2493), .Q(
        \REGISTERS[18][9] ) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n2512), .CK(net2483), .Q(
        \REGISTERS[16][9] ) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n2511), .CK(net2473), .Q(
        \REGISTERS[14][9] ) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n2510), .CK(net2468), .Q(
        \REGISTERS[13][9] ) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n2509), .CK(net2463), .Q(
        \REGISTERS[12][9] ) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n2508), .CK(net2458), .Q(
        \REGISTERS[11][9] ) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n2507), .CK(net2453), .Q(
        \REGISTERS[10][9] ) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n2506), .CK(net2448), .Q(\REGISTERS[9][9] ) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n2505), .CK(net2443), .Q(\REGISTERS[8][9] ) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n2504), .CK(net2503), .Q(
        \REGISTERS[20][25] ) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n2503), .CK(net2493), .Q(
        \REGISTERS[18][25] ) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n2502), .CK(net2483), .Q(
        \REGISTERS[16][25] ) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n2501), .CK(net2473), .Q(
        \REGISTERS[14][25] ) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n2500), .CK(net2468), .Q(
        \REGISTERS[13][25] ) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n2499), .CK(net2463), .Q(
        \REGISTERS[12][25] ) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n2498), .CK(net2458), .Q(
        \REGISTERS[11][25] ) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n2497), .CK(net2453), .Q(
        \REGISTERS[10][25] ) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n2496), .CK(net2448), .Q(
        \REGISTERS[9][25] ) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n2495), .CK(net2443), .Q(
        \REGISTERS[8][25] ) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n2494), .CK(net2503), .Q(
        \REGISTERS[20][27] ) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n2493), .CK(net2493), .Q(
        \REGISTERS[18][27] ) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n2492), .CK(net2483), .Q(
        \REGISTERS[16][27] ) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n2491), .CK(net2473), .Q(
        \REGISTERS[14][27] ) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n2490), .CK(net2468), .Q(
        \REGISTERS[13][27] ) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n2489), .CK(net2463), .Q(
        \REGISTERS[12][27] ) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n2488), .CK(net2458), .Q(
        \REGISTERS[11][27] ) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n2487), .CK(net2453), .Q(
        \REGISTERS[10][27] ) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n2486), .CK(net2448), .Q(
        \REGISTERS[9][27] ) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n2485), .CK(net2443), .Q(
        \REGISTERS[8][27] ) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n2484), .CK(net2503), .Q(
        \REGISTERS[20][14] ) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n2483), .CK(net2493), .Q(
        \REGISTERS[18][14] ) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n2482), .CK(net2483), .Q(
        \REGISTERS[16][14] ) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n2481), .CK(net2473), .Q(
        \REGISTERS[14][14] ) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n2480), .CK(net2468), .Q(
        \REGISTERS[13][14] ) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n2479), .CK(net2463), .Q(
        \REGISTERS[12][14] ) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n2478), .CK(net2458), .Q(
        \REGISTERS[11][14] ) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n2477), .CK(net2453), .Q(
        \REGISTERS[10][14] ) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n2476), .CK(net2448), .Q(
        \REGISTERS[9][14] ) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n2475), .CK(net2443), .Q(
        \REGISTERS[8][14] ) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n2474), .CK(net2503), .Q(
        \REGISTERS[20][19] ) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n2473), .CK(net2493), .Q(
        \REGISTERS[18][19] ) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n2472), .CK(net2483), .Q(
        \REGISTERS[16][19] ) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n2471), .CK(net2473), .Q(
        \REGISTERS[14][19] ) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n2470), .CK(net2468), .Q(
        \REGISTERS[13][19] ) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n2469), .CK(net2463), .Q(
        \REGISTERS[12][19] ) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n2468), .CK(net2458), .Q(
        \REGISTERS[11][19] ) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n2467), .CK(net2453), .Q(
        \REGISTERS[10][19] ) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n2466), .CK(net2448), .Q(
        \REGISTERS[9][19] ) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n2465), .CK(net2443), .Q(
        \REGISTERS[8][19] ) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n2464), .CK(net2503), .Q(
        \REGISTERS[20][4] ) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n2463), .CK(net2493), .Q(
        \REGISTERS[18][4] ) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n2462), .CK(net2483), .Q(
        \REGISTERS[16][4] ) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n2461), .CK(net2473), .Q(
        \REGISTERS[14][4] ) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n2460), .CK(net2468), .Q(
        \REGISTERS[13][4] ) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n2459), .CK(net2463), .Q(
        \REGISTERS[12][4] ) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n2458), .CK(net2458), .Q(
        \REGISTERS[11][4] ) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n2457), .CK(net2453), .Q(
        \REGISTERS[10][4] ) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n2456), .CK(net2448), .Q(\REGISTERS[9][4] ) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n2455), .CK(net2443), .Q(\REGISTERS[8][4] ) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n2454), .CK(net2503), .Q(
        \REGISTERS[20][11] ) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n2453), .CK(net2493), .Q(
        \REGISTERS[18][11] ) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n2452), .CK(net2483), .Q(
        \REGISTERS[16][11] ) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n2451), .CK(net2473), .Q(
        \REGISTERS[14][11] ) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n2450), .CK(net2468), .Q(
        \REGISTERS[13][11] ) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n2449), .CK(net2463), .Q(
        \REGISTERS[12][11] ) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n2448), .CK(net2458), .Q(
        \REGISTERS[11][11] ) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n2447), .CK(net2453), .Q(
        \REGISTERS[10][11] ) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n2446), .CK(net2448), .Q(
        \REGISTERS[9][11] ) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n2445), .CK(net2443), .Q(
        \REGISTERS[8][11] ) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n2444), .CK(net2503), .Q(
        \REGISTERS[20][12] ) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n2443), .CK(net2493), .Q(
        \REGISTERS[18][12] ) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n2442), .CK(net2483), .Q(
        \REGISTERS[16][12] ) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n2441), .CK(net2473), .Q(
        \REGISTERS[14][12] ) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n2440), .CK(net2468), .Q(
        \REGISTERS[13][12] ) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n2439), .CK(net2463), .Q(
        \REGISTERS[12][12] ) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n2438), .CK(net2458), .Q(
        \REGISTERS[11][12] ) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n2437), .CK(net2453), .Q(
        \REGISTERS[10][12] ) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n2436), .CK(net2448), .Q(
        \REGISTERS[9][12] ) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n2435), .CK(net2443), .Q(
        \REGISTERS[8][12] ) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n2434), .CK(net2503), .Q(
        \REGISTERS[20][2] ) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n2433), .CK(net2493), .Q(
        \REGISTERS[18][2] ) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n2432), .CK(net2483), .Q(
        \REGISTERS[16][2] ) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n2431), .CK(net2473), .Q(
        \REGISTERS[14][2] ) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n2430), .CK(net2468), .Q(
        \REGISTERS[13][2] ) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n2429), .CK(net2463), .Q(
        \REGISTERS[12][2] ) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n2428), .CK(net2458), .Q(
        \REGISTERS[11][2] ) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n2427), .CK(net2453), .Q(
        \REGISTERS[10][2] ) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n2426), .CK(net2448), .Q(\REGISTERS[9][2] ) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n2425), .CK(net2443), .Q(\REGISTERS[8][2] ) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n2424), .CK(net2558), .Q(
        \REGISTERS[31][7] ) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n2423), .CK(net2548), .Q(
        \REGISTERS[29][7] ) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n2422), .CK(net2538), .Q(
        \REGISTERS[27][7] ) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n2421), .CK(net2528), .Q(
        \REGISTERS[25][7] ) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n2420), .CK(net2518), .Q(
        \REGISTERS[23][7] ) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n2419), .CK(net2508), .Q(
        \REGISTERS[21][7] ) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n2418), .CK(net2503), .Q(
        \REGISTERS[20][7] ) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n2417), .CK(net2493), .Q(
        \REGISTERS[18][7] ) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n2416), .CK(net2483), .Q(
        \REGISTERS[16][7] ) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n2415), .CK(net2473), .Q(
        \REGISTERS[14][7] ) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n2414), .CK(net2468), .Q(
        \REGISTERS[13][7] ) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n2413), .CK(net2463), .Q(
        \REGISTERS[12][7] ) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n2412), .CK(net2458), .Q(
        \REGISTERS[11][7] ) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n2411), .CK(net2453), .Q(
        \REGISTERS[10][7] ) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n2410), .CK(net2448), .Q(\REGISTERS[9][7] ) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n2409), .CK(net2443), .Q(\REGISTERS[8][7] ) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n2408), .CK(net2503), .Q(
        \REGISTERS[20][16] ) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n2407), .CK(net2493), .Q(
        \REGISTERS[18][16] ) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n2406), .CK(net2483), .Q(
        \REGISTERS[16][16] ) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n2405), .CK(net2473), .Q(
        \REGISTERS[14][16] ) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n2404), .CK(net2468), .Q(
        \REGISTERS[13][16] ) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n2403), .CK(net2463), .Q(
        \REGISTERS[12][16] ) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n2402), .CK(net2458), .Q(
        \REGISTERS[11][16] ) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n2401), .CK(net2453), .Q(
        \REGISTERS[10][16] ) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n2400), .CK(net2448), .Q(
        \REGISTERS[9][16] ) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n2399), .CK(net2443), .Q(
        \REGISTERS[8][16] ) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n2398), .CK(net2503), .Q(
        \REGISTERS[20][17] ) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n2397), .CK(net2493), .Q(
        \REGISTERS[18][17] ) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n2396), .CK(net2483), .Q(
        \REGISTERS[16][17] ) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n2395), .CK(net2473), .Q(
        \REGISTERS[14][17] ) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n2394), .CK(net2468), .Q(
        \REGISTERS[13][17] ) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n2393), .CK(net2463), .Q(
        \REGISTERS[12][17] ) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n2392), .CK(net2458), .Q(
        \REGISTERS[11][17] ) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n2391), .CK(net2453), .Q(
        \REGISTERS[10][17] ) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n2390), .CK(net2448), .Q(
        \REGISTERS[9][17] ) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n2389), .CK(net2443), .Q(
        \REGISTERS[8][17] ) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n2388), .CK(net2558), .Q(
        \REGISTERS[31][30] ) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n2387), .CK(net2553), .Q(
        \REGISTERS[30][30] ) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n2386), .CK(net2548), .Q(
        \REGISTERS[29][30] ) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n2385), .CK(net2543), .Q(
        \REGISTERS[28][30] ) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n2384), .CK(net2538), .Q(
        \REGISTERS[27][30] ) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n2383), .CK(net2533), .Q(
        \REGISTERS[26][30] ) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n2382), .CK(net2528), .Q(
        \REGISTERS[25][30] ) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n2381), .CK(net2523), .Q(
        \REGISTERS[24][30] ) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n2380), .CK(net2518), .Q(
        \REGISTERS[23][30] ) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n2379), .CK(net2513), .Q(
        \REGISTERS[22][30] ) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n2378), .CK(net2508), .Q(
        \REGISTERS[21][30] ) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n2377), .CK(net2503), .Q(
        \REGISTERS[20][30] ) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n2376), .CK(net2498), .Q(
        \REGISTERS[19][30] ) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n2375), .CK(net2493), .Q(
        \REGISTERS[18][30] ) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n2374), .CK(net2488), .Q(
        \REGISTERS[17][30] ) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n2373), .CK(net2483), .Q(
        \REGISTERS[16][30] ) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n2372), .CK(net2478), .Q(
        \REGISTERS[15][30] ) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n2371), .CK(net2473), .Q(
        \REGISTERS[14][30] ) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n2370), .CK(net2468), .Q(
        \REGISTERS[13][30] ) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n2369), .CK(net2463), .Q(
        \REGISTERS[12][30] ) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n2368), .CK(net2458), .Q(
        \REGISTERS[11][30] ) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n2367), .CK(net2453), .Q(
        \REGISTERS[10][30] ) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n2366), .CK(net2448), .Q(
        \REGISTERS[9][30] ) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n2365), .CK(net2443), .Q(
        \REGISTERS[8][30] ) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n2364), .CK(net2438), .Q(
        \REGISTERS[7][30] ) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n2363), .CK(net2433), .Q(
        \REGISTERS[6][30] ) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n2362), .CK(net2428), .Q(
        \REGISTERS[5][30] ) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n2361), .CK(net2423), .Q(
        \REGISTERS[4][30] ) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n2360), .CK(net2418), .Q(
        \REGISTERS[3][30] ) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n2359), .CK(net2413), .Q(
        \REGISTERS[2][30] ) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n2358), .CK(net2408), .Q(
        \REGISTERS[1][30] ) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n2357), .CK(net2402), .Q(
        \REGISTERS[0][30] ) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n2356), .CK(net2558), .Q(
        \REGISTERS[31][1] ) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n2355), .CK(net2553), .Q(
        \REGISTERS[30][1] ) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n2354), .CK(net2548), .Q(
        \REGISTERS[29][1] ) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n2353), .CK(net2543), .Q(
        \REGISTERS[28][1] ) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n2352), .CK(net2538), .Q(
        \REGISTERS[27][1] ) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n2351), .CK(net2533), .Q(
        \REGISTERS[26][1] ) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n2350), .CK(net2528), .Q(
        \REGISTERS[25][1] ) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n2349), .CK(net2523), .Q(
        \REGISTERS[24][1] ) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n2348), .CK(net2518), .Q(
        \REGISTERS[23][1] ) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n2347), .CK(net2513), .Q(
        \REGISTERS[22][1] ) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n2346), .CK(net2508), .Q(
        \REGISTERS[21][1] ) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n2345), .CK(net2498), .Q(
        \REGISTERS[19][1] ) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n2344), .CK(net2488), .Q(
        \REGISTERS[17][1] ) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n2343), .CK(net2478), .Q(
        \REGISTERS[15][1] ) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n2342), .CK(net2438), .Q(\REGISTERS[7][1] ) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n2341), .CK(net2433), .Q(\REGISTERS[6][1] ) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n2340), .CK(net2428), .Q(\REGISTERS[5][1] ) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n2339), .CK(net2423), .Q(\REGISTERS[4][1] ) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n2338), .CK(net2418), .Q(\REGISTERS[3][1] ) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n2337), .CK(net2413), .Q(\REGISTERS[2][1] ) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n2336), .CK(net2408), .Q(\REGISTERS[1][1] ) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n2335), .CK(net2402), .Q(\REGISTERS[0][1] ) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n2334), .CK(net2558), .Q(
        \REGISTERS[31][22] ) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n2333), .CK(net2558), .Q(
        \REGISTERS[31][3] ) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n2332), .CK(net2553), .Q(
        \REGISTERS[30][22] ) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n2331), .CK(net2553), .Q(
        \REGISTERS[30][3] ) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n2330), .CK(net2548), .Q(
        \REGISTERS[29][22] ) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n2329), .CK(net2548), .Q(
        \REGISTERS[29][3] ) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n2328), .CK(net2543), .Q(
        \REGISTERS[28][22] ) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n2327), .CK(net2543), .Q(
        \REGISTERS[28][3] ) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n2326), .CK(net2538), .Q(
        \REGISTERS[27][22] ) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n2325), .CK(net2538), .Q(
        \REGISTERS[27][3] ) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n2324), .CK(net2533), .Q(
        \REGISTERS[26][22] ) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n2323), .CK(net2533), .Q(
        \REGISTERS[26][3] ) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n2322), .CK(net2528), .Q(
        \REGISTERS[25][22] ) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n2321), .CK(net2528), .Q(
        \REGISTERS[25][3] ) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n2320), .CK(net2523), .Q(
        \REGISTERS[24][22] ) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n2319), .CK(net2523), .Q(
        \REGISTERS[24][3] ) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n2318), .CK(net2518), .Q(
        \REGISTERS[23][22] ) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n2317), .CK(net2518), .Q(
        \REGISTERS[23][3] ) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n2316), .CK(net2513), .Q(
        \REGISTERS[22][22] ) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n2315), .CK(net2513), .Q(
        \REGISTERS[22][3] ) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n2314), .CK(net2508), .Q(
        \REGISTERS[21][22] ) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n2313), .CK(net2508), .Q(
        \REGISTERS[21][3] ) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n2312), .CK(net2498), .Q(
        \REGISTERS[19][22] ) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n2311), .CK(net2498), .Q(
        \REGISTERS[19][3] ) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n2310), .CK(net2488), .Q(
        \REGISTERS[17][22] ) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n2309), .CK(net2488), .Q(
        \REGISTERS[17][3] ) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n2308), .CK(net2478), .Q(
        \REGISTERS[15][22] ) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n2307), .CK(net2478), .Q(
        \REGISTERS[15][3] ) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n2306), .CK(net2438), .Q(
        \REGISTERS[7][22] ) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n2305), .CK(net2438), .Q(\REGISTERS[7][3] ) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n2304), .CK(net2433), .Q(
        \REGISTERS[6][22] ) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n2303), .CK(net2433), .Q(\REGISTERS[6][3] ) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n2302), .CK(net2428), .Q(
        \REGISTERS[5][22] ) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n2301), .CK(net2428), .Q(\REGISTERS[5][3] ) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n2300), .CK(net2423), .Q(
        \REGISTERS[4][22] ) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n2299), .CK(net2423), .Q(\REGISTERS[4][3] ) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n2298), .CK(net2418), .Q(
        \REGISTERS[3][22] ) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n2297), .CK(net2418), .Q(\REGISTERS[3][3] ) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n2296), .CK(net2413), .Q(
        \REGISTERS[2][22] ) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n2295), .CK(net2413), .Q(\REGISTERS[2][3] ) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n2294), .CK(net2408), .Q(
        \REGISTERS[1][22] ) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n2293), .CK(net2408), .Q(\REGISTERS[1][3] ) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n2292), .CK(net2402), .Q(
        \REGISTERS[0][22] ) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n2291), .CK(net2402), .Q(\REGISTERS[0][3] ) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n2290), .CK(net2558), .Q(
        \REGISTERS[31][28] ) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n2289), .CK(net2553), .Q(
        \REGISTERS[30][28] ) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n2288), .CK(net2548), .Q(
        \REGISTERS[29][28] ) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n2287), .CK(net2543), .Q(
        \REGISTERS[28][28] ) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n2286), .CK(net2538), .Q(
        \REGISTERS[27][28] ) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n2285), .CK(net2533), .Q(
        \REGISTERS[26][28] ) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n2284), .CK(net2528), .Q(
        \REGISTERS[25][28] ) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n2283), .CK(net2523), .Q(
        \REGISTERS[24][28] ) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n2282), .CK(net2518), .Q(
        \REGISTERS[23][28] ) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n2281), .CK(net2513), .Q(
        \REGISTERS[22][28] ) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n2280), .CK(net2508), .Q(
        \REGISTERS[21][28] ) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n2279), .CK(net2503), .Q(
        \REGISTERS[20][28] ) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n2278), .CK(net2498), .Q(
        \REGISTERS[19][28] ) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n2277), .CK(net2493), .Q(
        \REGISTERS[18][28] ) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n2276), .CK(net2488), .Q(
        \REGISTERS[17][28] ) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n2275), .CK(net2483), .Q(
        \REGISTERS[16][28] ) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n2274), .CK(net2478), .Q(
        \REGISTERS[15][28] ) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n2273), .CK(net2473), .Q(
        \REGISTERS[14][28] ) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n2272), .CK(net2468), .Q(
        \REGISTERS[13][28] ) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n2271), .CK(net2463), .Q(
        \REGISTERS[12][28] ) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n2270), .CK(net2458), .Q(
        \REGISTERS[11][28] ) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n2269), .CK(net2453), .Q(
        \REGISTERS[10][28] ) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n2268), .CK(net2448), .Q(
        \REGISTERS[9][28] ) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n2267), .CK(net2443), .Q(
        \REGISTERS[8][28] ) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n2266), .CK(net2438), .Q(
        \REGISTERS[7][28] ) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n2265), .CK(net2433), .Q(
        \REGISTERS[6][28] ) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n2264), .CK(net2428), .Q(
        \REGISTERS[5][28] ) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n2263), .CK(net2423), .Q(
        \REGISTERS[4][28] ) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n2262), .CK(net2418), .Q(
        \REGISTERS[3][28] ) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n2261), .CK(net2413), .Q(
        \REGISTERS[2][28] ) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n2260), .CK(net2408), .Q(
        \REGISTERS[1][28] ) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n2259), .CK(net2402), .Q(
        \REGISTERS[0][28] ) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n2258), .CK(net2558), .Q(
        \REGISTERS[31][5] ) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n2257), .CK(net2553), .Q(
        \REGISTERS[30][5] ) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n2256), .CK(net2548), .Q(
        \REGISTERS[29][5] ) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n2255), .CK(net2543), .Q(
        \REGISTERS[28][5] ) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n2254), .CK(net2538), .Q(
        \REGISTERS[27][5] ) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n2253), .CK(net2533), .Q(
        \REGISTERS[26][5] ) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n2252), .CK(net2528), .Q(
        \REGISTERS[25][5] ) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n2251), .CK(net2518), .Q(
        \REGISTERS[23][5] ) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n2250), .CK(net2513), .Q(
        \REGISTERS[22][5] ) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n2249), .CK(net2508), .Q(
        \REGISTERS[21][5] ) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n2248), .CK(net2498), .Q(
        \REGISTERS[19][5] ) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n2247), .CK(net2493), .Q(
        \REGISTERS[18][5] ) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n2246), .CK(net2488), .Q(
        \REGISTERS[17][5] ) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n2245), .CK(net2478), .Q(
        \REGISTERS[15][5] ) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n2244), .CK(net2438), .Q(\REGISTERS[7][5] ) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n2243), .CK(net2433), .Q(\REGISTERS[6][5] ) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n2242), .CK(net2428), .Q(\REGISTERS[5][5] ) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n2241), .CK(net2423), .Q(\REGISTERS[4][5] ) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n2240), .CK(net2418), .Q(\REGISTERS[3][5] ) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n2239), .CK(net2413), .Q(\REGISTERS[2][5] ) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n2238), .CK(net2408), .Q(\REGISTERS[1][5] ) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n2237), .CK(net2402), .Q(\REGISTERS[0][5] ) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n2236), .CK(net2558), .Q(
        \REGISTERS[31][6] ) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n2235), .CK(net2553), .Q(
        \REGISTERS[30][6] ) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n2234), .CK(net2548), .Q(
        \REGISTERS[29][6] ) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n2233), .CK(net2543), .Q(
        \REGISTERS[28][6] ) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n2232), .CK(net2538), .Q(
        \REGISTERS[27][6] ) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n2231), .CK(net2533), .Q(
        \REGISTERS[26][6] ) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n2230), .CK(net2528), .Q(
        \REGISTERS[25][6] ) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n2229), .CK(net2523), .Q(
        \REGISTERS[24][6] ) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n2228), .CK(net2518), .Q(
        \REGISTERS[23][6] ) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n2227), .CK(net2513), .Q(
        \REGISTERS[22][6] ) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n2226), .CK(net2508), .Q(
        \REGISTERS[21][6] ) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n2225), .CK(net2498), .Q(
        \REGISTERS[19][6] ) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n2224), .CK(net2488), .Q(
        \REGISTERS[17][6] ) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n2223), .CK(net2478), .Q(
        \REGISTERS[15][6] ) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n2222), .CK(net2438), .Q(\REGISTERS[7][6] ) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n2221), .CK(net2433), .Q(\REGISTERS[6][6] ) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n2220), .CK(net2428), .Q(\REGISTERS[5][6] ) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n2219), .CK(net2423), .Q(\REGISTERS[4][6] ) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n2218), .CK(net2418), .Q(\REGISTERS[3][6] ) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n2217), .CK(net2413), .Q(\REGISTERS[2][6] ) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n2216), .CK(net2408), .Q(\REGISTERS[1][6] ) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n2215), .CK(net2402), .Q(\REGISTERS[0][6] ) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n2214), .CK(net2558), .Q(
        \REGISTERS[31][31] ) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n2213), .CK(net2558), .Q(
        \REGISTERS[31][8] ) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n2212), .CK(net2553), .Q(
        \REGISTERS[30][31] ) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n2211), .CK(net2553), .Q(
        \REGISTERS[30][8] ) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n2210), .CK(net2548), .Q(
        \REGISTERS[29][31] ) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n2209), .CK(net2548), .Q(
        \REGISTERS[29][8] ) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n2208), .CK(net2543), .Q(
        \REGISTERS[28][31] ) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n2207), .CK(net2543), .Q(
        \REGISTERS[28][8] ) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n2206), .CK(net2538), .Q(
        \REGISTERS[27][31] ) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n2205), .CK(net2538), .Q(
        \REGISTERS[27][8] ) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n2204), .CK(net2533), .Q(
        \REGISTERS[26][31] ) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n2203), .CK(net2533), .Q(
        \REGISTERS[26][8] ) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n2202), .CK(net2528), .Q(
        \REGISTERS[25][31] ) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n2201), .CK(net2528), .Q(
        \REGISTERS[25][8] ) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n2200), .CK(net2523), .Q(
        \REGISTERS[24][31] ) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n2199), .CK(net2523), .Q(
        \REGISTERS[24][8] ) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n2198), .CK(net2518), .Q(
        \REGISTERS[23][31] ) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n2197), .CK(net2518), .Q(
        \REGISTERS[23][8] ) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n2196), .CK(net2513), .Q(
        \REGISTERS[22][31] ) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n2195), .CK(net2513), .Q(
        \REGISTERS[22][8] ) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n2194), .CK(net2508), .Q(
        \REGISTERS[21][31] ) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n2193), .CK(net2508), .Q(
        \REGISTERS[21][8] ) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n2192), .CK(net2498), .Q(
        \REGISTERS[19][31] ) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n2191), .CK(net2498), .Q(
        \REGISTERS[19][8] ) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n2190), .CK(net2488), .Q(
        \REGISTERS[17][31] ) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n2189), .CK(net2488), .Q(
        \REGISTERS[17][8] ) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n2188), .CK(net2478), .Q(
        \REGISTERS[15][31] ) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n2187), .CK(net2478), .Q(
        \REGISTERS[15][8] ) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n2186), .CK(net2438), .Q(
        \REGISTERS[7][31] ) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n2185), .CK(net2438), .Q(\REGISTERS[7][8] ) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n2184), .CK(net2433), .Q(
        \REGISTERS[6][31] ) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n2183), .CK(net2433), .Q(\REGISTERS[6][8] ) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n2182), .CK(net2428), .Q(
        \REGISTERS[5][31] ) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n2181), .CK(net2428), .Q(\REGISTERS[5][8] ) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n2180), .CK(net2423), .Q(
        \REGISTERS[4][31] ) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n2179), .CK(net2423), .Q(\REGISTERS[4][8] ) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n2178), .CK(net2418), .Q(
        \REGISTERS[3][31] ) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n2177), .CK(net2418), .Q(\REGISTERS[3][8] ) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n2176), .CK(net2413), .Q(
        \REGISTERS[2][31] ) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n2175), .CK(net2413), .Q(\REGISTERS[2][8] ) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n2174), .CK(net2408), .Q(
        \REGISTERS[1][31] ) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n2173), .CK(net2408), .Q(\REGISTERS[1][8] ) );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n2172), .CK(net2402), .Q(
        \REGISTERS[0][31] ) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n2171), .CK(net2402), .Q(\REGISTERS[0][8] ) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n2170), .CK(net2558), .Q(
        \REGISTERS[31][26] ) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n2169), .CK(net2558), .Q(
        \REGISTERS[31][20] ) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n2168), .CK(net2553), .Q(
        \REGISTERS[30][26] ) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n2167), .CK(net2553), .Q(
        \REGISTERS[30][20] ) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n2166), .CK(net2548), .Q(
        \REGISTERS[29][26] ) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n2165), .CK(net2548), .Q(
        \REGISTERS[29][20] ) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n2164), .CK(net2543), .Q(
        \REGISTERS[28][26] ) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n2163), .CK(net2543), .Q(
        \REGISTERS[28][20] ) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n2162), .CK(net2538), .Q(
        \REGISTERS[27][26] ) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n2161), .CK(net2538), .Q(
        \REGISTERS[27][20] ) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n2160), .CK(net2533), .Q(
        \REGISTERS[26][26] ) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n2159), .CK(net2533), .Q(
        \REGISTERS[26][20] ) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n2158), .CK(net2528), .Q(
        \REGISTERS[25][26] ) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n2157), .CK(net2528), .Q(
        \REGISTERS[25][20] ) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n2156), .CK(net2523), .Q(
        \REGISTERS[24][26] ) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n2155), .CK(net2523), .Q(
        \REGISTERS[24][20] ) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n2154), .CK(net2518), .Q(
        \REGISTERS[23][26] ) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n2153), .CK(net2518), .Q(
        \REGISTERS[23][20] ) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n2152), .CK(net2513), .Q(
        \REGISTERS[22][26] ) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n2151), .CK(net2513), .Q(
        \REGISTERS[22][20] ) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n2150), .CK(net2508), .Q(
        \REGISTERS[21][26] ) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n2149), .CK(net2508), .Q(
        \REGISTERS[21][20] ) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n2148), .CK(net2498), .Q(
        \REGISTERS[19][26] ) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n2147), .CK(net2498), .Q(
        \REGISTERS[19][20] ) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n2146), .CK(net2488), .Q(
        \REGISTERS[17][26] ) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n2145), .CK(net2488), .Q(
        \REGISTERS[17][20] ) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n2144), .CK(net2478), .Q(
        \REGISTERS[15][26] ) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n2143), .CK(net2478), .Q(
        \REGISTERS[15][20] ) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n2142), .CK(net2438), .Q(
        \REGISTERS[7][26] ) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n2141), .CK(net2438), .Q(
        \REGISTERS[7][20] ) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n2140), .CK(net2433), .Q(
        \REGISTERS[6][26] ) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n2139), .CK(net2433), .Q(
        \REGISTERS[6][20] ) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n2138), .CK(net2428), .Q(
        \REGISTERS[5][26] ) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n2137), .CK(net2428), .Q(
        \REGISTERS[5][20] ) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n2136), .CK(net2423), .Q(
        \REGISTERS[4][26] ) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n2135), .CK(net2423), .Q(
        \REGISTERS[4][20] ) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n2134), .CK(net2418), .Q(
        \REGISTERS[3][26] ) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n2133), .CK(net2418), .Q(
        \REGISTERS[3][20] ) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n2132), .CK(net2413), .Q(
        \REGISTERS[2][26] ) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n2131), .CK(net2413), .Q(
        \REGISTERS[2][20] ) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n2130), .CK(net2408), .Q(
        \REGISTERS[1][26] ) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n2129), .CK(net2408), .Q(
        \REGISTERS[1][20] ) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n2128), .CK(net2402), .Q(
        \REGISTERS[0][26] ) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n2127), .CK(net2402), .Q(
        \REGISTERS[0][20] ) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n2126), .CK(net2558), .Q(
        \REGISTERS[31][9] ) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n2125), .CK(net2553), .Q(
        \REGISTERS[30][9] ) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n2124), .CK(net2548), .Q(
        \REGISTERS[29][9] ) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n2123), .CK(net2543), .Q(
        \REGISTERS[28][9] ) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n2122), .CK(net2538), .Q(
        \REGISTERS[27][9] ) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n2121), .CK(net2533), .Q(
        \REGISTERS[26][9] ) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n2120), .CK(net2528), .Q(
        \REGISTERS[25][9] ) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n2119), .CK(net2523), .Q(
        \REGISTERS[24][9] ) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n2118), .CK(net2518), .Q(
        \REGISTERS[23][9] ) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n2117), .CK(net2513), .Q(
        \REGISTERS[22][9] ) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n2116), .CK(net2508), .Q(
        \REGISTERS[21][9] ) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n2115), .CK(net2498), .Q(
        \REGISTERS[19][9] ) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n2114), .CK(net2488), .Q(
        \REGISTERS[17][9] ) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n2113), .CK(net2478), .Q(
        \REGISTERS[15][9] ) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n2112), .CK(net2438), .Q(\REGISTERS[7][9] ) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n2111), .CK(net2433), .Q(\REGISTERS[6][9] ) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n2110), .CK(net2428), .Q(\REGISTERS[5][9] ) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n2109), .CK(net2423), .Q(\REGISTERS[4][9] ) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n2108), .CK(net2418), .Q(\REGISTERS[3][9] ) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n2107), .CK(net2413), .Q(\REGISTERS[2][9] ) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n2106), .CK(net2408), .Q(\REGISTERS[1][9] ) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n2105), .CK(net2402), .Q(\REGISTERS[0][9] ) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n2104), .CK(net2558), .Q(
        \REGISTERS[31][10] ) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n2103), .CK(net2553), .Q(
        \REGISTERS[30][10] ) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n2102), .CK(net2548), .Q(
        \REGISTERS[29][10] ) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n2101), .CK(net2543), .Q(
        \REGISTERS[28][10] ) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n2100), .CK(net2538), .Q(
        \REGISTERS[27][10] ) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n2099), .CK(net2533), .Q(
        \REGISTERS[26][10] ) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n2098), .CK(net2528), .Q(
        \REGISTERS[25][10] ) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n2097), .CK(net2523), .Q(
        \REGISTERS[24][10] ) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n2096), .CK(net2518), .Q(
        \REGISTERS[23][10] ) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n2095), .CK(net2513), .Q(
        \REGISTERS[22][10] ) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n2094), .CK(net2508), .Q(
        \REGISTERS[21][10] ) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n2093), .CK(net2503), .Q(
        \REGISTERS[20][10] ) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n2092), .CK(net2498), .Q(
        \REGISTERS[19][10] ) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n2091), .CK(net2493), .Q(
        \REGISTERS[18][10] ) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n2090), .CK(net2488), .Q(
        \REGISTERS[17][10] ) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n2089), .CK(net2483), .Q(
        \REGISTERS[16][10] ) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n2088), .CK(net2478), .Q(
        \REGISTERS[15][10] ) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n2087), .CK(net2473), .Q(
        \REGISTERS[14][10] ) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n2086), .CK(net2468), .Q(
        \REGISTERS[13][10] ) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n2085), .CK(net2463), .Q(
        \REGISTERS[12][10] ) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n2084), .CK(net2458), .Q(
        \REGISTERS[11][10] ) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n2083), .CK(net2453), .Q(
        \REGISTERS[10][10] ) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n2082), .CK(net2448), .Q(
        \REGISTERS[9][10] ) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n2081), .CK(net2443), .Q(
        \REGISTERS[8][10] ) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n2080), .CK(net2438), .Q(
        \REGISTERS[7][10] ) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n2079), .CK(net2433), .Q(
        \REGISTERS[6][10] ) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n2078), .CK(net2428), .Q(
        \REGISTERS[5][10] ) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n2077), .CK(net2423), .Q(
        \REGISTERS[4][10] ) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n2076), .CK(net2418), .Q(
        \REGISTERS[3][10] ) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n2075), .CK(net2413), .Q(
        \REGISTERS[2][10] ) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n2074), .CK(net2408), .Q(
        \REGISTERS[1][10] ) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n2073), .CK(net2402), .Q(
        \REGISTERS[0][10] ) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n2072), .CK(net2558), .Q(
        \REGISTERS[31][15] ) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n2071), .CK(net2553), .Q(
        \REGISTERS[30][15] ) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n2070), .CK(net2548), .Q(
        \REGISTERS[29][15] ) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n2069), .CK(net2543), .Q(
        \REGISTERS[28][15] ) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n2068), .CK(net2538), .Q(
        \REGISTERS[27][15] ) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n2067), .CK(net2533), .Q(
        \REGISTERS[26][15] ) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n2066), .CK(net2528), .Q(
        \REGISTERS[25][15] ) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n2065), .CK(net2523), .Q(
        \REGISTERS[24][15] ) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n2064), .CK(net2518), .Q(
        \REGISTERS[23][15] ) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n2063), .CK(net2513), .Q(
        \REGISTERS[22][15] ) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n2062), .CK(net2508), .Q(
        \REGISTERS[21][15] ) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n2061), .CK(net2503), .Q(
        \REGISTERS[20][15] ) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n2060), .CK(net2498), .Q(
        \REGISTERS[19][15] ) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n2059), .CK(net2493), .Q(
        \REGISTERS[18][15] ) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n2058), .CK(net2488), .Q(
        \REGISTERS[17][15] ) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n2057), .CK(net2483), .Q(
        \REGISTERS[16][15] ) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n2056), .CK(net2478), .Q(
        \REGISTERS[15][15] ) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n2055), .CK(net2473), .Q(
        \REGISTERS[14][15] ) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n2054), .CK(net2468), .Q(
        \REGISTERS[13][15] ) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n2053), .CK(net2463), .Q(
        \REGISTERS[12][15] ) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n2052), .CK(net2458), .Q(
        \REGISTERS[11][15] ) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n2051), .CK(net2453), .Q(
        \REGISTERS[10][15] ) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n2050), .CK(net2448), .Q(
        \REGISTERS[9][15] ) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n2049), .CK(net2443), .Q(
        \REGISTERS[8][15] ) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n2048), .CK(net2438), .Q(
        \REGISTERS[7][15] ) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n2047), .CK(net2433), .Q(
        \REGISTERS[6][15] ) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n2046), .CK(net2428), .Q(
        \REGISTERS[5][15] ) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n2045), .CK(net2423), .Q(
        \REGISTERS[4][15] ) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n2044), .CK(net2418), .Q(
        \REGISTERS[3][15] ) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n2043), .CK(net2413), .Q(
        \REGISTERS[2][15] ) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n2042), .CK(net2408), .Q(
        \REGISTERS[1][15] ) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n2041), .CK(net2402), .Q(
        \REGISTERS[0][15] ) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n2040), .CK(net2558), .Q(
        \REGISTERS[31][29] ) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n2039), .CK(net2553), .Q(
        \REGISTERS[30][29] ) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n2038), .CK(net2548), .Q(
        \REGISTERS[29][29] ) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n2037), .CK(net2543), .Q(
        \REGISTERS[28][29] ) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n2036), .CK(net2538), .Q(
        \REGISTERS[27][29] ) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n2035), .CK(net2533), .Q(
        \REGISTERS[26][29] ) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n2034), .CK(net2528), .Q(
        \REGISTERS[25][29] ) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n2033), .CK(net2523), .Q(
        \REGISTERS[24][29] ) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n2032), .CK(net2518), .Q(
        \REGISTERS[23][29] ) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n2031), .CK(net2513), .Q(
        \REGISTERS[22][29] ) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n2030), .CK(net2508), .Q(
        \REGISTERS[21][29] ) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n2029), .CK(net2503), .Q(
        \REGISTERS[20][29] ) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n2028), .CK(net2498), .Q(
        \REGISTERS[19][29] ) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n2027), .CK(net2493), .Q(
        \REGISTERS[18][29] ) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n2026), .CK(net2488), .Q(
        \REGISTERS[17][29] ) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n2025), .CK(net2483), .Q(
        \REGISTERS[16][29] ) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n2024), .CK(net2478), .Q(
        \REGISTERS[15][29] ) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n2023), .CK(net2473), .Q(
        \REGISTERS[14][29] ) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n2022), .CK(net2468), .Q(
        \REGISTERS[13][29] ) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n2021), .CK(net2463), .Q(
        \REGISTERS[12][29] ) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n2020), .CK(net2458), .Q(
        \REGISTERS[11][29] ) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n2019), .CK(net2453), .Q(
        \REGISTERS[10][29] ) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n2018), .CK(net2448), .Q(
        \REGISTERS[9][29] ) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n2017), .CK(net2443), .Q(
        \REGISTERS[8][29] ) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n2016), .CK(net2438), .Q(
        \REGISTERS[7][29] ) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n2015), .CK(net2433), .Q(
        \REGISTERS[6][29] ) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n2014), .CK(net2428), .Q(
        \REGISTERS[5][29] ) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n2013), .CK(net2423), .Q(
        \REGISTERS[4][29] ) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n2012), .CK(net2418), .Q(
        \REGISTERS[3][29] ) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n2011), .CK(net2413), .Q(
        \REGISTERS[2][29] ) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n2010), .CK(net2408), .Q(
        \REGISTERS[1][29] ) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n2009), .CK(net2402), .Q(
        \REGISTERS[0][29] ) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n2008), .CK(net2553), .Q(
        \REGISTERS[30][23] ) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n2007), .CK(net2543), .Q(
        \REGISTERS[28][23] ) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n2006), .CK(net2533), .Q(
        \REGISTERS[26][23] ) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n2005), .CK(net2523), .Q(
        \REGISTERS[24][23] ) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n2004), .CK(net2513), .Q(
        \REGISTERS[22][23] ) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n2003), .CK(net2498), .Q(
        \REGISTERS[19][23] ) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n2002), .CK(net2488), .Q(
        \REGISTERS[17][23] ) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n2001), .CK(net2478), .Q(
        \REGISTERS[15][23] ) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n2000), .CK(net2438), .Q(
        \REGISTERS[7][23] ) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n1999), .CK(net2433), .Q(
        \REGISTERS[6][23] ) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n1998), .CK(net2428), .Q(
        \REGISTERS[5][23] ) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n1997), .CK(net2423), .Q(
        \REGISTERS[4][23] ) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n1996), .CK(net2418), .Q(
        \REGISTERS[3][23] ) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n1995), .CK(net2413), .Q(
        \REGISTERS[2][23] ) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n1994), .CK(net2408), .Q(
        \REGISTERS[1][23] ) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n1993), .CK(net2402), .Q(
        \REGISTERS[0][23] ) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n1992), .CK(net2553), .Q(
        \REGISTERS[30][24] ) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n1991), .CK(net2543), .Q(
        \REGISTERS[28][24] ) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n1990), .CK(net2533), .Q(
        \REGISTERS[26][24] ) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n1989), .CK(net2523), .Q(
        \REGISTERS[24][24] ) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n1988), .CK(net2513), .Q(
        \REGISTERS[22][24] ) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n1987), .CK(net2498), .Q(
        \REGISTERS[19][24] ) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n1986), .CK(net2488), .Q(
        \REGISTERS[17][24] ) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n1985), .CK(net2478), .Q(
        \REGISTERS[15][24] ) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n1984), .CK(net2438), .Q(
        \REGISTERS[7][24] ) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n1983), .CK(net2433), .Q(
        \REGISTERS[6][24] ) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n1982), .CK(net2428), .Q(
        \REGISTERS[5][24] ) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n1981), .CK(net2423), .Q(
        \REGISTERS[4][24] ) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n1980), .CK(net2418), .Q(
        \REGISTERS[3][24] ) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n1979), .CK(net2413), .Q(
        \REGISTERS[2][24] ) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n1978), .CK(net2408), .Q(
        \REGISTERS[1][24] ) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n1977), .CK(net2402), .Q(
        \REGISTERS[0][24] ) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n1976), .CK(net2558), .Q(
        \REGISTERS[31][0] ) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n1975), .CK(net2553), .Q(
        \REGISTERS[30][0] ) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n1974), .CK(net2548), .Q(
        \REGISTERS[29][0] ) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n1973), .CK(net2543), .Q(
        \REGISTERS[28][0] ) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n1972), .CK(net2538), .Q(
        \REGISTERS[27][0] ) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n1971), .CK(net2533), .Q(
        \REGISTERS[26][0] ) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n1970), .CK(net2528), .Q(
        \REGISTERS[25][0] ) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n1969), .CK(net2523), .Q(
        \REGISTERS[24][0] ) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n1968), .CK(net2518), .Q(
        \REGISTERS[23][0] ) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n1967), .CK(net2513), .Q(
        \REGISTERS[22][0] ) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n1966), .CK(net2508), .Q(
        \REGISTERS[21][0] ) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n1965), .CK(net2503), .Q(
        \REGISTERS[20][0] ) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n1964), .CK(net2498), .Q(
        \REGISTERS[19][0] ) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n1963), .CK(net2493), .Q(
        \REGISTERS[18][0] ) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n1962), .CK(net2488), .Q(
        \REGISTERS[17][0] ) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n1961), .CK(net2483), .Q(
        \REGISTERS[16][0] ) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n1960), .CK(net2478), .Q(
        \REGISTERS[15][0] ) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n1959), .CK(net2473), .Q(
        \REGISTERS[14][0] ) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n1958), .CK(net2468), .Q(
        \REGISTERS[13][0] ) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n1957), .CK(net2463), .Q(
        \REGISTERS[12][0] ) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n1956), .CK(net2458), .Q(
        \REGISTERS[11][0] ) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n1955), .CK(net2453), .Q(
        \REGISTERS[10][0] ) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n1954), .CK(net2448), .Q(\REGISTERS[9][0] ) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n1953), .CK(net2443), .Q(\REGISTERS[8][0] ) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n1952), .CK(net2438), .Q(\REGISTERS[7][0] ) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n1951), .CK(net2433), .Q(\REGISTERS[6][0] ) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n1950), .CK(net2428), .Q(\REGISTERS[5][0] ) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n1949), .CK(net2423), .Q(\REGISTERS[4][0] ) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n1948), .CK(net2418), .Q(\REGISTERS[3][0] ) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n1947), .CK(net2413), .Q(\REGISTERS[2][0] ) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n1946), .CK(net2408), .Q(\REGISTERS[1][0] ) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n1945), .CK(net2402), .Q(\REGISTERS[0][0] ) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n1944), .CK(net2558), .Q(
        \REGISTERS[31][27] ) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n1943), .CK(net2553), .Q(
        \REGISTERS[30][27] ) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n1942), .CK(net2548), .Q(
        \REGISTERS[29][27] ) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n1941), .CK(net2543), .Q(
        \REGISTERS[28][27] ) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n1940), .CK(net2538), .Q(
        \REGISTERS[27][27] ) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n1939), .CK(net2533), .Q(
        \REGISTERS[26][27] ) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n1938), .CK(net2528), .Q(
        \REGISTERS[25][27] ) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n1937), .CK(net2523), .Q(
        \REGISTERS[24][27] ) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n1936), .CK(net2518), .Q(
        \REGISTERS[23][27] ) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n1935), .CK(net2513), .Q(
        \REGISTERS[22][27] ) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n1934), .CK(net2508), .Q(
        \REGISTERS[21][27] ) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n1933), .CK(net2498), .Q(
        \REGISTERS[19][27] ) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n1932), .CK(net2488), .Q(
        \REGISTERS[17][27] ) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n1931), .CK(net2478), .Q(
        \REGISTERS[15][27] ) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n1930), .CK(net2438), .Q(
        \REGISTERS[7][27] ) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n1929), .CK(net2433), .Q(
        \REGISTERS[6][27] ) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n1928), .CK(net2428), .Q(
        \REGISTERS[5][27] ) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n1927), .CK(net2423), .Q(
        \REGISTERS[4][27] ) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n1926), .CK(net2418), .Q(
        \REGISTERS[3][27] ) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n1925), .CK(net2413), .Q(
        \REGISTERS[2][27] ) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n1924), .CK(net2408), .Q(
        \REGISTERS[1][27] ) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n1923), .CK(net2402), .Q(
        \REGISTERS[0][27] ) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n1922), .CK(net2558), .Q(
        \REGISTERS[31][18] ) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n1921), .CK(net2553), .Q(
        \REGISTERS[30][18] ) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n1920), .CK(net2548), .Q(
        \REGISTERS[29][18] ) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n1919), .CK(net2543), .Q(
        \REGISTERS[28][18] ) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n1918), .CK(net2538), .Q(
        \REGISTERS[27][18] ) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n1917), .CK(net2533), .Q(
        \REGISTERS[26][18] ) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n1916), .CK(net2528), .Q(
        \REGISTERS[25][18] ) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n1915), .CK(net2523), .Q(
        \REGISTERS[24][18] ) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n1914), .CK(net2518), .Q(
        \REGISTERS[23][18] ) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n1913), .CK(net2513), .Q(
        \REGISTERS[22][18] ) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n1912), .CK(net2508), .Q(
        \REGISTERS[21][18] ) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n1911), .CK(net2498), .Q(
        \REGISTERS[19][18] ) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n1910), .CK(net2488), .Q(
        \REGISTERS[17][18] ) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n1909), .CK(net2478), .Q(
        \REGISTERS[15][18] ) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n1908), .CK(net2438), .Q(
        \REGISTERS[7][18] ) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n1907), .CK(net2433), .Q(
        \REGISTERS[6][18] ) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n1906), .CK(net2428), .Q(
        \REGISTERS[5][18] ) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n1905), .CK(net2423), .Q(
        \REGISTERS[4][18] ) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n1904), .CK(net2418), .Q(
        \REGISTERS[3][18] ) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n1903), .CK(net2413), .Q(
        \REGISTERS[2][18] ) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n1902), .CK(net2408), .Q(
        \REGISTERS[1][18] ) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n1901), .CK(net2402), .Q(
        \REGISTERS[0][18] ) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n1900), .CK(net2558), .Q(
        \REGISTERS[31][14] ) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n1899), .CK(net2553), .Q(
        \REGISTERS[30][14] ) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n1898), .CK(net2548), .Q(
        \REGISTERS[29][14] ) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n1897), .CK(net2543), .Q(
        \REGISTERS[28][14] ) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n1896), .CK(net2538), .Q(
        \REGISTERS[27][14] ) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n1895), .CK(net2533), .Q(
        \REGISTERS[26][14] ) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n1894), .CK(net2528), .Q(
        \REGISTERS[25][14] ) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n1893), .CK(net2523), .Q(
        \REGISTERS[24][14] ) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n1892), .CK(net2518), .Q(
        \REGISTERS[23][14] ) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n1891), .CK(net2513), .Q(
        \REGISTERS[22][14] ) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n1890), .CK(net2508), .Q(
        \REGISTERS[21][14] ) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n1889), .CK(net2498), .Q(
        \REGISTERS[19][14] ) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n1888), .CK(net2488), .Q(
        \REGISTERS[17][14] ) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n1887), .CK(net2478), .Q(
        \REGISTERS[15][14] ) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n1886), .CK(net2438), .Q(
        \REGISTERS[7][14] ) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n1885), .CK(net2433), .Q(
        \REGISTERS[6][14] ) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n1884), .CK(net2428), .Q(
        \REGISTERS[5][14] ) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n1883), .CK(net2423), .Q(
        \REGISTERS[4][14] ) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n1882), .CK(net2418), .Q(
        \REGISTERS[3][14] ) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n1881), .CK(net2413), .Q(
        \REGISTERS[2][14] ) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n1880), .CK(net2408), .Q(
        \REGISTERS[1][14] ) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n1879), .CK(net2402), .Q(
        \REGISTERS[0][14] ) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n1878), .CK(net2558), .Q(
        \REGISTERS[31][13] ) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n1877), .CK(net2553), .Q(
        \REGISTERS[30][13] ) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n1876), .CK(net2548), .Q(
        \REGISTERS[29][13] ) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n1875), .CK(net2543), .Q(
        \REGISTERS[28][13] ) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n1874), .CK(net2538), .Q(
        \REGISTERS[27][13] ) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n1873), .CK(net2533), .Q(
        \REGISTERS[26][13] ) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n1872), .CK(net2528), .Q(
        \REGISTERS[25][13] ) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n1871), .CK(net2523), .Q(
        \REGISTERS[24][13] ) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n1870), .CK(net2518), .Q(
        \REGISTERS[23][13] ) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n1869), .CK(net2513), .Q(
        \REGISTERS[22][13] ) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n1868), .CK(net2508), .Q(
        \REGISTERS[21][13] ) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n1867), .CK(net2498), .Q(
        \REGISTERS[19][13] ) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n1866), .CK(net2488), .Q(
        \REGISTERS[17][13] ) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n1865), .CK(net2478), .Q(
        \REGISTERS[15][13] ) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n1864), .CK(net2438), .Q(
        \REGISTERS[7][13] ) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n1863), .CK(net2433), .Q(
        \REGISTERS[6][13] ) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n1862), .CK(net2428), .Q(
        \REGISTERS[5][13] ) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n1861), .CK(net2423), .Q(
        \REGISTERS[4][13] ) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n1860), .CK(net2418), .Q(
        \REGISTERS[3][13] ) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n1859), .CK(net2413), .Q(
        \REGISTERS[2][13] ) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n1858), .CK(net2408), .Q(
        \REGISTERS[1][13] ) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n1857), .CK(net2402), .Q(
        \REGISTERS[0][13] ) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n1856), .CK(net2558), .Q(
        \REGISTERS[31][25] ) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n1855), .CK(net2553), .Q(
        \REGISTERS[30][25] ) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n1854), .CK(net2548), .Q(
        \REGISTERS[29][25] ) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n1853), .CK(net2543), .Q(
        \REGISTERS[28][25] ) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n1852), .CK(net2538), .Q(
        \REGISTERS[27][25] ) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n1851), .CK(net2533), .Q(
        \REGISTERS[26][25] ) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n1850), .CK(net2528), .Q(
        \REGISTERS[25][25] ) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n1849), .CK(net2523), .Q(
        \REGISTERS[24][25] ) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n1848), .CK(net2518), .Q(
        \REGISTERS[23][25] ) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n1847), .CK(net2513), .Q(
        \REGISTERS[22][25] ) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n1846), .CK(net2508), .Q(
        \REGISTERS[21][25] ) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n1845), .CK(net2498), .Q(
        \REGISTERS[19][25] ) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n1844), .CK(net2488), .Q(
        \REGISTERS[17][25] ) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n1843), .CK(net2478), .Q(
        \REGISTERS[15][25] ) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n1842), .CK(net2438), .Q(
        \REGISTERS[7][25] ) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n1841), .CK(net2433), .Q(
        \REGISTERS[6][25] ) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n1840), .CK(net2428), .Q(
        \REGISTERS[5][25] ) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n1839), .CK(net2423), .Q(
        \REGISTERS[4][25] ) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n1838), .CK(net2418), .Q(
        \REGISTERS[3][25] ) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n1837), .CK(net2413), .Q(
        \REGISTERS[2][25] ) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n1836), .CK(net2408), .Q(
        \REGISTERS[1][25] ) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n1835), .CK(net2402), .Q(
        \REGISTERS[0][25] ) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n1834), .CK(net2558), .Q(
        \REGISTERS[31][21] ) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n1833), .CK(net2553), .Q(
        \REGISTERS[30][21] ) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n1832), .CK(net2548), .Q(
        \REGISTERS[29][21] ) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n1831), .CK(net2543), .Q(
        \REGISTERS[28][21] ) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n1830), .CK(net2538), .Q(
        \REGISTERS[27][21] ) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n1829), .CK(net2533), .Q(
        \REGISTERS[26][21] ) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n1828), .CK(net2528), .Q(
        \REGISTERS[25][21] ) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n1827), .CK(net2523), .Q(
        \REGISTERS[24][21] ) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n1826), .CK(net2518), .Q(
        \REGISTERS[23][21] ) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n1825), .CK(net2513), .Q(
        \REGISTERS[22][21] ) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n1824), .CK(net2508), .Q(
        \REGISTERS[21][21] ) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n1823), .CK(net2503), .Q(
        \REGISTERS[20][21] ) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n1822), .CK(net2498), .Q(
        \REGISTERS[19][21] ) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n1821), .CK(net2493), .Q(
        \REGISTERS[18][21] ) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n1820), .CK(net2488), .Q(
        \REGISTERS[17][21] ) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n1819), .CK(net2483), .Q(
        \REGISTERS[16][21] ) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n1818), .CK(net2478), .Q(
        \REGISTERS[15][21] ) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n1817), .CK(net2473), .Q(
        \REGISTERS[14][21] ) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n1816), .CK(net2468), .Q(
        \REGISTERS[13][21] ) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n1815), .CK(net2463), .Q(
        \REGISTERS[12][21] ) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n1814), .CK(net2458), .Q(
        \REGISTERS[11][21] ) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n1813), .CK(net2453), .Q(
        \REGISTERS[10][21] ) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n1812), .CK(net2448), .Q(
        \REGISTERS[9][21] ) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n1811), .CK(net2443), .Q(
        \REGISTERS[8][21] ) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n1810), .CK(net2438), .Q(
        \REGISTERS[7][21] ) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n1809), .CK(net2433), .Q(
        \REGISTERS[6][21] ) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n1808), .CK(net2428), .Q(
        \REGISTERS[5][21] ) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n1807), .CK(net2423), .Q(
        \REGISTERS[4][21] ) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n1806), .CK(net2418), .Q(
        \REGISTERS[3][21] ) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n1805), .CK(net2413), .Q(
        \REGISTERS[2][21] ) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n1804), .CK(net2408), .Q(
        \REGISTERS[1][21] ) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n1803), .CK(net2402), .Q(
        \REGISTERS[0][21] ) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n1802), .CK(net2553), .Q(
        \REGISTERS[30][7] ) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n1801), .CK(net2543), .Q(
        \REGISTERS[28][7] ) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n1800), .CK(net2533), .Q(
        \REGISTERS[26][7] ) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n1799), .CK(net2523), .Q(
        \REGISTERS[24][7] ) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n1798), .CK(net2513), .Q(
        \REGISTERS[22][7] ) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n1797), .CK(net2498), .Q(
        \REGISTERS[19][7] ) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n1796), .CK(net2488), .Q(
        \REGISTERS[17][7] ) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n1795), .CK(net2478), .Q(
        \REGISTERS[15][7] ) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n1794), .CK(net2438), .Q(\REGISTERS[7][7] ) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n1793), .CK(net2433), .Q(\REGISTERS[6][7] ) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n1792), .CK(net2428), .Q(\REGISTERS[5][7] ) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n1791), .CK(net2423), .Q(\REGISTERS[4][7] ) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n1790), .CK(net2418), .Q(\REGISTERS[3][7] ) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n1789), .CK(net2413), .Q(\REGISTERS[2][7] ) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n1788), .CK(net2408), .Q(\REGISTERS[1][7] ) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n1787), .CK(net2402), .Q(\REGISTERS[0][7] ) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n1786), .CK(net2558), .Q(
        \REGISTERS[31][4] ) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n1785), .CK(net2553), .Q(
        \REGISTERS[30][4] ) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n1784), .CK(net2548), .Q(
        \REGISTERS[29][4] ) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n1783), .CK(net2543), .Q(
        \REGISTERS[28][4] ) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n1782), .CK(net2538), .Q(
        \REGISTERS[27][4] ) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n1781), .CK(net2533), .Q(
        \REGISTERS[26][4] ) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n1780), .CK(net2528), .Q(
        \REGISTERS[25][4] ) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n1779), .CK(net2523), .Q(
        \REGISTERS[24][4] ) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n1778), .CK(net2518), .Q(
        \REGISTERS[23][4] ) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n1777), .CK(net2513), .Q(
        \REGISTERS[22][4] ) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n1776), .CK(net2508), .Q(
        \REGISTERS[21][4] ) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n1775), .CK(net2498), .Q(
        \REGISTERS[19][4] ) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n1774), .CK(net2488), .Q(
        \REGISTERS[17][4] ) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n1773), .CK(net2478), .Q(
        \REGISTERS[15][4] ) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n1772), .CK(net2438), .Q(\REGISTERS[7][4] ) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n1771), .CK(net2433), .Q(\REGISTERS[6][4] ) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n1770), .CK(net2428), .Q(\REGISTERS[5][4] ) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n1769), .CK(net2423), .Q(\REGISTERS[4][4] ) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n1768), .CK(net2418), .Q(\REGISTERS[3][4] ) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n1767), .CK(net2413), .Q(\REGISTERS[2][4] ) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n1766), .CK(net2408), .Q(\REGISTERS[1][4] ) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n1765), .CK(net2402), .Q(\REGISTERS[0][4] ) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n1764), .CK(net2558), .Q(
        \REGISTERS[31][19] ) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n1763), .CK(net2553), .Q(
        \REGISTERS[30][19] ) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n1762), .CK(net2548), .Q(
        \REGISTERS[29][19] ) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n1761), .CK(net2543), .Q(
        \REGISTERS[28][19] ) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n1760), .CK(net2538), .Q(
        \REGISTERS[27][19] ) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n1759), .CK(net2533), .Q(
        \REGISTERS[26][19] ) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n1758), .CK(net2528), .Q(
        \REGISTERS[25][19] ) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n1757), .CK(net2523), .Q(
        \REGISTERS[24][19] ) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n1756), .CK(net2518), .Q(
        \REGISTERS[23][19] ) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n1755), .CK(net2513), .Q(
        \REGISTERS[22][19] ) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n1754), .CK(net2508), .Q(
        \REGISTERS[21][19] ) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n1753), .CK(net2498), .Q(
        \REGISTERS[19][19] ) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n1752), .CK(net2488), .Q(
        \REGISTERS[17][19] ) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n1751), .CK(net2478), .Q(
        \REGISTERS[15][19] ) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n1750), .CK(net2438), .Q(
        \REGISTERS[7][19] ) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n1749), .CK(net2433), .Q(
        \REGISTERS[6][19] ) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n1748), .CK(net2428), .Q(
        \REGISTERS[5][19] ) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n1747), .CK(net2423), .Q(
        \REGISTERS[4][19] ) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n1746), .CK(net2418), .Q(
        \REGISTERS[3][19] ) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n1745), .CK(net2413), .Q(
        \REGISTERS[2][19] ) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n1744), .CK(net2408), .Q(
        \REGISTERS[1][19] ) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n1743), .CK(net2402), .Q(
        \REGISTERS[0][19] ) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n1742), .CK(net2558), .Q(
        \REGISTERS[31][2] ) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n1741), .CK(net2553), .Q(
        \REGISTERS[30][2] ) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n1740), .CK(net2548), .Q(
        \REGISTERS[29][2] ) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n1739), .CK(net2543), .Q(
        \REGISTERS[28][2] ) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n1738), .CK(net2538), .Q(
        \REGISTERS[27][2] ) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n1737), .CK(net2533), .Q(
        \REGISTERS[26][2] ) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n1736), .CK(net2528), .Q(
        \REGISTERS[25][2] ) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n1735), .CK(net2523), .Q(
        \REGISTERS[24][2] ) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n1734), .CK(net2518), .Q(
        \REGISTERS[23][2] ) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n1733), .CK(net2513), .Q(
        \REGISTERS[22][2] ) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n1732), .CK(net2508), .Q(
        \REGISTERS[21][2] ) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n1731), .CK(net2498), .Q(
        \REGISTERS[19][2] ) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n1730), .CK(net2488), .Q(
        \REGISTERS[17][2] ) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n1729), .CK(net2478), .Q(
        \REGISTERS[15][2] ) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n1728), .CK(net2438), .Q(\REGISTERS[7][2] ) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n1727), .CK(net2433), .Q(\REGISTERS[6][2] ) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n1726), .CK(net2428), .Q(\REGISTERS[5][2] ) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n1725), .CK(net2423), .Q(\REGISTERS[4][2] ) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n1724), .CK(net2418), .Q(\REGISTERS[3][2] ) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n1723), .CK(net2413), .Q(\REGISTERS[2][2] ) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n1722), .CK(net2408), .Q(\REGISTERS[1][2] ) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n1721), .CK(net2402), .Q(\REGISTERS[0][2] ) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n1720), .CK(net2558), .Q(
        \REGISTERS[31][16] ) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n1719), .CK(net2553), .Q(
        \REGISTERS[30][16] ) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n1718), .CK(net2548), .Q(
        \REGISTERS[29][16] ) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n1717), .CK(net2543), .Q(
        \REGISTERS[28][16] ) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n1716), .CK(net2538), .Q(
        \REGISTERS[27][16] ) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n1715), .CK(net2533), .Q(
        \REGISTERS[26][16] ) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n1714), .CK(net2528), .Q(
        \REGISTERS[25][16] ) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n1713), .CK(net2523), .Q(
        \REGISTERS[24][16] ) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n1712), .CK(net2518), .Q(
        \REGISTERS[23][16] ) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n1711), .CK(net2513), .Q(
        \REGISTERS[22][16] ) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n1710), .CK(net2508), .Q(
        \REGISTERS[21][16] ) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n1709), .CK(net2498), .Q(
        \REGISTERS[19][16] ) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n1708), .CK(net2488), .Q(
        \REGISTERS[17][16] ) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n1707), .CK(net2478), .Q(
        \REGISTERS[15][16] ) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n1706), .CK(net2438), .Q(
        \REGISTERS[7][16] ) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n1705), .CK(net2433), .Q(
        \REGISTERS[6][16] ) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n1704), .CK(net2428), .Q(
        \REGISTERS[5][16] ) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n1703), .CK(net2423), .Q(
        \REGISTERS[4][16] ) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n1702), .CK(net2418), .Q(
        \REGISTERS[3][16] ) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n1701), .CK(net2413), .Q(
        \REGISTERS[2][16] ) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n1700), .CK(net2408), .Q(
        \REGISTERS[1][16] ) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n1699), .CK(net2402), .Q(
        \REGISTERS[0][16] ) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n1698), .CK(net2558), .Q(
        \REGISTERS[31][17] ) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n1697), .CK(net2553), .Q(
        \REGISTERS[30][17] ) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n1696), .CK(net2548), .Q(
        \REGISTERS[29][17] ) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n1695), .CK(net2543), .Q(
        \REGISTERS[28][17] ) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n1694), .CK(net2538), .Q(
        \REGISTERS[27][17] ) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n1693), .CK(net2533), .Q(
        \REGISTERS[26][17] ) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n1692), .CK(net2528), .Q(
        \REGISTERS[25][17] ) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n1691), .CK(net2523), .Q(
        \REGISTERS[24][17] ) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n1690), .CK(net2518), .Q(
        \REGISTERS[23][17] ) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n1689), .CK(net2513), .Q(
        \REGISTERS[22][17] ) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n1688), .CK(net2508), .Q(
        \REGISTERS[21][17] ) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n1687), .CK(net2498), .Q(
        \REGISTERS[19][17] ) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n1686), .CK(net2488), .Q(
        \REGISTERS[17][17] ) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n1685), .CK(net2478), .Q(
        \REGISTERS[15][17] ) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n1684), .CK(net2438), .Q(
        \REGISTERS[7][17] ) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n1683), .CK(net2433), .Q(
        \REGISTERS[6][17] ) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n1682), .CK(net2428), .Q(
        \REGISTERS[5][17] ) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n1681), .CK(net2423), .Q(
        \REGISTERS[4][17] ) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n1680), .CK(net2418), .Q(
        \REGISTERS[3][17] ) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n1679), .CK(net2413), .Q(
        \REGISTERS[2][17] ) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n1678), .CK(net2408), .Q(
        \REGISTERS[1][17] ) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n1677), .CK(net2402), .Q(
        \REGISTERS[0][17] ) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n1676), .CK(net2558), .Q(
        \REGISTERS[31][12] ) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n1675), .CK(net2553), .Q(
        \REGISTERS[30][12] ) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n1674), .CK(net2548), .Q(
        \REGISTERS[29][12] ) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n1673), .CK(net2543), .Q(
        \REGISTERS[28][12] ) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n1672), .CK(net2538), .Q(
        \REGISTERS[27][12] ) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n1671), .CK(net2533), .Q(
        \REGISTERS[26][12] ) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n1670), .CK(net2528), .Q(
        \REGISTERS[25][12] ) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n1669), .CK(net2523), .Q(
        \REGISTERS[24][12] ) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n1668), .CK(net2518), .Q(
        \REGISTERS[23][12] ) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n1667), .CK(net2513), .Q(
        \REGISTERS[22][12] ) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n1666), .CK(net2508), .Q(
        \REGISTERS[21][12] ) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n1665), .CK(net2498), .Q(
        \REGISTERS[19][12] ) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n1664), .CK(net2488), .Q(
        \REGISTERS[17][12] ) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n1663), .CK(net2478), .Q(
        \REGISTERS[15][12] ) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n1662), .CK(net2438), .Q(
        \REGISTERS[7][12] ) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n1661), .CK(net2433), .Q(
        \REGISTERS[6][12] ) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n1660), .CK(net2428), .Q(
        \REGISTERS[5][12] ) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n1659), .CK(net2423), .Q(
        \REGISTERS[4][12] ) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n1658), .CK(net2418), .Q(
        \REGISTERS[3][12] ) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n1657), .CK(net2413), .Q(
        \REGISTERS[2][12] ) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n1656), .CK(net2408), .Q(
        \REGISTERS[1][12] ) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n1655), .CK(net2402), .Q(
        \REGISTERS[0][12] ) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n1654), .CK(net2558), .Q(
        \REGISTERS[31][11] ) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n1653), .CK(net2553), .Q(
        \REGISTERS[30][11] ) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n1652), .CK(net2548), .Q(
        \REGISTERS[29][11] ) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n1651), .CK(net2543), .Q(
        \REGISTERS[28][11] ) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n1650), .CK(net2538), .Q(
        \REGISTERS[27][11] ) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n1649), .CK(net2533), .Q(
        \REGISTERS[26][11] ) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n1648), .CK(net2528), .Q(
        \REGISTERS[25][11] ) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n1647), .CK(net2523), .Q(
        \REGISTERS[24][11] ) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n1646), .CK(net2518), .Q(
        \REGISTERS[23][11] ) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n1645), .CK(net2513), .Q(
        \REGISTERS[22][11] ) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n1644), .CK(net2508), .Q(
        \REGISTERS[21][11] ) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n1643), .CK(net2498), .Q(
        \REGISTERS[19][11] ) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n1642), .CK(net2488), .Q(
        \REGISTERS[17][11] ) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n1641), .CK(net2478), .Q(
        \REGISTERS[15][11] ) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n1640), .CK(net2438), .Q(
        \REGISTERS[7][11] ) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n1639), .CK(net2433), .Q(
        \REGISTERS[6][11] ) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n1638), .CK(net2428), .Q(
        \REGISTERS[5][11] ) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n1637), .CK(net2423), .Q(
        \REGISTERS[4][11] ) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n1636), .CK(net2418), .Q(
        \REGISTERS[3][11] ) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n1635), .CK(net2413), .Q(
        \REGISTERS[2][11] ) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n1634), .CK(net2408), .Q(
        \REGISTERS[1][11] ) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n1633), .CK(net2402), .Q(
        \REGISTERS[0][11] ) );
  CLKBUF_X2 U3 ( .A(n1632), .Z(n147) );
  CLKBUF_X2 U4 ( .A(n144), .Z(n146) );
  CLKBUF_X2 U5 ( .A(n152), .Z(n143) );
  CLKBUF_X2 U6 ( .A(n150), .Z(n152) );
  INV_X1 U7 ( .A(n153), .ZN(n1631) );
  INV_X2 U8 ( .A(n1631), .ZN(n1632) );
  CLKBUF_X1 U9 ( .A(n146), .Z(n153) );
  CLKBUF_X2 U10 ( .A(RST), .Z(n138) );
  CLKBUF_X2 U11 ( .A(RST), .Z(n141) );
  CLKBUF_X2 U12 ( .A(RST), .Z(n148) );
  CLKBUF_X2 U13 ( .A(n154), .Z(n142) );
  CLKBUF_X2 U14 ( .A(RST), .Z(n137) );
  CLKBUF_X2 U15 ( .A(RST), .Z(n140) );
  CLKBUF_X2 U16 ( .A(RST), .Z(n155) );
  CLKBUF_X2 U17 ( .A(RST), .Z(n139) );
  CLKBUF_X2 U18 ( .A(RST), .Z(n154) );
  CLKBUF_X2 U19 ( .A(RST), .Z(n144) );
  CLKBUF_X2 U20 ( .A(RST), .Z(n151) );
  CLKBUF_X2 U21 ( .A(n149), .Z(n145) );
  CLKBUF_X2 U22 ( .A(RST), .Z(n150) );
  CLKBUF_X2 U24 ( .A(n156), .Z(n149) );
  CLKBUF_X2 U25 ( .A(RST), .Z(n156) );
  AND2_X1 U26 ( .A1(n113), .A2(RST), .ZN(n1633) );
  AND2_X1 U27 ( .A1(n113), .A2(n156), .ZN(n1634) );
  AND2_X1 U28 ( .A1(n113), .A2(n155), .ZN(n1635) );
  AND2_X1 U29 ( .A1(n113), .A2(n147), .ZN(n1636) );
  AND2_X1 U30 ( .A1(n113), .A2(n1632), .ZN(n1637) );
  AND2_X1 U31 ( .A1(n113), .A2(RST), .ZN(n1638) );
  AND2_X1 U32 ( .A1(n113), .A2(n151), .ZN(n1639) );
  AND2_X1 U33 ( .A1(n113), .A2(RST), .ZN(n1640) );
  AND2_X1 U35 ( .A1(n113), .A2(RST), .ZN(n1641) );
  AND2_X1 U36 ( .A1(n113), .A2(n151), .ZN(n1642) );
  AND2_X1 U37 ( .A1(n113), .A2(RST), .ZN(n1643) );
  AND2_X1 U38 ( .A1(n113), .A2(RST), .ZN(n1644) );
  AND2_X1 U39 ( .A1(n113), .A2(RST), .ZN(n1645) );
  AND2_X1 U40 ( .A1(n113), .A2(n137), .ZN(n1646) );
  AND2_X1 U41 ( .A1(n113), .A2(RST), .ZN(n1647) );
  AND2_X1 U43 ( .A1(n113), .A2(n138), .ZN(n1648) );
  AND2_X1 U44 ( .A1(n113), .A2(RST), .ZN(n1649) );
  AND2_X1 U45 ( .A1(n113), .A2(RST), .ZN(n1650) );
  AND2_X1 U46 ( .A1(n113), .A2(n139), .ZN(n1651) );
  AND2_X1 U47 ( .A1(n113), .A2(n137), .ZN(n1652) );
  AND2_X1 U48 ( .A1(n113), .A2(n147), .ZN(n1653) );
  AND2_X1 U49 ( .A1(n113), .A2(RST), .ZN(n1654) );
  AND2_X1 U51 ( .A1(n111), .A2(RST), .ZN(n1655) );
  AND2_X1 U52 ( .A1(n111), .A2(n156), .ZN(n1656) );
  AND2_X1 U53 ( .A1(n111), .A2(n155), .ZN(n1657) );
  AND2_X1 U54 ( .A1(n111), .A2(RST), .ZN(n1658) );
  AND2_X1 U92 ( .A1(n111), .A2(n1632), .ZN(n1659) );
  AND2_X1 U142 ( .A1(n111), .A2(n143), .ZN(n1660) );
  AND2_X1 U143 ( .A1(n111), .A2(n151), .ZN(n1661) );
  AND2_X1 U144 ( .A1(n111), .A2(n156), .ZN(n1662) );
  AND2_X1 U148 ( .A1(n111), .A2(n146), .ZN(n1663) );
  AND2_X1 U149 ( .A1(n111), .A2(n152), .ZN(n1664) );
  AND2_X1 U150 ( .A1(n111), .A2(RST), .ZN(n1665) );
  AND2_X1 U151 ( .A1(n111), .A2(RST), .ZN(n1666) );
  AND2_X1 U154 ( .A1(n111), .A2(RST), .ZN(n1667) );
  AND2_X1 U155 ( .A1(n111), .A2(n139), .ZN(n1668) );
  AND2_X1 U156 ( .A1(n111), .A2(RST), .ZN(n1669) );
  AND2_X1 U158 ( .A1(n111), .A2(n137), .ZN(n1670) );
  AND2_X1 U160 ( .A1(n111), .A2(n140), .ZN(n1671) );
  AND2_X1 U161 ( .A1(n111), .A2(RST), .ZN(n1672) );
  AND2_X1 U163 ( .A1(n111), .A2(n139), .ZN(n1673) );
  AND2_X1 U164 ( .A1(n111), .A2(n137), .ZN(n1674) );
  AND2_X1 U165 ( .A1(n111), .A2(n142), .ZN(n1675) );
  AND2_X1 U166 ( .A1(n111), .A2(RST), .ZN(n1676) );
  AND2_X1 U904 ( .A1(n101), .A2(RST), .ZN(n1677) );
  AND2_X1 U1662 ( .A1(n101), .A2(n156), .ZN(n1678) );
  AND2_X1 U1731 ( .A1(n101), .A2(n155), .ZN(n1679) );
  AND2_X1 U1732 ( .A1(n101), .A2(RST), .ZN(n1680) );
  AND2_X1 U1733 ( .A1(n101), .A2(n1632), .ZN(n1681) );
  AND2_X1 U1734 ( .A1(n101), .A2(n152), .ZN(n1682) );
  AND2_X1 U1735 ( .A1(n101), .A2(n151), .ZN(n1683) );
  AND2_X1 U1736 ( .A1(n101), .A2(n148), .ZN(n1684) );
  AND2_X1 U1737 ( .A1(n101), .A2(RST), .ZN(n1685) );
  AND2_X1 U1738 ( .A1(n101), .A2(RST), .ZN(n1686) );
  AND2_X1 U1739 ( .A1(n101), .A2(n138), .ZN(n1687) );
  AND2_X1 U1740 ( .A1(n101), .A2(RST), .ZN(n1688) );
  AND2_X1 U1741 ( .A1(n101), .A2(n141), .ZN(n1689) );
  AND2_X1 U1742 ( .A1(n101), .A2(RST), .ZN(n1690) );
  AND2_X1 U1743 ( .A1(n101), .A2(RST), .ZN(n1691) );
  AND2_X1 U1744 ( .A1(n101), .A2(n139), .ZN(n1692) );
  AND2_X1 U1745 ( .A1(n101), .A2(n151), .ZN(n1693) );
  AND2_X1 U1746 ( .A1(n101), .A2(RST), .ZN(n1694) );
  AND2_X1 U1747 ( .A1(n101), .A2(n139), .ZN(n1695) );
  AND2_X1 U1748 ( .A1(n101), .A2(n137), .ZN(n1696) );
  AND2_X1 U1749 ( .A1(n101), .A2(RST), .ZN(n1697) );
  AND2_X1 U1750 ( .A1(n101), .A2(n152), .ZN(n1698) );
  AND2_X1 U1751 ( .A1(n103), .A2(RST), .ZN(n1699) );
  AND2_X1 U1752 ( .A1(n103), .A2(n156), .ZN(n1700) );
  AND2_X1 U1753 ( .A1(n103), .A2(n155), .ZN(n1701) );
  AND2_X1 U1754 ( .A1(n103), .A2(n142), .ZN(n1702) );
  AND2_X1 U1755 ( .A1(n103), .A2(n1632), .ZN(n1703) );
  AND2_X1 U1756 ( .A1(n103), .A2(n146), .ZN(n1704) );
  AND2_X1 U1757 ( .A1(n103), .A2(n151), .ZN(n1705) );
  AND2_X1 U1758 ( .A1(n103), .A2(n148), .ZN(n1706) );
  AND2_X1 U1759 ( .A1(n103), .A2(n154), .ZN(n1707) );
  AND2_X1 U1760 ( .A1(n103), .A2(n149), .ZN(n1708) );
  AND2_X1 U1761 ( .A1(n103), .A2(n139), .ZN(n1709) );
  AND2_X1 U1762 ( .A1(n103), .A2(RST), .ZN(n1710) );
  AND2_X1 U1763 ( .A1(n103), .A2(RST), .ZN(n1711) );
  AND2_X1 U1764 ( .A1(n103), .A2(n141), .ZN(n1712) );
  AND2_X1 U1765 ( .A1(n103), .A2(n141), .ZN(n1713) );
  AND2_X1 U1766 ( .A1(n103), .A2(n140), .ZN(n1714) );
  AND2_X1 U1767 ( .A1(n103), .A2(RST), .ZN(n1715) );
  AND2_X1 U1768 ( .A1(n103), .A2(RST), .ZN(n1716) );
  AND2_X1 U1769 ( .A1(n103), .A2(n139), .ZN(n1717) );
  AND2_X1 U1770 ( .A1(n103), .A2(n137), .ZN(n1718) );
  AND2_X1 U1771 ( .A1(n103), .A2(RST), .ZN(n1719) );
  AND2_X1 U1772 ( .A1(n103), .A2(n143), .ZN(n1720) );
  AND2_X1 U1773 ( .A1(n131), .A2(n155), .ZN(n1721) );
  AND2_X1 U1774 ( .A1(n131), .A2(n145), .ZN(n1722) );
  AND2_X1 U1775 ( .A1(n131), .A2(n154), .ZN(n1723) );
  AND2_X1 U1776 ( .A1(n131), .A2(RST), .ZN(n1724) );
  AND2_X1 U1777 ( .A1(n131), .A2(n152), .ZN(n1725) );
  AND2_X1 U1778 ( .A1(n131), .A2(RST), .ZN(n1726) );
  AND2_X1 U1779 ( .A1(n131), .A2(n150), .ZN(n1727) );
  AND2_X1 U1780 ( .A1(n131), .A2(RST), .ZN(n1728) );
  AND2_X1 U1781 ( .A1(n131), .A2(RST), .ZN(n1729) );
  AND2_X1 U1782 ( .A1(n131), .A2(n140), .ZN(n1730) );
  AND2_X1 U1783 ( .A1(n131), .A2(n152), .ZN(n1731) );
  AND2_X1 U1784 ( .A1(n131), .A2(n139), .ZN(n1732) );
  AND2_X1 U1785 ( .A1(n131), .A2(RST), .ZN(n1733) );
  AND2_X1 U1786 ( .A1(n131), .A2(n141), .ZN(n1734) );
  AND2_X1 U1787 ( .A1(n131), .A2(n145), .ZN(n1735) );
  AND2_X1 U1788 ( .A1(n131), .A2(RST), .ZN(n1736) );
  AND2_X1 U1789 ( .A1(n131), .A2(n141), .ZN(n1737) );
  AND2_X1 U1790 ( .A1(n131), .A2(n140), .ZN(n1738) );
  AND2_X1 U1791 ( .A1(n131), .A2(n138), .ZN(n1739) );
  AND2_X1 U1792 ( .A1(n131), .A2(n142), .ZN(n1740) );
  AND2_X1 U1793 ( .A1(n131), .A2(n143), .ZN(n1741) );
  AND2_X1 U1794 ( .A1(n131), .A2(RST), .ZN(n1742) );
  AND2_X1 U1795 ( .A1(n97), .A2(RST), .ZN(n1743) );
  AND2_X1 U1796 ( .A1(n97), .A2(n156), .ZN(n1744) );
  AND2_X1 U1797 ( .A1(n97), .A2(n155), .ZN(n1745) );
  AND2_X1 U1798 ( .A1(n97), .A2(n155), .ZN(n1746) );
  AND2_X1 U1799 ( .A1(n97), .A2(n1632), .ZN(n1747) );
  AND2_X1 U1800 ( .A1(n97), .A2(n143), .ZN(n1748) );
  AND2_X1 U1801 ( .A1(n97), .A2(n151), .ZN(n1749) );
  AND2_X1 U1802 ( .A1(n97), .A2(n143), .ZN(n1750) );
  AND2_X1 U1803 ( .A1(n97), .A2(n150), .ZN(n1751) );
  AND2_X1 U1804 ( .A1(n97), .A2(n1632), .ZN(n1752) );
  AND2_X1 U1805 ( .A1(n97), .A2(RST), .ZN(n1753) );
  AND2_X1 U1806 ( .A1(n97), .A2(RST), .ZN(n1754) );
  AND2_X1 U1807 ( .A1(n97), .A2(n140), .ZN(n1755) );
  AND2_X1 U1808 ( .A1(n97), .A2(n139), .ZN(n1756) );
  AND2_X1 U1809 ( .A1(n97), .A2(n144), .ZN(n1757) );
  AND2_X1 U1810 ( .A1(n97), .A2(n155), .ZN(n1758) );
  AND2_X1 U1811 ( .A1(n97), .A2(RST), .ZN(n1759) );
  AND2_X1 U1812 ( .A1(n97), .A2(RST), .ZN(n1760) );
  AND2_X1 U1813 ( .A1(n97), .A2(n139), .ZN(n1761) );
  AND2_X1 U1814 ( .A1(n97), .A2(n137), .ZN(n1762) );
  AND2_X1 U1815 ( .A1(n97), .A2(n145), .ZN(n1763) );
  AND2_X1 U1816 ( .A1(n97), .A2(n149), .ZN(n1764) );
  AND2_X1 U1817 ( .A1(n127), .A2(RST), .ZN(n1765) );
  AND2_X1 U1818 ( .A1(n127), .A2(RST), .ZN(n1766) );
  AND2_X1 U1819 ( .A1(n127), .A2(n154), .ZN(n1767) );
  AND2_X1 U1820 ( .A1(n127), .A2(n151), .ZN(n1768) );
  AND2_X1 U1821 ( .A1(n127), .A2(n152), .ZN(n1769) );
  AND2_X1 U1822 ( .A1(n127), .A2(n156), .ZN(n1770) );
  AND2_X1 U1823 ( .A1(n127), .A2(n150), .ZN(n1771) );
  AND2_X1 U1824 ( .A1(n127), .A2(n152), .ZN(n1772) );
  AND2_X1 U1825 ( .A1(n127), .A2(RST), .ZN(n1773) );
  AND2_X1 U1826 ( .A1(n127), .A2(n138), .ZN(n1774) );
  AND2_X1 U1827 ( .A1(n127), .A2(n154), .ZN(n1775) );
  AND2_X1 U1828 ( .A1(n127), .A2(RST), .ZN(n1776) );
  AND2_X1 U1829 ( .A1(n127), .A2(RST), .ZN(n1777) );
  AND2_X1 U1830 ( .A1(n127), .A2(n143), .ZN(n1778) );
  AND2_X1 U1831 ( .A1(n127), .A2(RST), .ZN(n1779) );
  AND2_X1 U1832 ( .A1(n127), .A2(RST), .ZN(n1780) );
  AND2_X1 U1833 ( .A1(n127), .A2(n141), .ZN(n1781) );
  AND2_X1 U1834 ( .A1(n127), .A2(n140), .ZN(n1782) );
  AND2_X1 U1835 ( .A1(n127), .A2(n138), .ZN(n1783) );
  AND2_X1 U1836 ( .A1(n127), .A2(n150), .ZN(n1784) );
  AND2_X1 U1837 ( .A1(n127), .A2(n150), .ZN(n1785) );
  AND2_X1 U1838 ( .A1(n127), .A2(n147), .ZN(n1786) );
  AND2_X1 U1839 ( .A1(n121), .A2(RST), .ZN(n1787) );
  AND2_X1 U1840 ( .A1(n121), .A2(n156), .ZN(n1788) );
  AND2_X1 U1841 ( .A1(n121), .A2(n155), .ZN(n1789) );
  AND2_X1 U1842 ( .A1(n121), .A2(RST), .ZN(n1790) );
  AND2_X1 U1843 ( .A1(n121), .A2(n1632), .ZN(n1791) );
  AND2_X1 U1844 ( .A1(n121), .A2(n156), .ZN(n1792) );
  AND2_X1 U1845 ( .A1(n121), .A2(n151), .ZN(n1793) );
  AND2_X1 U1846 ( .A1(n121), .A2(n1632), .ZN(n1794) );
  AND2_X1 U1847 ( .A1(n121), .A2(n152), .ZN(n1795) );
  AND2_X1 U1848 ( .A1(n121), .A2(n147), .ZN(n1796) );
  AND2_X1 U1849 ( .A1(n121), .A2(n139), .ZN(n1797) );
  AND2_X1 U1850 ( .A1(n121), .A2(n139), .ZN(n1798) );
  AND2_X1 U1851 ( .A1(n121), .A2(n139), .ZN(n1799) );
  AND2_X1 U1852 ( .A1(n121), .A2(n141), .ZN(n1800) );
  AND2_X1 U1853 ( .A1(n121), .A2(n139), .ZN(n1801) );
  AND2_X1 U1854 ( .A1(n121), .A2(RST), .ZN(n1802) );
  AND2_X1 U1855 ( .A1(DATAIN[21]), .A2(n142), .ZN(n1803) );
  AND2_X1 U1856 ( .A1(DATAIN[21]), .A2(n144), .ZN(n1804) );
  AND2_X1 U1857 ( .A1(DATAIN[21]), .A2(n148), .ZN(n1805) );
  AND2_X1 U1858 ( .A1(DATAIN[21]), .A2(n154), .ZN(n1806) );
  AND2_X1 U1859 ( .A1(DATAIN[21]), .A2(n150), .ZN(n1807) );
  AND2_X1 U1860 ( .A1(DATAIN[21]), .A2(n152), .ZN(n1808) );
  AND2_X1 U1861 ( .A1(DATAIN[21]), .A2(RST), .ZN(n1809) );
  AND2_X1 U1862 ( .A1(DATAIN[21]), .A2(n150), .ZN(n1810) );
  AND2_X1 U1863 ( .A1(DATAIN[21]), .A2(n143), .ZN(n1811) );
  AND2_X1 U1864 ( .A1(DATAIN[21]), .A2(RST), .ZN(n1812) );
  AND2_X1 U1865 ( .A1(DATAIN[21]), .A2(n148), .ZN(n1813) );
  AND2_X1 U1866 ( .A1(DATAIN[21]), .A2(RST), .ZN(n1814) );
  AND2_X1 U1867 ( .A1(DATAIN[21]), .A2(n154), .ZN(n1815) );
  AND2_X1 U1868 ( .A1(DATAIN[21]), .A2(n146), .ZN(n1816) );
  AND2_X1 U1869 ( .A1(DATAIN[21]), .A2(n144), .ZN(n1817) );
  AND2_X1 U1870 ( .A1(DATAIN[21]), .A2(n143), .ZN(n1818) );
  AND2_X1 U1871 ( .A1(DATAIN[21]), .A2(RST), .ZN(n1819) );
  AND2_X1 U1872 ( .A1(DATAIN[21]), .A2(n142), .ZN(n1820) );
  AND2_X1 U1873 ( .A1(DATAIN[21]), .A2(RST), .ZN(n1821) );
  AND2_X1 U1874 ( .A1(DATAIN[21]), .A2(n156), .ZN(n1822) );
  AND2_X1 U1875 ( .A1(DATAIN[21]), .A2(n144), .ZN(n1823) );
  AND2_X1 U1876 ( .A1(DATAIN[21]), .A2(RST), .ZN(n1824) );
  AND2_X1 U1877 ( .A1(DATAIN[21]), .A2(n138), .ZN(n1825) );
  AND2_X1 U1878 ( .A1(DATAIN[21]), .A2(RST), .ZN(n1826) );
  AND2_X1 U1879 ( .A1(DATAIN[21]), .A2(n150), .ZN(n1827) );
  AND2_X1 U1880 ( .A1(DATAIN[21]), .A2(n141), .ZN(n1828) );
  AND2_X1 U1881 ( .A1(DATAIN[21]), .A2(n143), .ZN(n1829) );
  AND2_X1 U1882 ( .A1(DATAIN[21]), .A2(n141), .ZN(n1830) );
  AND2_X1 U1883 ( .A1(DATAIN[21]), .A2(n140), .ZN(n1831) );
  AND2_X1 U1884 ( .A1(DATAIN[21]), .A2(n138), .ZN(n1832) );
  AND2_X1 U1885 ( .A1(DATAIN[21]), .A2(RST), .ZN(n1833) );
  AND2_X1 U1886 ( .A1(DATAIN[21]), .A2(RST), .ZN(n1834) );
  AND2_X1 U1887 ( .A1(n85), .A2(n156), .ZN(n1835) );
  AND2_X1 U1888 ( .A1(n85), .A2(n155), .ZN(n1836) );
  AND2_X1 U1889 ( .A1(n85), .A2(n152), .ZN(n1837) );
  AND2_X1 U1890 ( .A1(n85), .A2(n154), .ZN(n1838) );
  AND2_X1 U1891 ( .A1(n85), .A2(n146), .ZN(n1839) );
  AND2_X1 U1892 ( .A1(n85), .A2(n152), .ZN(n1840) );
  AND2_X1 U1893 ( .A1(n85), .A2(RST), .ZN(n1841) );
  AND2_X1 U1894 ( .A1(n85), .A2(n150), .ZN(n1842) );
  AND2_X1 U1895 ( .A1(n85), .A2(n143), .ZN(n1843) );
  AND2_X1 U1896 ( .A1(n85), .A2(n142), .ZN(n1844) );
  AND2_X1 U1897 ( .A1(n85), .A2(RST), .ZN(n1845) );
  AND2_X1 U1898 ( .A1(n85), .A2(RST), .ZN(n1846) );
  AND2_X1 U1899 ( .A1(n85), .A2(RST), .ZN(n1847) );
  AND2_X1 U1900 ( .A1(n85), .A2(n141), .ZN(n1848) );
  AND2_X1 U1901 ( .A1(n85), .A2(n139), .ZN(n1849) );
  AND2_X1 U1902 ( .A1(n85), .A2(n154), .ZN(n1850) );
  AND2_X1 U1903 ( .A1(n85), .A2(n139), .ZN(n1851) );
  AND2_X1 U1904 ( .A1(n85), .A2(n141), .ZN(n1852) );
  AND2_X1 U1905 ( .A1(n85), .A2(n140), .ZN(n1853) );
  AND2_X1 U1906 ( .A1(n85), .A2(n138), .ZN(n1854) );
  AND2_X1 U1907 ( .A1(n85), .A2(RST), .ZN(n1855) );
  AND2_X1 U1908 ( .A1(n85), .A2(n1632), .ZN(n1856) );
  AND2_X1 U1909 ( .A1(n109), .A2(RST), .ZN(n1857) );
  AND2_X1 U1910 ( .A1(n109), .A2(n156), .ZN(n1858) );
  AND2_X1 U1911 ( .A1(n109), .A2(n155), .ZN(n1859) );
  AND2_X1 U1912 ( .A1(n109), .A2(n144), .ZN(n1860) );
  AND2_X1 U1913 ( .A1(n109), .A2(n1632), .ZN(n1861) );
  AND2_X1 U1914 ( .A1(n109), .A2(n145), .ZN(n1862) );
  AND2_X1 U1915 ( .A1(n109), .A2(n151), .ZN(n1863) );
  AND2_X1 U1916 ( .A1(n109), .A2(n155), .ZN(n1864) );
  AND2_X1 U1917 ( .A1(n109), .A2(n143), .ZN(n1865) );
  AND2_X1 U1918 ( .A1(n109), .A2(n142), .ZN(n1866) );
  AND2_X1 U1919 ( .A1(n109), .A2(n141), .ZN(n1867) );
  AND2_X1 U1920 ( .A1(n109), .A2(RST), .ZN(n1868) );
  AND2_X1 U1921 ( .A1(n109), .A2(RST), .ZN(n1869) );
  AND2_X1 U1922 ( .A1(n109), .A2(RST), .ZN(n1870) );
  AND2_X1 U1923 ( .A1(n109), .A2(RST), .ZN(n1871) );
  AND2_X1 U1924 ( .A1(n109), .A2(RST), .ZN(n1872) );
  AND2_X1 U1925 ( .A1(n109), .A2(n151), .ZN(n1873) );
  AND2_X1 U1926 ( .A1(n109), .A2(RST), .ZN(n1874) );
  AND2_X1 U1927 ( .A1(n109), .A2(n139), .ZN(n1875) );
  AND2_X1 U1928 ( .A1(n109), .A2(n137), .ZN(n1876) );
  AND2_X1 U1929 ( .A1(n109), .A2(n156), .ZN(n1877) );
  AND2_X1 U1930 ( .A1(n109), .A2(n145), .ZN(n1878) );
  AND2_X1 U1931 ( .A1(n107), .A2(RST), .ZN(n1879) );
  AND2_X1 U1932 ( .A1(n107), .A2(n156), .ZN(n1880) );
  AND2_X1 U1933 ( .A1(n107), .A2(n155), .ZN(n1881) );
  AND2_X1 U1934 ( .A1(n107), .A2(n151), .ZN(n1882) );
  AND2_X1 U1935 ( .A1(n107), .A2(n1632), .ZN(n1883) );
  AND2_X1 U1936 ( .A1(n107), .A2(n150), .ZN(n1884) );
  AND2_X1 U1937 ( .A1(n107), .A2(n151), .ZN(n1885) );
  AND2_X1 U1938 ( .A1(n107), .A2(RST), .ZN(n1886) );
  AND2_X1 U1939 ( .A1(n107), .A2(n150), .ZN(n1887) );
  AND2_X1 U1940 ( .A1(n107), .A2(n155), .ZN(n1888) );
  AND2_X1 U1941 ( .A1(n107), .A2(RST), .ZN(n1889) );
  AND2_X1 U1942 ( .A1(n107), .A2(RST), .ZN(n1890) );
  AND2_X1 U1943 ( .A1(n107), .A2(RST), .ZN(n1891) );
  AND2_X1 U1944 ( .A1(n107), .A2(RST), .ZN(n1892) );
  AND2_X1 U1945 ( .A1(n107), .A2(RST), .ZN(n1893) );
  AND2_X1 U1946 ( .A1(n107), .A2(n140), .ZN(n1894) );
  AND2_X1 U1947 ( .A1(n107), .A2(n137), .ZN(n1895) );
  AND2_X1 U1948 ( .A1(n107), .A2(RST), .ZN(n1896) );
  AND2_X1 U1949 ( .A1(n107), .A2(n139), .ZN(n1897) );
  AND2_X1 U1950 ( .A1(n107), .A2(n137), .ZN(n1898) );
  AND2_X1 U1951 ( .A1(n107), .A2(n149), .ZN(n1899) );
  AND2_X1 U1952 ( .A1(n107), .A2(RST), .ZN(n1900) );
  AND2_X1 U1953 ( .A1(n99), .A2(RST), .ZN(n1901) );
  AND2_X1 U1954 ( .A1(n99), .A2(n156), .ZN(n1902) );
  AND2_X1 U1955 ( .A1(n99), .A2(n155), .ZN(n1903) );
  AND2_X1 U1956 ( .A1(n99), .A2(n156), .ZN(n1904) );
  AND2_X1 U1957 ( .A1(n99), .A2(n1632), .ZN(n1905) );
  AND2_X1 U1958 ( .A1(n99), .A2(RST), .ZN(n1906) );
  AND2_X1 U1959 ( .A1(n99), .A2(n151), .ZN(n1907) );
  AND2_X1 U1960 ( .A1(n99), .A2(n146), .ZN(n1908) );
  AND2_X1 U1961 ( .A1(n99), .A2(n145), .ZN(n1909) );
  AND2_X1 U1962 ( .A1(n99), .A2(n150), .ZN(n1910) );
  AND2_X1 U1963 ( .A1(n99), .A2(n137), .ZN(n1911) );
  AND2_X1 U1964 ( .A1(n99), .A2(RST), .ZN(n1912) );
  AND2_X1 U1965 ( .A1(n99), .A2(RST), .ZN(n1913) );
  AND2_X1 U1966 ( .A1(n99), .A2(n140), .ZN(n1914) );
  AND2_X1 U1967 ( .A1(n99), .A2(n138), .ZN(n1915) );
  AND2_X1 U1968 ( .A1(n99), .A2(n1632), .ZN(n1916) );
  AND2_X1 U1969 ( .A1(n99), .A2(n155), .ZN(n1917) );
  AND2_X1 U1970 ( .A1(n99), .A2(RST), .ZN(n1918) );
  AND2_X1 U1971 ( .A1(n99), .A2(n139), .ZN(n1919) );
  AND2_X1 U1972 ( .A1(n99), .A2(n137), .ZN(n1920) );
  AND2_X1 U1973 ( .A1(n99), .A2(RST), .ZN(n1921) );
  AND2_X1 U1974 ( .A1(n99), .A2(n150), .ZN(n1922) );
  AND2_X1 U1975 ( .A1(n81), .A2(RST), .ZN(n1923) );
  AND2_X1 U1976 ( .A1(n81), .A2(n146), .ZN(n1924) );
  AND2_X1 U1977 ( .A1(n81), .A2(n155), .ZN(n1925) );
  AND2_X1 U1978 ( .A1(n81), .A2(n154), .ZN(n1926) );
  AND2_X1 U1979 ( .A1(n81), .A2(n146), .ZN(n1927) );
  AND2_X1 U1980 ( .A1(n81), .A2(n152), .ZN(n1928) );
  AND2_X1 U1981 ( .A1(n81), .A2(n145), .ZN(n1929) );
  AND2_X1 U1982 ( .A1(n81), .A2(n150), .ZN(n1930) );
  AND2_X1 U1983 ( .A1(n81), .A2(n143), .ZN(n1931) );
  AND2_X1 U1984 ( .A1(n81), .A2(n142), .ZN(n1932) );
  AND2_X1 U1985 ( .A1(n81), .A2(RST), .ZN(n1933) );
  AND2_X1 U1986 ( .A1(n81), .A2(RST), .ZN(n1934) );
  AND2_X1 U1987 ( .A1(n81), .A2(RST), .ZN(n1935) );
  AND2_X1 U1988 ( .A1(n81), .A2(n140), .ZN(n1936) );
  AND2_X1 U1989 ( .A1(n81), .A2(RST), .ZN(n1937) );
  AND2_X1 U1990 ( .A1(n81), .A2(n140), .ZN(n1938) );
  AND2_X1 U1991 ( .A1(n81), .A2(n137), .ZN(n1939) );
  AND2_X1 U1992 ( .A1(n81), .A2(n141), .ZN(n1940) );
  AND2_X1 U1993 ( .A1(n81), .A2(n140), .ZN(n1941) );
  AND2_X1 U1994 ( .A1(n81), .A2(n138), .ZN(n1942) );
  AND2_X1 U1995 ( .A1(n81), .A2(n155), .ZN(n1943) );
  AND2_X1 U1996 ( .A1(n81), .A2(RST), .ZN(n1944) );
  AND2_X1 U1997 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1945) );
  AND2_X1 U1998 ( .A1(DATAIN[0]), .A2(n154), .ZN(n1946) );
  AND2_X1 U1999 ( .A1(DATAIN[0]), .A2(n154), .ZN(n1947) );
  AND2_X1 U2000 ( .A1(DATAIN[0]), .A2(n148), .ZN(n1948) );
  AND2_X1 U2001 ( .A1(DATAIN[0]), .A2(n152), .ZN(n1949) );
  AND2_X1 U2002 ( .A1(DATAIN[0]), .A2(n154), .ZN(n1950) );
  AND2_X1 U2003 ( .A1(DATAIN[0]), .A2(n150), .ZN(n1951) );
  AND2_X1 U2004 ( .A1(DATAIN[0]), .A2(n148), .ZN(n1952) );
  AND2_X1 U2005 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1953) );
  AND2_X1 U2006 ( .A1(DATAIN[0]), .A2(n148), .ZN(n1954) );
  AND2_X1 U2007 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1955) );
  AND2_X1 U2008 ( .A1(DATAIN[0]), .A2(n149), .ZN(n1956) );
  AND2_X1 U2009 ( .A1(DATAIN[0]), .A2(n146), .ZN(n1957) );
  AND2_X1 U2010 ( .A1(DATAIN[0]), .A2(n144), .ZN(n1958) );
  AND2_X1 U2011 ( .A1(DATAIN[0]), .A2(n143), .ZN(n1959) );
  AND2_X1 U2012 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1960) );
  AND2_X1 U2013 ( .A1(DATAIN[0]), .A2(n142), .ZN(n1961) );
  AND2_X1 U2014 ( .A1(DATAIN[0]), .A2(n141), .ZN(n1962) );
  AND2_X1 U2015 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1963) );
  AND2_X1 U2016 ( .A1(DATAIN[0]), .A2(n148), .ZN(n1964) );
  AND2_X1 U2017 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1965) );
  AND2_X1 U2018 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1966) );
  AND2_X1 U2019 ( .A1(DATAIN[0]), .A2(n137), .ZN(n1967) );
  AND2_X1 U2020 ( .A1(DATAIN[0]), .A2(n152), .ZN(n1968) );
  AND2_X1 U2021 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1969) );
  AND2_X1 U2022 ( .A1(DATAIN[0]), .A2(n138), .ZN(n1970) );
  AND2_X1 U2023 ( .A1(DATAIN[0]), .A2(n141), .ZN(n1971) );
  AND2_X1 U2024 ( .A1(DATAIN[0]), .A2(n140), .ZN(n1972) );
  AND2_X1 U2025 ( .A1(DATAIN[0]), .A2(n138), .ZN(n1973) );
  AND2_X1 U2026 ( .A1(DATAIN[0]), .A2(n148), .ZN(n1974) );
  AND2_X1 U2027 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1975) );
  AND2_X1 U2028 ( .A1(DATAIN[0]), .A2(RST), .ZN(n1976) );
  AND2_X1 U2029 ( .A1(n87), .A2(n154), .ZN(n1977) );
  AND2_X1 U2030 ( .A1(n87), .A2(n142), .ZN(n1978) );
  AND2_X1 U2031 ( .A1(n87), .A2(n151), .ZN(n1979) );
  AND2_X1 U2032 ( .A1(n87), .A2(n154), .ZN(n1980) );
  AND2_X1 U2033 ( .A1(n87), .A2(RST), .ZN(n1981) );
  AND2_X1 U2034 ( .A1(n87), .A2(n152), .ZN(n1982) );
  AND2_X1 U2035 ( .A1(n87), .A2(n147), .ZN(n1983) );
  AND2_X1 U2036 ( .A1(n87), .A2(n150), .ZN(n1984) );
  AND2_X1 U2037 ( .A1(n87), .A2(n143), .ZN(n1985) );
  AND2_X1 U2038 ( .A1(n87), .A2(n142), .ZN(n1986) );
  AND2_X1 U2039 ( .A1(n87), .A2(n143), .ZN(n1987) );
  AND2_X1 U2040 ( .A1(n87), .A2(RST), .ZN(n1988) );
  AND2_X1 U2041 ( .A1(n87), .A2(RST), .ZN(n1989) );
  AND2_X1 U2042 ( .A1(n87), .A2(n141), .ZN(n1990) );
  AND2_X1 U2043 ( .A1(n87), .A2(n140), .ZN(n1991) );
  AND2_X1 U2044 ( .A1(n87), .A2(RST), .ZN(n1992) );
  AND2_X1 U2045 ( .A1(n89), .A2(n150), .ZN(n1993) );
  AND2_X1 U2046 ( .A1(n89), .A2(n152), .ZN(n1994) );
  AND2_X1 U2047 ( .A1(n89), .A2(n144), .ZN(n1995) );
  AND2_X1 U2048 ( .A1(n89), .A2(n154), .ZN(n1996) );
  AND2_X1 U2049 ( .A1(n89), .A2(n154), .ZN(n1997) );
  AND2_X1 U2050 ( .A1(n89), .A2(n152), .ZN(n1998) );
  AND2_X1 U2051 ( .A1(n89), .A2(n148), .ZN(n1999) );
  AND2_X1 U2052 ( .A1(n89), .A2(n150), .ZN(n2000) );
  AND2_X1 U2053 ( .A1(n89), .A2(n143), .ZN(n2001) );
  AND2_X1 U2054 ( .A1(n89), .A2(n142), .ZN(n2002) );
  AND2_X1 U2055 ( .A1(n89), .A2(RST), .ZN(n2003) );
  AND2_X1 U2056 ( .A1(n89), .A2(RST), .ZN(n2004) );
  AND2_X1 U2057 ( .A1(n89), .A2(n156), .ZN(n2005) );
  AND2_X1 U2058 ( .A1(n89), .A2(n146), .ZN(n2006) );
  AND2_X1 U2059 ( .A1(n89), .A2(n140), .ZN(n2007) );
  AND2_X1 U2060 ( .A1(n89), .A2(RST), .ZN(n2008) );
  AND2_X1 U2061 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2009) );
  AND2_X1 U2062 ( .A1(DATAIN[29]), .A2(n150), .ZN(n2010) );
  AND2_X1 U2063 ( .A1(DATAIN[29]), .A2(n143), .ZN(n2011) );
  AND2_X1 U2064 ( .A1(DATAIN[29]), .A2(n154), .ZN(n2012) );
  AND2_X1 U2065 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2013) );
  AND2_X1 U2066 ( .A1(DATAIN[29]), .A2(n152), .ZN(n2014) );
  AND2_X1 U2067 ( .A1(DATAIN[29]), .A2(n151), .ZN(n2015) );
  AND2_X1 U2068 ( .A1(DATAIN[29]), .A2(n150), .ZN(n2016) );
  AND2_X1 U2069 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2017) );
  AND2_X1 U2070 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2018) );
  AND2_X1 U2071 ( .A1(DATAIN[29]), .A2(n148), .ZN(n2019) );
  AND2_X1 U2072 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2020) );
  AND2_X1 U2073 ( .A1(DATAIN[29]), .A2(n146), .ZN(n2021) );
  AND2_X1 U2074 ( .A1(DATAIN[29]), .A2(n146), .ZN(n2022) );
  AND2_X1 U2075 ( .A1(DATAIN[29]), .A2(n144), .ZN(n2023) );
  AND2_X1 U2076 ( .A1(DATAIN[29]), .A2(n143), .ZN(n2024) );
  AND2_X1 U2077 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2025) );
  AND2_X1 U2078 ( .A1(DATAIN[29]), .A2(n142), .ZN(n2026) );
  AND2_X1 U2079 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2027) );
  AND2_X1 U2080 ( .A1(DATAIN[29]), .A2(n143), .ZN(n2028) );
  AND2_X1 U2081 ( .A1(DATAIN[29]), .A2(n145), .ZN(n2029) );
  AND2_X1 U2082 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2030) );
  AND2_X1 U2083 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2031) );
  AND2_X1 U2084 ( .A1(DATAIN[29]), .A2(n138), .ZN(n2032) );
  AND2_X1 U2085 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2033) );
  AND2_X1 U2086 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2034) );
  AND2_X1 U2087 ( .A1(DATAIN[29]), .A2(n140), .ZN(n2035) );
  AND2_X1 U2088 ( .A1(DATAIN[29]), .A2(n141), .ZN(n2036) );
  AND2_X1 U2089 ( .A1(DATAIN[29]), .A2(n140), .ZN(n2037) );
  AND2_X1 U2090 ( .A1(DATAIN[29]), .A2(n138), .ZN(n2038) );
  AND2_X1 U2091 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2039) );
  AND2_X1 U2092 ( .A1(DATAIN[29]), .A2(RST), .ZN(n2040) );
  AND2_X1 U2093 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2041) );
  AND2_X1 U2094 ( .A1(DATAIN[15]), .A2(n156), .ZN(n2042) );
  AND2_X1 U2095 ( .A1(DATAIN[15]), .A2(n155), .ZN(n2043) );
  AND2_X1 U2096 ( .A1(DATAIN[15]), .A2(n152), .ZN(n2044) );
  AND2_X1 U2097 ( .A1(DATAIN[15]), .A2(n1632), .ZN(n2045) );
  AND2_X1 U2098 ( .A1(DATAIN[15]), .A2(n156), .ZN(n2046) );
  AND2_X1 U2099 ( .A1(DATAIN[15]), .A2(n151), .ZN(n2047) );
  AND2_X1 U2100 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2048) );
  AND2_X1 U2101 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2049) );
  AND2_X1 U2102 ( .A1(DATAIN[15]), .A2(n149), .ZN(n2050) );
  AND2_X1 U2103 ( .A1(DATAIN[15]), .A2(n147), .ZN(n2051) );
  AND2_X1 U2104 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2052) );
  AND2_X1 U2105 ( .A1(DATAIN[15]), .A2(n155), .ZN(n2053) );
  AND2_X1 U2106 ( .A1(DATAIN[15]), .A2(n145), .ZN(n2054) );
  AND2_X1 U2107 ( .A1(DATAIN[15]), .A2(n149), .ZN(n2055) );
  AND2_X1 U2108 ( .A1(DATAIN[15]), .A2(n1632), .ZN(n2056) );
  AND2_X1 U2109 ( .A1(DATAIN[15]), .A2(n146), .ZN(n2057) );
  AND2_X1 U2110 ( .A1(DATAIN[15]), .A2(n145), .ZN(n2058) );
  AND2_X1 U2111 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2059) );
  AND2_X1 U2112 ( .A1(DATAIN[15]), .A2(n140), .ZN(n2060) );
  AND2_X1 U2113 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2061) );
  AND2_X1 U2114 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2062) );
  AND2_X1 U2115 ( .A1(DATAIN[15]), .A2(n141), .ZN(n2063) );
  AND2_X1 U2116 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2064) );
  AND2_X1 U2117 ( .A1(DATAIN[15]), .A2(n156), .ZN(n2065) );
  AND2_X1 U2118 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2066) );
  AND2_X1 U2119 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2067) );
  AND2_X1 U2120 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2068) );
  AND2_X1 U2121 ( .A1(DATAIN[15]), .A2(n139), .ZN(n2069) );
  AND2_X1 U2122 ( .A1(DATAIN[15]), .A2(n137), .ZN(n2070) );
  AND2_X1 U2123 ( .A1(DATAIN[15]), .A2(n137), .ZN(n2071) );
  AND2_X1 U2124 ( .A1(DATAIN[15]), .A2(RST), .ZN(n2072) );
  AND2_X1 U2125 ( .A1(DATAIN[10]), .A2(RST), .ZN(n2073) );
  AND2_X1 U2126 ( .A1(DATAIN[10]), .A2(n156), .ZN(n2074) );
  AND2_X1 U2127 ( .A1(DATAIN[10]), .A2(n155), .ZN(n2075) );
  AND2_X1 U2128 ( .A1(DATAIN[10]), .A2(n148), .ZN(n2076) );
  AND2_X1 U2129 ( .A1(DATAIN[10]), .A2(n1632), .ZN(n2077) );
  AND2_X1 U2130 ( .A1(DATAIN[10]), .A2(RST), .ZN(n2078) );
  AND2_X1 U2131 ( .A1(DATAIN[10]), .A2(n151), .ZN(n2079) );
  AND2_X1 U2132 ( .A1(DATAIN[10]), .A2(RST), .ZN(n2080) );
  AND2_X1 U2133 ( .A1(DATAIN[10]), .A2(n144), .ZN(n2081) );
  AND2_X1 U2134 ( .A1(DATAIN[10]), .A2(n149), .ZN(n2082) );
  AND2_X1 U2135 ( .A1(DATAIN[10]), .A2(n147), .ZN(n2083) );
  AND2_X1 U2136 ( .A1(DATAIN[10]), .A2(RST), .ZN(n2084) );
  AND2_X1 U2137 ( .A1(DATAIN[10]), .A2(n154), .ZN(n2085) );
  AND2_X1 U2138 ( .A1(DATAIN[10]), .A2(n145), .ZN(n2086) );
  AND2_X1 U2139 ( .A1(DATAIN[10]), .A2(n143), .ZN(n2087) );
  AND2_X1 U2140 ( .A1(DATAIN[10]), .A2(n149), .ZN(n2088) );
  AND2_X1 U2141 ( .A1(DATAIN[10]), .A2(n142), .ZN(n2089) );
  AND2_X1 U2142 ( .A1(DATAIN[10]), .A2(n144), .ZN(n2090) );
  AND2_X1 U2143 ( .A1(DATAIN[10]), .A2(n149), .ZN(n2091) );
  AND2_X1 U2144 ( .A1(DATAIN[10]), .A2(RST), .ZN(n2092) );
  AND2_X1 U2145 ( .A1(DATAIN[10]), .A2(n150), .ZN(n2093) );
  AND2_X1 U2146 ( .A1(DATAIN[10]), .A2(RST), .ZN(n2094) );
  AND2_X1 U2147 ( .A1(DATAIN[10]), .A2(RST), .ZN(n2095) );
  AND2_X1 U2148 ( .A1(DATAIN[10]), .A2(n137), .ZN(n2096) );
  AND2_X1 U2149 ( .A1(DATAIN[10]), .A2(n137), .ZN(n2097) );
  AND2_X1 U2150 ( .A1(DATAIN[10]), .A2(n139), .ZN(n2098) );
  AND2_X1 U2151 ( .A1(DATAIN[10]), .A2(n137), .ZN(n2099) );
  AND2_X1 U2152 ( .A1(DATAIN[10]), .A2(RST), .ZN(n2100) );
  AND2_X1 U2153 ( .A1(DATAIN[10]), .A2(n139), .ZN(n2101) );
  AND2_X1 U2154 ( .A1(DATAIN[10]), .A2(n137), .ZN(n2102) );
  AND2_X1 U2155 ( .A1(DATAIN[10]), .A2(n148), .ZN(n2103) );
  AND2_X1 U2156 ( .A1(DATAIN[10]), .A2(RST), .ZN(n2104) );
  AND2_X1 U2157 ( .A1(n117), .A2(RST), .ZN(n2105) );
  AND2_X1 U2158 ( .A1(n117), .A2(n156), .ZN(n2106) );
  AND2_X1 U2159 ( .A1(n117), .A2(n155), .ZN(n2107) );
  AND2_X1 U2160 ( .A1(n117), .A2(RST), .ZN(n2108) );
  AND2_X1 U2161 ( .A1(n117), .A2(n1632), .ZN(n2109) );
  AND2_X1 U2162 ( .A1(n117), .A2(RST), .ZN(n2110) );
  AND2_X1 U2163 ( .A1(n117), .A2(n151), .ZN(n2111) );
  AND2_X1 U2164 ( .A1(n117), .A2(n142), .ZN(n2112) );
  AND2_X1 U2165 ( .A1(n117), .A2(n155), .ZN(n2113) );
  AND2_X1 U2166 ( .A1(n117), .A2(RST), .ZN(n2114) );
  AND2_X1 U2167 ( .A1(n117), .A2(n137), .ZN(n2115) );
  AND2_X1 U2168 ( .A1(n117), .A2(RST), .ZN(n2116) );
  AND2_X1 U2169 ( .A1(n117), .A2(n137), .ZN(n2117) );
  AND2_X1 U2170 ( .A1(n117), .A2(n138), .ZN(n2118) );
  AND2_X1 U2171 ( .A1(n117), .A2(n152), .ZN(n2119) );
  AND2_X1 U2172 ( .A1(n117), .A2(n141), .ZN(n2120) );
  AND2_X1 U2173 ( .A1(n117), .A2(n138), .ZN(n2121) );
  AND2_X1 U2174 ( .A1(n117), .A2(RST), .ZN(n2122) );
  AND2_X1 U2175 ( .A1(n117), .A2(n139), .ZN(n2123) );
  AND2_X1 U2176 ( .A1(n117), .A2(n137), .ZN(n2124) );
  AND2_X1 U2177 ( .A1(n117), .A2(RST), .ZN(n2125) );
  AND2_X1 U2178 ( .A1(n117), .A2(n140), .ZN(n2126) );
  AND2_X1 U2179 ( .A1(n95), .A2(RST), .ZN(n2127) );
  AND2_X1 U2180 ( .A1(n83), .A2(RST), .ZN(n2128) );
  AND2_X1 U2181 ( .A1(n95), .A2(n156), .ZN(n2129) );
  AND2_X1 U2182 ( .A1(n83), .A2(RST), .ZN(n2130) );
  AND2_X1 U2183 ( .A1(n95), .A2(n155), .ZN(n2131) );
  AND2_X1 U2184 ( .A1(n83), .A2(n142), .ZN(n2132) );
  AND2_X1 U2185 ( .A1(n95), .A2(RST), .ZN(n2133) );
  AND2_X1 U2186 ( .A1(n83), .A2(n154), .ZN(n2134) );
  AND2_X1 U2187 ( .A1(n95), .A2(n1632), .ZN(n2135) );
  AND2_X1 U2188 ( .A1(n83), .A2(RST), .ZN(n2136) );
  AND2_X1 U2189 ( .A1(n95), .A2(RST), .ZN(n2137) );
  AND2_X1 U2190 ( .A1(n83), .A2(n152), .ZN(n2138) );
  AND2_X1 U2191 ( .A1(n95), .A2(n151), .ZN(n2139) );
  AND2_X1 U2192 ( .A1(n83), .A2(RST), .ZN(n2140) );
  AND2_X1 U2193 ( .A1(n95), .A2(RST), .ZN(n2141) );
  AND2_X1 U2194 ( .A1(n83), .A2(n150), .ZN(n2142) );
  AND2_X1 U2195 ( .A1(n95), .A2(RST), .ZN(n2143) );
  AND2_X1 U2196 ( .A1(n83), .A2(n143), .ZN(n2144) );
  AND2_X1 U2197 ( .A1(n95), .A2(n154), .ZN(n2145) );
  AND2_X1 U2198 ( .A1(n83), .A2(n142), .ZN(n2146) );
  AND2_X1 U2199 ( .A1(n95), .A2(RST), .ZN(n2147) );
  AND2_X1 U2200 ( .A1(n83), .A2(RST), .ZN(n2148) );
  AND2_X1 U2201 ( .A1(n95), .A2(RST), .ZN(n2149) );
  AND2_X1 U2202 ( .A1(n83), .A2(RST), .ZN(n2150) );
  AND2_X1 U2203 ( .A1(n95), .A2(n139), .ZN(n2151) );
  AND2_X1 U2204 ( .A1(n83), .A2(RST), .ZN(n2152) );
  AND2_X1 U2205 ( .A1(n95), .A2(n138), .ZN(n2153) );
  AND2_X1 U2206 ( .A1(n83), .A2(RST), .ZN(n2154) );
  AND2_X1 U2207 ( .A1(n95), .A2(n150), .ZN(n2155) );
  AND2_X1 U2208 ( .A1(n83), .A2(n1632), .ZN(n2156) );
  AND2_X1 U2209 ( .A1(n95), .A2(n151), .ZN(n2157) );
  AND2_X1 U2210 ( .A1(n83), .A2(n149), .ZN(n2158) );
  AND2_X1 U2211 ( .A1(n95), .A2(RST), .ZN(n2159) );
  AND2_X1 U2212 ( .A1(n83), .A2(n138), .ZN(n2160) );
  AND2_X1 U2213 ( .A1(n95), .A2(RST), .ZN(n2161) );
  AND2_X1 U2214 ( .A1(n83), .A2(n141), .ZN(n2162) );
  AND2_X1 U2215 ( .A1(n95), .A2(n139), .ZN(n2163) );
  AND2_X1 U2216 ( .A1(n83), .A2(n140), .ZN(n2164) );
  AND2_X1 U2217 ( .A1(n95), .A2(n137), .ZN(n2165) );
  AND2_X1 U2218 ( .A1(n83), .A2(n138), .ZN(n2166) );
  AND2_X1 U2219 ( .A1(n95), .A2(RST), .ZN(n2167) );
  AND2_X1 U2220 ( .A1(n83), .A2(n151), .ZN(n2168) );
  AND2_X1 U2221 ( .A1(n95), .A2(n156), .ZN(n2169) );
  AND2_X1 U2222 ( .A1(n83), .A2(n156), .ZN(n2170) );
  AND2_X1 U2223 ( .A1(n119), .A2(RST), .ZN(n2171) );
  AND2_X1 U2224 ( .A1(n73), .A2(n149), .ZN(n2172) );
  AND2_X1 U2225 ( .A1(n119), .A2(n156), .ZN(n2173) );
  AND2_X1 U2226 ( .A1(n73), .A2(n154), .ZN(n2174) );
  AND2_X1 U2227 ( .A1(n119), .A2(n155), .ZN(n2175) );
  AND2_X1 U2228 ( .A1(n73), .A2(n1632), .ZN(n2176) );
  AND2_X1 U2229 ( .A1(n119), .A2(n149), .ZN(n2177) );
  AND2_X1 U2230 ( .A1(n73), .A2(n154), .ZN(n2178) );
  AND2_X1 U2231 ( .A1(n119), .A2(n1632), .ZN(n2179) );
  AND2_X1 U2232 ( .A1(n73), .A2(RST), .ZN(n2180) );
  AND2_X1 U2233 ( .A1(n119), .A2(n155), .ZN(n2181) );
  AND2_X1 U2234 ( .A1(n73), .A2(n152), .ZN(n2182) );
  AND2_X1 U2235 ( .A1(n119), .A2(n151), .ZN(n2183) );
  AND2_X1 U2236 ( .A1(n73), .A2(n1632), .ZN(n2184) );
  AND2_X1 U2237 ( .A1(n119), .A2(n154), .ZN(n2185) );
  AND2_X1 U2238 ( .A1(n73), .A2(n150), .ZN(n2186) );
  AND2_X1 U2239 ( .A1(n119), .A2(n142), .ZN(n2187) );
  AND2_X1 U2240 ( .A1(n73), .A2(n143), .ZN(n2188) );
  AND2_X1 U2241 ( .A1(n119), .A2(RST), .ZN(n2189) );
  AND2_X1 U2242 ( .A1(n73), .A2(n142), .ZN(n2190) );
  AND2_X1 U2243 ( .A1(n119), .A2(n138), .ZN(n2191) );
  AND2_X1 U2244 ( .A1(n73), .A2(n146), .ZN(n2192) );
  AND2_X1 U2245 ( .A1(n119), .A2(RST), .ZN(n2193) );
  AND2_X1 U2246 ( .A1(n73), .A2(RST), .ZN(n2194) );
  AND2_X1 U2247 ( .A1(n119), .A2(n138), .ZN(n2195) );
  AND2_X1 U2248 ( .A1(n73), .A2(n141), .ZN(n2196) );
  AND2_X1 U2249 ( .A1(n119), .A2(n139), .ZN(n2197) );
  AND2_X1 U2250 ( .A1(n73), .A2(n138), .ZN(n2198) );
  AND2_X1 U2251 ( .A1(n119), .A2(n146), .ZN(n2199) );
  AND2_X1 U2252 ( .A1(n73), .A2(n149), .ZN(n2200) );
  AND2_X1 U2253 ( .A1(n119), .A2(n145), .ZN(n2201) );
  AND2_X1 U2254 ( .A1(n73), .A2(RST), .ZN(n2202) );
  AND2_X1 U2255 ( .A1(n119), .A2(n139), .ZN(n2203) );
  AND2_X1 U2256 ( .A1(n73), .A2(RST), .ZN(n2204) );
  AND2_X1 U2257 ( .A1(n119), .A2(RST), .ZN(n2205) );
  AND2_X1 U2258 ( .A1(n73), .A2(n141), .ZN(n2206) );
  AND2_X1 U2259 ( .A1(n119), .A2(n139), .ZN(n2207) );
  AND2_X1 U2260 ( .A1(n73), .A2(n140), .ZN(n2208) );
  AND2_X1 U2261 ( .A1(n119), .A2(n137), .ZN(n2209) );
  AND2_X1 U2262 ( .A1(n73), .A2(n138), .ZN(n2210) );
  AND2_X1 U2263 ( .A1(n119), .A2(RST), .ZN(n2211) );
  AND2_X1 U2264 ( .A1(n73), .A2(RST), .ZN(n2212) );
  AND2_X1 U2265 ( .A1(n119), .A2(n1632), .ZN(n2213) );
  AND2_X1 U2266 ( .A1(n73), .A2(n145), .ZN(n2214) );
  AND2_X1 U2267 ( .A1(n123), .A2(RST), .ZN(n2215) );
  AND2_X1 U2268 ( .A1(n123), .A2(n156), .ZN(n2216) );
  AND2_X1 U2269 ( .A1(n123), .A2(n155), .ZN(n2217) );
  AND2_X1 U2270 ( .A1(n123), .A2(n154), .ZN(n2218) );
  AND2_X1 U2271 ( .A1(n123), .A2(n1632), .ZN(n2219) );
  AND2_X1 U2272 ( .A1(n123), .A2(RST), .ZN(n2220) );
  AND2_X1 U2273 ( .A1(n123), .A2(n151), .ZN(n2221) );
  AND2_X1 U2274 ( .A1(n123), .A2(n151), .ZN(n2222) );
  AND2_X1 U2275 ( .A1(n123), .A2(n151), .ZN(n2223) );
  AND2_X1 U2276 ( .A1(n123), .A2(n148), .ZN(n2224) );
  AND2_X1 U2277 ( .A1(n123), .A2(n140), .ZN(n2225) );
  AND2_X1 U2278 ( .A1(n123), .A2(RST), .ZN(n2226) );
  AND2_X1 U2279 ( .A1(n123), .A2(n140), .ZN(n2227) );
  AND2_X1 U2280 ( .A1(n123), .A2(RST), .ZN(n2228) );
  AND2_X1 U2281 ( .A1(n123), .A2(n139), .ZN(n2229) );
  AND2_X1 U2282 ( .A1(n123), .A2(n1632), .ZN(n2230) );
  AND2_X1 U2283 ( .A1(n123), .A2(n154), .ZN(n2231) );
  AND2_X1 U2284 ( .A1(n123), .A2(RST), .ZN(n2232) );
  AND2_X1 U2285 ( .A1(n123), .A2(n139), .ZN(n2233) );
  AND2_X1 U2286 ( .A1(n123), .A2(n137), .ZN(n2234) );
  AND2_X1 U2287 ( .A1(n123), .A2(RST), .ZN(n2235) );
  AND2_X1 U2288 ( .A1(n123), .A2(n146), .ZN(n2236) );
  AND2_X1 U2289 ( .A1(n125), .A2(RST), .ZN(n2237) );
  AND2_X1 U2290 ( .A1(n125), .A2(n156), .ZN(n2238) );
  AND2_X1 U2291 ( .A1(n125), .A2(n155), .ZN(n2239) );
  AND2_X1 U2292 ( .A1(n125), .A2(RST), .ZN(n2240) );
  AND2_X1 U2293 ( .A1(n125), .A2(n1632), .ZN(n2241) );
  AND2_X1 U2294 ( .A1(n125), .A2(RST), .ZN(n2242) );
  AND2_X1 U2295 ( .A1(n125), .A2(n151), .ZN(n2243) );
  AND2_X1 U2296 ( .A1(n125), .A2(n144), .ZN(n2244) );
  AND2_X1 U2297 ( .A1(n125), .A2(n144), .ZN(n2245) );
  AND2_X1 U2298 ( .A1(n125), .A2(n149), .ZN(n2246) );
  AND2_X1 U2299 ( .A1(n125), .A2(RST), .ZN(n2247) );
  AND2_X1 U2300 ( .A1(n125), .A2(RST), .ZN(n2248) );
  AND2_X1 U2301 ( .A1(n125), .A2(n137), .ZN(n2249) );
  AND2_X1 U2302 ( .A1(n125), .A2(RST), .ZN(n2250) );
  AND2_X1 U2303 ( .A1(n125), .A2(n141), .ZN(n2251) );
  AND2_X1 U2304 ( .A1(n125), .A2(n143), .ZN(n2252) );
  AND2_X1 U2305 ( .A1(n125), .A2(n144), .ZN(n2253) );
  AND2_X1 U2306 ( .A1(n125), .A2(RST), .ZN(n2254) );
  AND2_X1 U2307 ( .A1(n125), .A2(n139), .ZN(n2255) );
  AND2_X1 U2308 ( .A1(n125), .A2(n137), .ZN(n2256) );
  AND2_X1 U2309 ( .A1(n125), .A2(n155), .ZN(n2257) );
  AND2_X1 U2310 ( .A1(n125), .A2(n142), .ZN(n2258) );
  AND2_X1 U2311 ( .A1(DATAIN[28]), .A2(n149), .ZN(n2259) );
  AND2_X1 U2312 ( .A1(DATAIN[28]), .A2(n143), .ZN(n2260) );
  AND2_X1 U2313 ( .A1(DATAIN[28]), .A2(n146), .ZN(n2261) );
  AND2_X1 U2314 ( .A1(DATAIN[28]), .A2(n154), .ZN(n2262) );
  AND2_X1 U2315 ( .A1(DATAIN[28]), .A2(n156), .ZN(n2263) );
  AND2_X1 U2316 ( .A1(DATAIN[28]), .A2(n152), .ZN(n2264) );
  AND2_X1 U2317 ( .A1(DATAIN[28]), .A2(n144), .ZN(n2265) );
  AND2_X1 U2318 ( .A1(DATAIN[28]), .A2(n150), .ZN(n2266) );
  AND2_X1 U2319 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2267) );
  AND2_X1 U2320 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2268) );
  AND2_X1 U2321 ( .A1(DATAIN[28]), .A2(n148), .ZN(n2269) );
  AND2_X1 U2322 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2270) );
  AND2_X1 U2323 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2271) );
  AND2_X1 U2324 ( .A1(DATAIN[28]), .A2(n146), .ZN(n2272) );
  AND2_X1 U2325 ( .A1(DATAIN[28]), .A2(n144), .ZN(n2273) );
  AND2_X1 U2326 ( .A1(DATAIN[28]), .A2(n143), .ZN(n2274) );
  AND2_X1 U2327 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2275) );
  AND2_X1 U2328 ( .A1(DATAIN[28]), .A2(n142), .ZN(n2276) );
  AND2_X1 U2329 ( .A1(DATAIN[28]), .A2(n140), .ZN(n2277) );
  AND2_X1 U2330 ( .A1(DATAIN[28]), .A2(n156), .ZN(n2278) );
  AND2_X1 U2331 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2279) );
  AND2_X1 U2332 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2280) );
  AND2_X1 U2333 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2281) );
  AND2_X1 U2334 ( .A1(DATAIN[28]), .A2(n139), .ZN(n2282) );
  AND2_X1 U2335 ( .A1(DATAIN[28]), .A2(n147), .ZN(n2283) );
  AND2_X1 U2336 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2284) );
  AND2_X1 U2337 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2285) );
  AND2_X1 U2338 ( .A1(DATAIN[28]), .A2(n141), .ZN(n2286) );
  AND2_X1 U2339 ( .A1(DATAIN[28]), .A2(n140), .ZN(n2287) );
  AND2_X1 U2340 ( .A1(DATAIN[28]), .A2(n138), .ZN(n2288) );
  AND2_X1 U2341 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2289) );
  AND2_X1 U2342 ( .A1(DATAIN[28]), .A2(RST), .ZN(n2290) );
  AND2_X1 U2343 ( .A1(n129), .A2(RST), .ZN(n2291) );
  AND2_X1 U2344 ( .A1(n91), .A2(n155), .ZN(n2292) );
  AND2_X1 U2345 ( .A1(n129), .A2(n142), .ZN(n2293) );
  AND2_X1 U2346 ( .A1(n91), .A2(n151), .ZN(n2294) );
  AND2_X1 U2347 ( .A1(n129), .A2(n154), .ZN(n2295) );
  AND2_X1 U2348 ( .A1(n91), .A2(n147), .ZN(n2296) );
  AND2_X1 U2349 ( .A1(n129), .A2(n144), .ZN(n2297) );
  AND2_X1 U2350 ( .A1(n91), .A2(n154), .ZN(n2298) );
  AND2_X1 U2351 ( .A1(n129), .A2(n152), .ZN(n2299) );
  AND2_X1 U2352 ( .A1(n91), .A2(n1632), .ZN(n2300) );
  AND2_X1 U2353 ( .A1(n129), .A2(RST), .ZN(n2301) );
  AND2_X1 U2354 ( .A1(n91), .A2(n152), .ZN(n2302) );
  AND2_X1 U2355 ( .A1(n129), .A2(n150), .ZN(n2303) );
  AND2_X1 U2356 ( .A1(n91), .A2(n149), .ZN(n2304) );
  AND2_X1 U2357 ( .A1(n129), .A2(RST), .ZN(n2305) );
  AND2_X1 U2358 ( .A1(n91), .A2(n150), .ZN(n2306) );
  AND2_X1 U2359 ( .A1(n129), .A2(RST), .ZN(n2307) );
  AND2_X1 U2360 ( .A1(n91), .A2(n143), .ZN(n2308) );
  AND2_X1 U2361 ( .A1(n129), .A2(n139), .ZN(n2309) );
  AND2_X1 U2362 ( .A1(n91), .A2(n142), .ZN(n2310) );
  AND2_X1 U2363 ( .A1(n129), .A2(RST), .ZN(n2311) );
  AND2_X1 U2364 ( .A1(n91), .A2(n144), .ZN(n2312) );
  AND2_X1 U2365 ( .A1(n129), .A2(n138), .ZN(n2313) );
  AND2_X1 U2366 ( .A1(n91), .A2(RST), .ZN(n2314) );
  AND2_X1 U2367 ( .A1(n129), .A2(RST), .ZN(n2315) );
  AND2_X1 U2368 ( .A1(n91), .A2(n137), .ZN(n2316) );
  AND2_X1 U2369 ( .A1(n129), .A2(n1632), .ZN(n2317) );
  AND2_X1 U2370 ( .A1(n91), .A2(RST), .ZN(n2318) );
  AND2_X1 U2371 ( .A1(n129), .A2(n146), .ZN(n2319) );
  AND2_X1 U2372 ( .A1(n91), .A2(n154), .ZN(n2320) );
  AND2_X1 U2373 ( .A1(n129), .A2(n151), .ZN(n2321) );
  AND2_X1 U2374 ( .A1(n91), .A2(RST), .ZN(n2322) );
  AND2_X1 U2375 ( .A1(n129), .A2(n141), .ZN(n2323) );
  AND2_X1 U2376 ( .A1(n91), .A2(n1632), .ZN(n2324) );
  AND2_X1 U2377 ( .A1(n129), .A2(n140), .ZN(n2325) );
  AND2_X1 U2378 ( .A1(n91), .A2(n141), .ZN(n2326) );
  AND2_X1 U2379 ( .A1(n129), .A2(n138), .ZN(n2327) );
  AND2_X1 U2380 ( .A1(n91), .A2(n140), .ZN(n2328) );
  AND2_X1 U2381 ( .A1(n129), .A2(n149), .ZN(n2329) );
  AND2_X1 U2382 ( .A1(n91), .A2(n138), .ZN(n2330) );
  AND2_X1 U2383 ( .A1(n129), .A2(n152), .ZN(n2331) );
  AND2_X1 U2384 ( .A1(n91), .A2(n140), .ZN(n2332) );
  AND2_X1 U2385 ( .A1(n129), .A2(n145), .ZN(n2333) );
  AND2_X1 U2386 ( .A1(n91), .A2(n148), .ZN(n2334) );
  AND2_X1 U2387 ( .A1(n133), .A2(n145), .ZN(n2335) );
  AND2_X1 U2388 ( .A1(n133), .A2(RST), .ZN(n2336) );
  AND2_X1 U2389 ( .A1(n133), .A2(n154), .ZN(n2337) );
  AND2_X1 U2390 ( .A1(n133), .A2(n147), .ZN(n2338) );
  AND2_X1 U2391 ( .A1(n133), .A2(n152), .ZN(n2339) );
  AND2_X1 U2392 ( .A1(n133), .A2(n142), .ZN(n2340) );
  AND2_X1 U2393 ( .A1(n133), .A2(n150), .ZN(n2341) );
  AND2_X1 U2394 ( .A1(n133), .A2(n147), .ZN(n2342) );
  AND2_X1 U2395 ( .A1(n133), .A2(RST), .ZN(n2343) );
  AND2_X1 U2396 ( .A1(n133), .A2(RST), .ZN(n2344) );
  AND2_X1 U2397 ( .A1(n133), .A2(n1632), .ZN(n2345) );
  AND2_X1 U2398 ( .A1(n133), .A2(n140), .ZN(n2346) );
  AND2_X1 U2399 ( .A1(n133), .A2(RST), .ZN(n2347) );
  AND2_X1 U2400 ( .A1(n133), .A2(n152), .ZN(n2348) );
  AND2_X1 U2401 ( .A1(n133), .A2(RST), .ZN(n2349) );
  AND2_X1 U2402 ( .A1(n133), .A2(n146), .ZN(n2350) );
  AND2_X1 U2403 ( .A1(n133), .A2(n141), .ZN(n2351) );
  AND2_X1 U2404 ( .A1(n133), .A2(n140), .ZN(n2352) );
  AND2_X1 U2405 ( .A1(n133), .A2(n138), .ZN(n2353) );
  AND2_X1 U2406 ( .A1(n133), .A2(n147), .ZN(n2354) );
  AND2_X1 U2407 ( .A1(n133), .A2(RST), .ZN(n2355) );
  AND2_X1 U2408 ( .A1(n133), .A2(RST), .ZN(n2356) );
  AND2_X1 U2409 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2357) );
  AND2_X1 U2410 ( .A1(DATAIN[30]), .A2(n1632), .ZN(n2358) );
  AND2_X1 U2411 ( .A1(DATAIN[30]), .A2(n150), .ZN(n2359) );
  AND2_X1 U2412 ( .A1(DATAIN[30]), .A2(n154), .ZN(n2360) );
  AND2_X1 U2413 ( .A1(DATAIN[30]), .A2(n149), .ZN(n2361) );
  AND2_X1 U2414 ( .A1(DATAIN[30]), .A2(n152), .ZN(n2362) );
  AND2_X1 U2415 ( .A1(DATAIN[30]), .A2(n152), .ZN(n2363) );
  AND2_X1 U2416 ( .A1(DATAIN[30]), .A2(n150), .ZN(n2364) );
  AND2_X1 U2417 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2365) );
  AND2_X1 U2418 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2366) );
  AND2_X1 U2419 ( .A1(DATAIN[30]), .A2(n148), .ZN(n2367) );
  AND2_X1 U2420 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2368) );
  AND2_X1 U2421 ( .A1(DATAIN[30]), .A2(n143), .ZN(n2369) );
  AND2_X1 U2422 ( .A1(DATAIN[30]), .A2(n146), .ZN(n2370) );
  AND2_X1 U2423 ( .A1(DATAIN[30]), .A2(n144), .ZN(n2371) );
  AND2_X1 U2424 ( .A1(DATAIN[30]), .A2(n143), .ZN(n2372) );
  AND2_X1 U2425 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2373) );
  AND2_X1 U2426 ( .A1(DATAIN[30]), .A2(n142), .ZN(n2374) );
  AND2_X1 U2427 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2375) );
  AND2_X1 U2428 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2376) );
  AND2_X1 U2429 ( .A1(DATAIN[30]), .A2(n143), .ZN(n2377) );
  AND2_X1 U2430 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2378) );
  AND2_X1 U2431 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2379) );
  AND2_X1 U2432 ( .A1(DATAIN[30]), .A2(n137), .ZN(n2380) );
  AND2_X1 U2433 ( .A1(DATAIN[30]), .A2(n148), .ZN(n2381) );
  AND2_X1 U2434 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2382) );
  AND2_X1 U2435 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2383) );
  AND2_X1 U2436 ( .A1(DATAIN[30]), .A2(n141), .ZN(n2384) );
  AND2_X1 U2437 ( .A1(DATAIN[30]), .A2(n140), .ZN(n2385) );
  AND2_X1 U2438 ( .A1(DATAIN[30]), .A2(n138), .ZN(n2386) );
  AND2_X1 U2439 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2387) );
  AND2_X1 U2440 ( .A1(DATAIN[30]), .A2(RST), .ZN(n2388) );
  AND2_X1 U2441 ( .A1(DATAIN[17]), .A2(n156), .ZN(n2389) );
  AND2_X1 U2442 ( .A1(DATAIN[17]), .A2(n149), .ZN(n2390) );
  AND2_X1 U2443 ( .A1(DATAIN[17]), .A2(n147), .ZN(n2391) );
  AND2_X1 U2444 ( .A1(DATAIN[17]), .A2(RST), .ZN(n2392) );
  AND2_X1 U2445 ( .A1(DATAIN[17]), .A2(n150), .ZN(n2393) );
  AND2_X1 U2446 ( .A1(DATAIN[17]), .A2(n145), .ZN(n2394) );
  AND2_X1 U2447 ( .A1(DATAIN[17]), .A2(n147), .ZN(n2395) );
  AND2_X1 U2448 ( .A1(DATAIN[17]), .A2(n150), .ZN(n2396) );
  AND2_X1 U2449 ( .A1(DATAIN[17]), .A2(RST), .ZN(n2397) );
  AND2_X1 U2450 ( .A1(DATAIN[17]), .A2(n148), .ZN(n2398) );
  AND2_X1 U2451 ( .A1(DATAIN[16]), .A2(RST), .ZN(n2399) );
  AND2_X1 U2452 ( .A1(DATAIN[16]), .A2(n149), .ZN(n2400) );
  AND2_X1 U2453 ( .A1(DATAIN[16]), .A2(n147), .ZN(n2401) );
  AND2_X1 U2454 ( .A1(DATAIN[16]), .A2(RST), .ZN(n2402) );
  AND2_X1 U2455 ( .A1(DATAIN[16]), .A2(n155), .ZN(n2403) );
  AND2_X1 U2456 ( .A1(DATAIN[16]), .A2(n145), .ZN(n2404) );
  AND2_X1 U2457 ( .A1(DATAIN[16]), .A2(n148), .ZN(n2405) );
  AND2_X1 U2458 ( .A1(DATAIN[16]), .A2(n143), .ZN(n2406) );
  AND2_X1 U2459 ( .A1(DATAIN[16]), .A2(n145), .ZN(n2407) );
  AND2_X1 U2460 ( .A1(DATAIN[16]), .A2(n151), .ZN(n2408) );
  AND2_X1 U2461 ( .A1(DATAIN[7]), .A2(n147), .ZN(n2409) );
  AND2_X1 U2462 ( .A1(DATAIN[7]), .A2(n149), .ZN(n2410) );
  AND2_X1 U2463 ( .A1(DATAIN[7]), .A2(n147), .ZN(n2411) );
  AND2_X1 U2464 ( .A1(DATAIN[7]), .A2(RST), .ZN(n2412) );
  AND2_X1 U2465 ( .A1(DATAIN[7]), .A2(n150), .ZN(n2413) );
  AND2_X1 U2466 ( .A1(DATAIN[7]), .A2(n145), .ZN(n2414) );
  AND2_X1 U2467 ( .A1(DATAIN[7]), .A2(n147), .ZN(n2415) );
  AND2_X1 U2468 ( .A1(DATAIN[7]), .A2(n144), .ZN(n2416) );
  AND2_X1 U2469 ( .A1(DATAIN[7]), .A2(RST), .ZN(n2417) );
  AND2_X1 U2470 ( .A1(DATAIN[7]), .A2(n148), .ZN(n2418) );
  AND2_X1 U2471 ( .A1(DATAIN[7]), .A2(n141), .ZN(n2419) );
  AND2_X1 U2472 ( .A1(DATAIN[7]), .A2(n140), .ZN(n2420) );
  AND2_X1 U2473 ( .A1(DATAIN[7]), .A2(n146), .ZN(n2421) );
  AND2_X1 U2474 ( .A1(DATAIN[7]), .A2(RST), .ZN(n2422) );
  AND2_X1 U2475 ( .A1(DATAIN[7]), .A2(n137), .ZN(n2423) );
  AND2_X1 U2476 ( .A1(DATAIN[7]), .A2(n146), .ZN(n2424) );
  AND2_X1 U2477 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2425) );
  AND2_X1 U2478 ( .A1(DATAIN[2]), .A2(n148), .ZN(n2426) );
  AND2_X1 U2479 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2427) );
  AND2_X1 U2480 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2428) );
  AND2_X1 U2481 ( .A1(DATAIN[2]), .A2(n146), .ZN(n2429) );
  AND2_X1 U2482 ( .A1(DATAIN[2]), .A2(n144), .ZN(n2430) );
  AND2_X1 U2483 ( .A1(DATAIN[2]), .A2(n143), .ZN(n2431) );
  AND2_X1 U2484 ( .A1(DATAIN[2]), .A2(n142), .ZN(n2432) );
  AND2_X1 U2485 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2433) );
  AND2_X1 U2486 ( .A1(DATAIN[2]), .A2(RST), .ZN(n2434) );
  AND2_X1 U2487 ( .A1(DATAIN[12]), .A2(n152), .ZN(n2435) );
  AND2_X1 U2488 ( .A1(DATAIN[12]), .A2(n149), .ZN(n2436) );
  AND2_X1 U2489 ( .A1(DATAIN[12]), .A2(n147), .ZN(n2437) );
  AND2_X1 U2490 ( .A1(DATAIN[12]), .A2(RST), .ZN(n2438) );
  AND2_X1 U2491 ( .A1(DATAIN[12]), .A2(RST), .ZN(n2439) );
  AND2_X1 U2492 ( .A1(DATAIN[12]), .A2(n145), .ZN(n2440) );
  AND2_X1 U2493 ( .A1(DATAIN[12]), .A2(RST), .ZN(n2441) );
  AND2_X1 U2494 ( .A1(DATAIN[12]), .A2(RST), .ZN(n2442) );
  AND2_X1 U2495 ( .A1(DATAIN[12]), .A2(n138), .ZN(n2443) );
  AND2_X1 U2496 ( .A1(DATAIN[12]), .A2(n147), .ZN(n2444) );
  AND2_X1 U2497 ( .A1(DATAIN[11]), .A2(n151), .ZN(n2445) );
  AND2_X1 U2498 ( .A1(DATAIN[11]), .A2(n149), .ZN(n2446) );
  AND2_X1 U2499 ( .A1(DATAIN[11]), .A2(n147), .ZN(n2447) );
  AND2_X1 U2500 ( .A1(DATAIN[11]), .A2(RST), .ZN(n2448) );
  AND2_X1 U2501 ( .A1(DATAIN[11]), .A2(n142), .ZN(n2449) );
  AND2_X1 U2502 ( .A1(DATAIN[11]), .A2(n145), .ZN(n2450) );
  AND2_X1 U2503 ( .A1(DATAIN[11]), .A2(RST), .ZN(n2451) );
  AND2_X1 U2504 ( .A1(DATAIN[11]), .A2(n155), .ZN(n2452) );
  AND2_X1 U2505 ( .A1(DATAIN[11]), .A2(RST), .ZN(n2453) );
  AND2_X1 U2506 ( .A1(DATAIN[11]), .A2(n145), .ZN(n2454) );
  AND2_X1 U2507 ( .A1(DATAIN[4]), .A2(RST), .ZN(n2455) );
  AND2_X1 U2508 ( .A1(DATAIN[4]), .A2(n148), .ZN(n2456) );
  AND2_X1 U2509 ( .A1(DATAIN[4]), .A2(RST), .ZN(n2457) );
  AND2_X1 U2510 ( .A1(DATAIN[4]), .A2(n152), .ZN(n2458) );
  AND2_X1 U2511 ( .A1(DATAIN[4]), .A2(n146), .ZN(n2459) );
  AND2_X1 U2512 ( .A1(DATAIN[4]), .A2(n144), .ZN(n2460) );
  AND2_X1 U2513 ( .A1(DATAIN[4]), .A2(n143), .ZN(n2461) );
  AND2_X1 U2514 ( .A1(DATAIN[4]), .A2(n142), .ZN(n2462) );
  AND2_X1 U2515 ( .A1(DATAIN[4]), .A2(RST), .ZN(n2463) );
  AND2_X1 U2516 ( .A1(DATAIN[4]), .A2(RST), .ZN(n2464) );
  AND2_X1 U2517 ( .A1(DATAIN[19]), .A2(RST), .ZN(n2465) );
  AND2_X1 U2518 ( .A1(DATAIN[19]), .A2(n149), .ZN(n2466) );
  AND2_X1 U2519 ( .A1(DATAIN[19]), .A2(n147), .ZN(n2467) );
  AND2_X1 U2520 ( .A1(DATAIN[19]), .A2(RST), .ZN(n2468) );
  AND2_X1 U2521 ( .A1(DATAIN[19]), .A2(n149), .ZN(n2469) );
  AND2_X1 U2522 ( .A1(DATAIN[19]), .A2(n145), .ZN(n2470) );
  AND2_X1 U2523 ( .A1(DATAIN[19]), .A2(RST), .ZN(n2471) );
  AND2_X1 U2524 ( .A1(DATAIN[19]), .A2(n154), .ZN(n2472) );
  AND2_X1 U2525 ( .A1(DATAIN[19]), .A2(n145), .ZN(n2473) );
  AND2_X1 U2526 ( .A1(DATAIN[19]), .A2(n145), .ZN(n2474) );
  AND2_X1 U2527 ( .A1(DATAIN[14]), .A2(n142), .ZN(n2475) );
  AND2_X1 U2528 ( .A1(DATAIN[14]), .A2(n149), .ZN(n2476) );
  AND2_X1 U2529 ( .A1(DATAIN[14]), .A2(n147), .ZN(n2477) );
  AND2_X1 U2530 ( .A1(DATAIN[14]), .A2(RST), .ZN(n2478) );
  AND2_X1 U2531 ( .A1(DATAIN[14]), .A2(n156), .ZN(n2479) );
  AND2_X1 U2532 ( .A1(DATAIN[14]), .A2(n145), .ZN(n2480) );
  AND2_X1 U2533 ( .A1(DATAIN[14]), .A2(RST), .ZN(n2481) );
  AND2_X1 U2534 ( .A1(DATAIN[14]), .A2(RST), .ZN(n2482) );
  AND2_X1 U2535 ( .A1(DATAIN[14]), .A2(n138), .ZN(n2483) );
  AND2_X1 U2536 ( .A1(DATAIN[14]), .A2(RST), .ZN(n2484) );
  AND2_X1 U2537 ( .A1(DATAIN[27]), .A2(n142), .ZN(n2485) );
  AND2_X1 U2538 ( .A1(DATAIN[27]), .A2(RST), .ZN(n2486) );
  AND2_X1 U2539 ( .A1(DATAIN[27]), .A2(n148), .ZN(n2487) );
  AND2_X1 U2540 ( .A1(DATAIN[27]), .A2(RST), .ZN(n2488) );
  AND2_X1 U2541 ( .A1(DATAIN[27]), .A2(RST), .ZN(n2489) );
  AND2_X1 U2542 ( .A1(DATAIN[27]), .A2(n146), .ZN(n2490) );
  AND2_X1 U2543 ( .A1(DATAIN[27]), .A2(n144), .ZN(n2491) );
  AND2_X1 U2544 ( .A1(DATAIN[27]), .A2(RST), .ZN(n2492) );
  AND2_X1 U2545 ( .A1(DATAIN[27]), .A2(n137), .ZN(n2493) );
  AND2_X1 U2546 ( .A1(DATAIN[27]), .A2(RST), .ZN(n2494) );
  AND2_X1 U2547 ( .A1(DATAIN[25]), .A2(n156), .ZN(n2495) );
  AND2_X1 U2548 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2496) );
  AND2_X1 U2549 ( .A1(DATAIN[25]), .A2(n148), .ZN(n2497) );
  AND2_X1 U2550 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2498) );
  AND2_X1 U2551 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2499) );
  AND2_X1 U2552 ( .A1(DATAIN[25]), .A2(n146), .ZN(n2500) );
  AND2_X1 U2553 ( .A1(DATAIN[25]), .A2(n144), .ZN(n2501) );
  AND2_X1 U2554 ( .A1(DATAIN[25]), .A2(RST), .ZN(n2502) );
  AND2_X1 U2555 ( .A1(DATAIN[25]), .A2(n139), .ZN(n2503) );
  AND2_X1 U2556 ( .A1(DATAIN[25]), .A2(n141), .ZN(n2504) );
  AND2_X1 U2557 ( .A1(DATAIN[9]), .A2(RST), .ZN(n2505) );
  AND2_X1 U2558 ( .A1(DATAIN[9]), .A2(n149), .ZN(n2506) );
  AND2_X1 U2559 ( .A1(DATAIN[9]), .A2(n147), .ZN(n2507) );
  AND2_X1 U2560 ( .A1(DATAIN[9]), .A2(RST), .ZN(n2508) );
  AND2_X1 U2561 ( .A1(DATAIN[9]), .A2(n1632), .ZN(n2509) );
  AND2_X1 U2562 ( .A1(DATAIN[9]), .A2(n145), .ZN(n2510) );
  AND2_X1 U2563 ( .A1(DATAIN[9]), .A2(n146), .ZN(n2511) );
  AND2_X1 U2564 ( .A1(DATAIN[9]), .A2(n152), .ZN(n2512) );
  AND2_X1 U2565 ( .A1(DATAIN[9]), .A2(RST), .ZN(n2513) );
  AND2_X1 U2566 ( .A1(DATAIN[9]), .A2(n146), .ZN(n2514) );
  AND2_X1 U2567 ( .A1(DATAIN[13]), .A2(n1632), .ZN(n2515) );
  AND2_X1 U2568 ( .A1(DATAIN[13]), .A2(n149), .ZN(n2516) );
  AND2_X1 U2569 ( .A1(DATAIN[13]), .A2(n147), .ZN(n2517) );
  AND2_X1 U2570 ( .A1(DATAIN[13]), .A2(RST), .ZN(n2518) );
  AND2_X1 U2571 ( .A1(DATAIN[13]), .A2(RST), .ZN(n2519) );
  AND2_X1 U2572 ( .A1(DATAIN[13]), .A2(n145), .ZN(n2520) );
  AND2_X1 U2573 ( .A1(DATAIN[13]), .A2(RST), .ZN(n2521) );
  AND2_X1 U2574 ( .A1(DATAIN[13]), .A2(RST), .ZN(n2522) );
  AND2_X1 U2575 ( .A1(DATAIN[13]), .A2(n1632), .ZN(n2523) );
  AND2_X1 U2576 ( .A1(DATAIN[13]), .A2(n141), .ZN(n2524) );
  AND2_X1 U2577 ( .A1(DATAIN[8]), .A2(RST), .ZN(n2525) );
  AND2_X1 U2578 ( .A1(DATAIN[31]), .A2(RST), .ZN(n2526) );
  AND2_X1 U2579 ( .A1(DATAIN[8]), .A2(n149), .ZN(n2527) );
  AND2_X1 U2580 ( .A1(DATAIN[31]), .A2(RST), .ZN(n2528) );
  AND2_X1 U2581 ( .A1(DATAIN[8]), .A2(n147), .ZN(n2529) );
  AND2_X1 U2582 ( .A1(DATAIN[31]), .A2(n148), .ZN(n2530) );
  AND2_X1 U2583 ( .A1(DATAIN[8]), .A2(RST), .ZN(n2531) );
  AND2_X1 U2584 ( .A1(DATAIN[31]), .A2(RST), .ZN(n2532) );
  AND2_X1 U2585 ( .A1(DATAIN[8]), .A2(n152), .ZN(n2533) );
  AND2_X1 U2586 ( .A1(DATAIN[31]), .A2(RST), .ZN(n2534) );
  AND2_X1 U2587 ( .A1(DATAIN[8]), .A2(n145), .ZN(n2535) );
  AND2_X1 U2588 ( .A1(DATAIN[31]), .A2(n146), .ZN(n2536) );
  AND2_X1 U2589 ( .A1(DATAIN[8]), .A2(n147), .ZN(n2537) );
  AND2_X1 U2590 ( .A1(DATAIN[31]), .A2(n144), .ZN(n2538) );
  AND2_X1 U2591 ( .A1(DATAIN[8]), .A2(n151), .ZN(n2539) );
  AND2_X1 U2592 ( .A1(DATAIN[31]), .A2(RST), .ZN(n2540) );
  AND2_X1 U2593 ( .A1(DATAIN[8]), .A2(RST), .ZN(n2541) );
  AND2_X1 U2594 ( .A1(DATAIN[31]), .A2(RST), .ZN(n2542) );
  AND2_X1 U2595 ( .A1(DATAIN[8]), .A2(n147), .ZN(n2543) );
  AND2_X1 U2596 ( .A1(DATAIN[31]), .A2(RST), .ZN(n2544) );
  AND2_X1 U2597 ( .A1(DATAIN[18]), .A2(n155), .ZN(n2545) );
  AND2_X1 U2598 ( .A1(DATAIN[18]), .A2(n149), .ZN(n2546) );
  AND2_X1 U2599 ( .A1(DATAIN[18]), .A2(n147), .ZN(n2547) );
  AND2_X1 U2600 ( .A1(DATAIN[18]), .A2(RST), .ZN(n2548) );
  AND2_X1 U2601 ( .A1(DATAIN[18]), .A2(RST), .ZN(n2549) );
  AND2_X1 U2602 ( .A1(DATAIN[18]), .A2(n145), .ZN(n2550) );
  AND2_X1 U2603 ( .A1(DATAIN[18]), .A2(RST), .ZN(n2551) );
  AND2_X1 U2604 ( .A1(DATAIN[18]), .A2(n1632), .ZN(n2552) );
  AND2_X1 U2605 ( .A1(DATAIN[18]), .A2(n149), .ZN(n2553) );
  AND2_X1 U2606 ( .A1(DATAIN[18]), .A2(RST), .ZN(n2554) );
  AND2_X1 U2607 ( .A1(DATAIN[5]), .A2(n149), .ZN(n2555) );
  AND2_X1 U2608 ( .A1(DATAIN[5]), .A2(n149), .ZN(n2556) );
  AND2_X1 U2609 ( .A1(DATAIN[5]), .A2(n147), .ZN(n2557) );
  AND2_X1 U2610 ( .A1(DATAIN[5]), .A2(RST), .ZN(n2558) );
  AND2_X1 U2611 ( .A1(DATAIN[5]), .A2(n144), .ZN(n2559) );
  AND2_X1 U2612 ( .A1(DATAIN[5]), .A2(n145), .ZN(n2560) );
  AND2_X1 U2613 ( .A1(DATAIN[5]), .A2(n156), .ZN(n2561) );
  AND2_X1 U2614 ( .A1(DATAIN[5]), .A2(n148), .ZN(n2562) );
  AND2_X1 U2615 ( .A1(DATAIN[5]), .A2(n145), .ZN(n2563) );
  AND2_X1 U2616 ( .A1(DATAIN[5]), .A2(n143), .ZN(n2564) );
  AND2_X1 U2617 ( .A1(DATAIN[1]), .A2(RST), .ZN(n2565) );
  AND2_X1 U2618 ( .A1(DATAIN[1]), .A2(n148), .ZN(n2566) );
  AND2_X1 U2619 ( .A1(DATAIN[1]), .A2(RST), .ZN(n2567) );
  AND2_X1 U2620 ( .A1(DATAIN[1]), .A2(RST), .ZN(n2568) );
  AND2_X1 U2621 ( .A1(DATAIN[1]), .A2(n146), .ZN(n2569) );
  AND2_X1 U2622 ( .A1(DATAIN[1]), .A2(n144), .ZN(n2570) );
  AND2_X1 U2623 ( .A1(DATAIN[1]), .A2(n143), .ZN(n2571) );
  AND2_X1 U2624 ( .A1(DATAIN[1]), .A2(n142), .ZN(n2572) );
  AND2_X1 U2625 ( .A1(DATAIN[1]), .A2(n144), .ZN(n2573) );
  AND2_X1 U2626 ( .A1(DATAIN[1]), .A2(RST), .ZN(n2574) );
  AND2_X1 U2627 ( .A1(DATAIN[3]), .A2(RST), .ZN(n2575) );
  AND2_X1 U2628 ( .A1(DATAIN[22]), .A2(RST), .ZN(n2576) );
  AND2_X1 U2629 ( .A1(DATAIN[3]), .A2(n148), .ZN(n2577) );
  AND2_X1 U2630 ( .A1(DATAIN[22]), .A2(RST), .ZN(n2578) );
  AND2_X1 U2631 ( .A1(DATAIN[3]), .A2(RST), .ZN(n2579) );
  AND2_X1 U2632 ( .A1(DATAIN[22]), .A2(n148), .ZN(n2580) );
  AND2_X1 U2633 ( .A1(DATAIN[3]), .A2(n144), .ZN(n2581) );
  AND2_X1 U2634 ( .A1(DATAIN[22]), .A2(RST), .ZN(n2582) );
  AND2_X1 U2635 ( .A1(DATAIN[3]), .A2(n146), .ZN(n2583) );
  AND2_X1 U2636 ( .A1(DATAIN[22]), .A2(RST), .ZN(n2584) );
  AND2_X1 U2637 ( .A1(DATAIN[3]), .A2(n144), .ZN(n2585) );
  AND2_X1 U2638 ( .A1(DATAIN[22]), .A2(n146), .ZN(n2586) );
  AND2_X1 U2639 ( .A1(DATAIN[3]), .A2(n143), .ZN(n2587) );
  AND2_X1 U2640 ( .A1(DATAIN[22]), .A2(n144), .ZN(n2588) );
  AND2_X1 U2641 ( .A1(DATAIN[3]), .A2(n142), .ZN(n2589) );
  AND2_X1 U2642 ( .A1(DATAIN[22]), .A2(RST), .ZN(n2590) );
  AND2_X1 U2643 ( .A1(DATAIN[3]), .A2(RST), .ZN(n2591) );
  AND2_X1 U2644 ( .A1(DATAIN[22]), .A2(n141), .ZN(n2592) );
  AND2_X1 U2645 ( .A1(DATAIN[3]), .A2(RST), .ZN(n2593) );
  AND2_X1 U2646 ( .A1(DATAIN[22]), .A2(RST), .ZN(n2594) );
  AND2_X1 U2647 ( .A1(DATAIN[6]), .A2(RST), .ZN(n2595) );
  AND2_X1 U2648 ( .A1(DATAIN[6]), .A2(n149), .ZN(n2596) );
  AND2_X1 U2649 ( .A1(DATAIN[6]), .A2(n147), .ZN(n2597) );
  AND2_X1 U2650 ( .A1(DATAIN[6]), .A2(RST), .ZN(n2598) );
  AND2_X1 U2651 ( .A1(DATAIN[6]), .A2(n151), .ZN(n2599) );
  AND2_X1 U2652 ( .A1(DATAIN[6]), .A2(n145), .ZN(n2600) );
  AND2_X1 U2653 ( .A1(DATAIN[6]), .A2(n156), .ZN(n2601) );
  AND2_X1 U2654 ( .A1(DATAIN[6]), .A2(n147), .ZN(n2602) );
  AND2_X1 U2655 ( .A1(DATAIN[6]), .A2(n155), .ZN(n2603) );
  AND2_X1 U2656 ( .A1(DATAIN[6]), .A2(n152), .ZN(n2604) );
  AND2_X1 U2657 ( .A1(DATAIN[26]), .A2(n148), .ZN(n2605) );
  AND2_X1 U2658 ( .A1(DATAIN[26]), .A2(RST), .ZN(n2606) );
  AND2_X1 U2659 ( .A1(DATAIN[26]), .A2(n148), .ZN(n2607) );
  AND2_X1 U2660 ( .A1(DATAIN[26]), .A2(RST), .ZN(n2608) );
  AND2_X1 U2661 ( .A1(DATAIN[26]), .A2(RST), .ZN(n2609) );
  AND2_X1 U2662 ( .A1(DATAIN[26]), .A2(n146), .ZN(n2610) );
  AND2_X1 U2663 ( .A1(DATAIN[26]), .A2(n144), .ZN(n2611) );
  AND2_X1 U2664 ( .A1(DATAIN[26]), .A2(RST), .ZN(n2612) );
  AND2_X1 U2665 ( .A1(DATAIN[26]), .A2(n138), .ZN(n2613) );
  AND2_X1 U2666 ( .A1(DATAIN[26]), .A2(RST), .ZN(n2614) );
  AND2_X1 U2667 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2615) );
  AND2_X1 U2668 ( .A1(DATAIN[20]), .A2(n149), .ZN(n2616) );
  AND2_X1 U2669 ( .A1(DATAIN[20]), .A2(n147), .ZN(n2617) );
  AND2_X1 U2670 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2618) );
  AND2_X1 U2671 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2619) );
  AND2_X1 U2672 ( .A1(DATAIN[20]), .A2(n145), .ZN(n2620) );
  AND2_X1 U2673 ( .A1(DATAIN[20]), .A2(n145), .ZN(n2621) );
  AND2_X1 U2674 ( .A1(DATAIN[20]), .A2(RST), .ZN(n2622) );
  AND2_X1 U2675 ( .A1(DATAIN[20]), .A2(n142), .ZN(n2623) );
  AND2_X1 U2676 ( .A1(DATAIN[20]), .A2(n150), .ZN(n2624) );
  AND2_X1 U2677 ( .A1(DATAIN[24]), .A2(n150), .ZN(n2625) );
  AND2_X1 U2678 ( .A1(DATAIN[24]), .A2(RST), .ZN(n2626) );
  AND2_X1 U2679 ( .A1(DATAIN[24]), .A2(n148), .ZN(n2627) );
  AND2_X1 U2680 ( .A1(DATAIN[24]), .A2(RST), .ZN(n2628) );
  AND2_X1 U2681 ( .A1(DATAIN[24]), .A2(RST), .ZN(n2629) );
  AND2_X1 U2682 ( .A1(DATAIN[24]), .A2(n146), .ZN(n2630) );
  AND2_X1 U2683 ( .A1(DATAIN[24]), .A2(n144), .ZN(n2631) );
  AND2_X1 U2684 ( .A1(DATAIN[24]), .A2(RST), .ZN(n2632) );
  AND2_X1 U2685 ( .A1(DATAIN[24]), .A2(n140), .ZN(n2633) );
  AND2_X1 U2686 ( .A1(DATAIN[24]), .A2(n143), .ZN(n2634) );
  AND2_X1 U2687 ( .A1(DATAIN[24]), .A2(RST), .ZN(n2635) );
  AND2_X1 U2688 ( .A1(DATAIN[24]), .A2(n137), .ZN(n2636) );
  AND2_X1 U2689 ( .A1(DATAIN[24]), .A2(n137), .ZN(n2637) );
  AND2_X1 U2690 ( .A1(DATAIN[24]), .A2(n141), .ZN(n2638) );
  AND2_X1 U2691 ( .A1(DATAIN[24]), .A2(n138), .ZN(n2639) );
  AND2_X1 U2692 ( .A1(DATAIN[24]), .A2(n142), .ZN(n2640) );
  AND2_X1 U2693 ( .A1(DATAIN[23]), .A2(n145), .ZN(n2641) );
  AND2_X1 U2694 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2642) );
  AND2_X1 U2695 ( .A1(DATAIN[23]), .A2(n148), .ZN(n2643) );
  AND2_X1 U2696 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2644) );
  AND2_X1 U2697 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2645) );
  AND2_X1 U2698 ( .A1(DATAIN[23]), .A2(n146), .ZN(n2646) );
  AND2_X1 U2699 ( .A1(DATAIN[23]), .A2(n144), .ZN(n2647) );
  AND2_X1 U2700 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2648) );
  AND2_X1 U2701 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2649) );
  AND2_X1 U2702 ( .A1(DATAIN[23]), .A2(n154), .ZN(n2650) );
  AND2_X1 U2703 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2651) );
  AND2_X1 U2704 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2652) );
  AND2_X1 U2705 ( .A1(DATAIN[23]), .A2(RST), .ZN(n2653) );
  AND2_X1 U2706 ( .A1(DATAIN[23]), .A2(n141), .ZN(n2654) );
  AND2_X1 U2707 ( .A1(DATAIN[23]), .A2(n138), .ZN(n2655) );
  AND2_X1 U2708 ( .A1(DATAIN[23]), .A2(n147), .ZN(n2656) );
  INV_X2 U2709 ( .A(DATAIN[29]), .ZN(n2665) );
  INV_X2 U2710 ( .A(DATAIN[30]), .ZN(n2664) );
  INV_X2 U2711 ( .A(DATAIN[10]), .ZN(n2661) );
  INV_X2 U2712 ( .A(DATAIN[15]), .ZN(n2658) );
  BUF_X2 U2713 ( .A(n82), .Z(n2657) );
  INV_X4 U2714 ( .A(n126), .ZN(n125) );
  BUF_X2 U2715 ( .A(n124), .Z(n2659) );
  BUF_X2 U2716 ( .A(n108), .Z(n2660) );
  INV_X1 U2717 ( .A(DATAIN[2]), .ZN(n132) );
  INV_X1 U2718 ( .A(DATAIN[3]), .ZN(n130) );
  INV_X1 U2719 ( .A(DATAIN[22]), .ZN(n92) );
  INV_X1 U2720 ( .A(DATAIN[31]), .ZN(n74) );
  INV_X1 U2721 ( .A(DATAIN[9]), .ZN(n118) );
  INV_X1 U2722 ( .A(DATAIN[8]), .ZN(n120) );
  BUF_X2 U2723 ( .A(n126), .Z(n2662) );
  INV_X2 U2724 ( .A(DATAIN[0]), .ZN(n2677) );
  INV_X1 U2725 ( .A(DATAIN[19]), .ZN(n98) );
  INV_X1 U2726 ( .A(DATAIN[16]), .ZN(n104) );
  INV_X1 U2727 ( .A(DATAIN[17]), .ZN(n102) );
  CLKBUF_X1 U2728 ( .A(DATAIN[21]), .Z(n2663) );
  INV_X2 U2729 ( .A(n2663), .ZN(n94) );
  INV_X4 U2730 ( .A(n120), .ZN(n119) );
  INV_X4 U2731 ( .A(n74), .ZN(n73) );
  INV_X4 U2732 ( .A(n98), .ZN(n97) );
  INV_X4 U2733 ( .A(n128), .ZN(n127) );
  INV_X4 U2734 ( .A(n118), .ZN(n117) );
  INV_X4 U2735 ( .A(n130), .ZN(n129) );
  INV_X4 U2736 ( .A(n92), .ZN(n91) );
  CLKBUF_X1 U2737 ( .A(n112), .Z(n2666) );
  INV_X2 U2738 ( .A(DATAIN[12]), .ZN(n112) );
  CLKBUF_X1 U2739 ( .A(n102), .Z(n2667) );
  CLKBUF_X1 U2740 ( .A(n104), .Z(n2668) );
  CLKBUF_X1 U2741 ( .A(n132), .Z(n2669) );
  CLKBUF_X1 U2742 ( .A(n130), .Z(n2670) );
  CLKBUF_X1 U2743 ( .A(n74), .Z(n2671) );
  CLKBUF_X1 U2744 ( .A(n92), .Z(n2672) );
  CLKBUF_X1 U2745 ( .A(n98), .Z(n2673) );
  CLKBUF_X1 U2746 ( .A(n118), .Z(n2674) );
  CLKBUF_X1 U2747 ( .A(n120), .Z(n2675) );
  CLKBUF_X1 U2748 ( .A(n128), .Z(n2676) );
  INV_X2 U2749 ( .A(DATAIN[4]), .ZN(n128) );
  AOI22_X2 U2750 ( .A1(n1532), .A2(n71), .B1(n70), .B2(n2678), .ZN(N407) );
  AOI22_X2 U2751 ( .A1(n798), .A2(n35), .B1(n34), .B2(n2678), .ZN(N275) );
  INV_X2 U2752 ( .A(DATAIN[28]), .ZN(n2678) );
  INV_X2 U2753 ( .A(n110), .ZN(n109) );
  INV_X2 U2754 ( .A(n134), .ZN(n133) );
  INV_X2 U2755 ( .A(n86), .ZN(n85) );
  INV_X2 U2756 ( .A(n96), .ZN(n95) );
  INV_X2 U2757 ( .A(n114), .ZN(n113) );
  INV_X2 U2758 ( .A(n84), .ZN(n83) );
  INV_X2 U2759 ( .A(n132), .ZN(n131) );
  INV_X2 U2760 ( .A(n104), .ZN(n103) );
  INV_X2 U2761 ( .A(n102), .ZN(n101) );
  INV_X2 U2762 ( .A(n112), .ZN(n111) );
  INV_X2 U2763 ( .A(n108), .ZN(n107) );
  INV_X2 U2764 ( .A(n124), .ZN(n123) );
  INV_X2 U2765 ( .A(n82), .ZN(n81) );
endmodule


module SNPS_CLOCK_GATE_HIGH_FFD_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2314, net2316, net2318, net2319, net2322, net2325;
  assign net2314 = EN;
  assign net2316 = CLK;
  assign ENCLK = net2318;
  assign net2325 = TE;

  DLL_X1 latch ( .D(net2319), .GN(net2316), .Q(net2322) );
  OR2_X1 test_or ( .A1(net2314), .A2(net2325), .ZN(net2319) );
  AND2_X1 main_gate ( .A1(net2322), .A2(net2316), .ZN(net2318) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_12 ( CLK, EN, ENCLK, TE
 );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2350, net2352, net2354, net2355, net2358, net2361;
  assign net2350 = EN;
  assign net2352 = CLK;
  assign ENCLK = net2354;
  assign net2361 = TE;

  DLL_X1 latch ( .D(net2355), .GN(net2352), .Q(net2358) );
  OR2_X1 test_or ( .A1(net2350), .A2(net2361), .ZN(net2355) );
  AND2_X2 main_gate ( .A1(net2358), .A2(net2352), .ZN(net2354) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_11 ( CLK, EN, ENCLK, TE
 );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2350, net2352, net2354, net2355, net2358, net2361;
  assign net2350 = EN;
  assign net2352 = CLK;
  assign ENCLK = net2354;
  assign net2361 = TE;

  DLL_X1 latch ( .D(net2355), .GN(net2352), .Q(net2358) );
  AND2_X1 main_gate ( .A1(net2358), .A2(net2352), .ZN(net2354) );
  OR2_X1 test_or ( .A1(net2350), .A2(net2361), .ZN(net2355) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_10 ( CLK, EN, ENCLK, TE
 );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2350, net2352, net2354, net2355, net2358, net2361;
  assign net2350 = EN;
  assign net2352 = CLK;
  assign ENCLK = net2354;
  assign net2361 = TE;

  DLL_X1 latch ( .D(net2355), .GN(net2352), .Q(net2358) );
  AND2_X1 main_gate ( .A1(net2358), .A2(net2352), .ZN(net2354) );
  OR2_X1 test_or ( .A1(net2350), .A2(net2361), .ZN(net2355) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2350, net2352, net2354, net2355, net2358, net2361;
  assign net2350 = EN;
  assign net2352 = CLK;
  assign ENCLK = net2354;
  assign net2361 = TE;

  DLL_X1 latch ( .D(net2355), .GN(net2352), .Q(net2358) );
  OR2_X1 test_or ( .A1(net2350), .A2(net2361), .ZN(net2355) );
  AND2_X1 main_gate ( .A1(net2358), .A2(net2352), .ZN(net2354) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2350, net2352, net2354, net2355, net2358, net2361;
  assign net2350 = EN;
  assign net2352 = CLK;
  assign ENCLK = net2354;
  assign net2361 = TE;

  DLL_X1 latch ( .D(net2355), .GN(net2352), .Q(net2358) );
  OR2_X1 test_or ( .A1(net2350), .A2(net2361), .ZN(net2355) );
  AND2_X1 main_gate ( .A1(net2358), .A2(net2352), .ZN(net2354) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2350, net2352, net2354, net2355, net2358, net2361;
  assign net2350 = EN;
  assign net2352 = CLK;
  assign ENCLK = net2354;
  assign net2361 = TE;

  DLL_X1 latch ( .D(net2355), .GN(net2352), .Q(net2358) );
  OR2_X1 test_or ( .A1(net2350), .A2(net2361), .ZN(net2355) );
  AND2_X1 main_gate ( .A1(net2358), .A2(net2352), .ZN(net2354) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2350, net2352, net2354, net2355, net2358, net2361;
  assign net2350 = EN;
  assign net2352 = CLK;
  assign ENCLK = net2354;
  assign net2361 = TE;

  DLL_X1 latch ( .D(net2355), .GN(net2352), .Q(net2358) );
  OR2_X1 test_or ( .A1(net2350), .A2(net2361), .ZN(net2355) );
  AND2_X1 main_gate ( .A1(net2358), .A2(net2352), .ZN(net2354) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2350, net2352, net2354, net2355, net2358, net2361;
  assign net2350 = EN;
  assign net2352 = CLK;
  assign ENCLK = net2354;
  assign net2361 = TE;

  DLL_X1 latch ( .D(net2355), .GN(net2352), .Q(net2358) );
  OR2_X1 test_or ( .A1(net2350), .A2(net2361), .ZN(net2355) );
  AND2_X1 main_gate ( .A1(net2358), .A2(net2352), .ZN(net2354) );
endmodule


module SNPS_CLOCK_GATE_HIGH_FFD_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2314, net2316, net2318, net2319, net2322, net2325;
  assign net2314 = EN;
  assign net2316 = CLK;
  assign ENCLK = net2318;
  assign net2325 = TE;

  DLL_X1 latch ( .D(net2319), .GN(net2316), .Q(net2322) );
  OR2_X1 test_or ( .A1(net2314), .A2(net2325), .ZN(net2319) );
  AND2_X1 main_gate ( .A1(net2322), .A2(net2316), .ZN(net2318) );
endmodule


module SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net2350, net2352, net2354, net2355, net2358, net2361;
  assign net2350 = EN;
  assign net2352 = CLK;
  assign ENCLK = net2354;
  assign net2361 = TE;

  DLL_X1 latch ( .D(net2355), .GN(net2352), .Q(net2358) );
  OR2_X1 test_or ( .A1(net2350), .A2(net2361), .ZN(net2355) );
  AND2_X1 main_gate ( .A1(net2358), .A2(net2352), .ZN(net2354) );
endmodule


module DLX_WIDTH32 ( CLK, RST, IROM_ADDR, IROM_DATA, DRAM_EN, DRAM_RW, 
        DRAM_ADDR, DRAM_DATA_IN, DRAM_DATA_OUT );
  output [11:0] IROM_ADDR;
  input [31:0] IROM_DATA;
  output [11:0] DRAM_ADDR;
  input [31:0] DRAM_DATA_IN;
  output [31:0] DRAM_DATA_OUT;
  input CLK, RST;
  output DRAM_EN, DRAM_RW;
  wire   w_IF_EN, w_RF_RD1, w_EX_EN, w_MuxA_SEL, w_MuxB_SEL, w_JUMP_EQ,
         w_JUMP_LINK, w_RF_WE_EX, w_SIGN_LD, w_WB_EN, w_RF_WE, \PC/N34 ,
         \PC/N33 , \PC/N32 , \PC/N31 , \PC/N30 , \PC/N29 , \PC/N28 , \PC/N27 ,
         \PC/N26 , \PC/N25 , \PC/N24 , \PC/N23 , \PC/N22 , \PC/N21 , \PC/N20 ,
         \PC/N19 , \PC/N18 , \PC/N17 , \PC/N16 , \PC/N15 , \PC/N14 , \PC/N13 ,
         \PC/N12 , \PC/N11 , \PC/N10 , \PC/N9 , \PC/N8 , \PC/N7 , \PC/N6 ,
         \PC/N5 , \PC/N4 , \PC/N3 , \PC/N2 , \CU/N79 , \CU/N78 , \CU/N77 ,
         \CU/N76 , \CU/N75 , \CU/N74 , \CU/N73 , \CU/N72 , \CU/N71 , \CU/N70 ,
         \CU/N69 , \CU/N68 , \CU/N67 , \CU/N66 , \CU/N65 , \CU/N64 , \CU/N63 ,
         \CU/N62 , \CU/N61 , \CU/N60 , \CU/N59 , \CU/N58 , \CU/N57 , \CU/N56 ,
         \CU/N55 , \CU/N54 , \CU/N53 , \CU/N52 , \CU/N51 , \CU/N50 , \CU/N49 ,
         \CU/N48 , \CU/N47 , \CU/N46 , \CU/N45 , \CU/N44 , \CU/N43 , \CU/N42 ,
         \CU/N41 , \CU/N40 , \CU/N39 , \CU/cw2[2] , \CU/cw2[1] , \CU/cw1[11] ,
         \CU/cw1[10] , \CU/cw1[9] , \CU/cw1[8] , \CU/cw1[7] , \CU/cw1[6] ,
         \CU/cw1[5] , \CU/cw1[4] , \CU/cw1[3] , \CU/cw1[2] , \CU/cw1[1] ,
         \CU/JUMP3 , \CU/JUMP2 , \CU/JUMP1 , \DP/RegLMD_out[31] ,
         \DP/RegLMD_out[30] , \DP/RegLMD_out[29] , \DP/RegLMD_out[28] ,
         \DP/RegLMD_out[27] , \DP/RegLMD_out[26] , \DP/RegLMD_out[25] ,
         \DP/RegLMD_out[24] , \DP/RegLMD_out[23] , \DP/RegLMD_out[22] ,
         \DP/RegLMD_out[21] , \DP/RegLMD_out[20] , \DP/RegLMD_out[19] ,
         \DP/RegLMD_out[18] , \DP/RegLMD_out[17] , \DP/RegLMD_out[16] ,
         \DP/RegLMD_out[15] , \DP/RegLMD_out[14] , \DP/RegLMD_out[13] ,
         \DP/RegLMD_out[12] , \DP/RegLMD_out[11] , \DP/RegLMD_out[10] ,
         \DP/RegLMD_out[9] , \DP/RegLMD_out[8] , \DP/RegLMD_out[7] ,
         \DP/RegLMD_out[6] , \DP/RegLMD_out[5] , \DP/RegLMD_out[4] ,
         \DP/RegLMD_out[3] , \DP/RegLMD_out[2] , \DP/RegLMD_out[1] ,
         \DP/RegLMD_out[0] , \DP/RegALU2_out[31] , \DP/RegALU2_out[30] ,
         \DP/RegALU2_out[29] , \DP/RegALU2_out[28] , \DP/RegALU2_out[27] ,
         \DP/RegALU2_out[26] , \DP/RegALU2_out[25] , \DP/RegALU2_out[24] ,
         \DP/RegALU2_out[23] , \DP/RegALU2_out[22] , \DP/RegALU2_out[21] ,
         \DP/RegALU2_out[20] , \DP/RegALU2_out[19] , \DP/RegALU2_out[18] ,
         \DP/RegALU2_out[17] , \DP/RegALU2_out[16] , \DP/RegALU2_out[15] ,
         \DP/RegALU2_out[14] , \DP/RegALU2_out[13] , \DP/RegALU2_out[12] ,
         \DP/RegALU2_out[11] , \DP/RegALU2_out[10] , \DP/RegALU2_out[9] ,
         \DP/RegALU2_out[8] , \DP/RegALU2_out[7] , \DP/RegALU2_out[6] ,
         \DP/RegALU2_out[5] , \DP/RegALU2_out[4] , \DP/RegALU2_out[3] ,
         \DP/RegALU2_out[2] , \DP/RegALU2_out[1] , \DP/RegALU2_out[0] ,
         \DP/LOAD8[7] , \DP/LOAD8[6] , \DP/LOAD8[5] , \DP/LOAD8[4] ,
         \DP/LOAD8[3] , \DP/LOAD8[2] , \DP/LOAD8[1] , \DP/LOAD8[0] ,
         \DP/LOAD16[15] , \DP/LOAD16[14] , \DP/LOAD16[13] , \DP/LOAD16[12] ,
         \DP/LOAD16[11] , \DP/LOAD16[10] , \DP/LOAD16[9] , \DP/LOAD16[8] ,
         \DP/FwdD , \DP/RD2[0] , \DP/RD2[1] , \DP/RD2[2] , \DP/RegME_out[31] ,
         \DP/RegME_out[30] , \DP/RegME_out[29] , \DP/RegME_out[28] ,
         \DP/RegME_out[27] , \DP/RegME_out[26] , \DP/RegME_out[25] ,
         \DP/RegME_out[24] , \DP/RegME_out[23] , \DP/RegME_out[22] ,
         \DP/RegME_out[21] , \DP/RegME_out[20] , \DP/RegME_out[19] ,
         \DP/RegME_out[18] , \DP/RegME_out[17] , \DP/RegME_out[16] ,
         \DP/RegME_out[15] , \DP/RegME_out[14] , \DP/RegME_out[13] ,
         \DP/RegME_out[12] , \DP/RegME_out[11] , \DP/RegME_out[10] ,
         \DP/RegME_out[9] , \DP/RegME_out[8] , \DP/RegME_out[7] ,
         \DP/RegME_out[6] , \DP/RegME_out[5] , \DP/RegME_out[4] ,
         \DP/RegME_out[3] , \DP/RegME_out[2] , \DP/RegME_out[1] ,
         \DP/RegME_out[0] , \DP/NPC3[31] , \DP/NPC3[30] , \DP/NPC3[29] ,
         \DP/NPC3[28] , \DP/NPC3[27] , \DP/NPC3[26] , \DP/NPC3[25] ,
         \DP/NPC3[24] , \DP/NPC3[23] , \DP/NPC3[22] , \DP/NPC3[21] ,
         \DP/NPC3[20] , \DP/NPC3[19] , \DP/NPC3[18] , \DP/NPC3[17] ,
         \DP/NPC3[16] , \DP/NPC3[15] , \DP/NPC3[14] , \DP/NPC3[13] ,
         \DP/NPC3[12] , \DP/NPC3[11] , \DP/NPC3[10] , \DP/NPC3[9] ,
         \DP/NPC3[8] , \DP/NPC3[7] , \DP/NPC3[6] , \DP/NPC3[5] , \DP/NPC3[4] ,
         \DP/NPC3[3] , \DP/NPC3[2] , \DP/NPC3[1] , \DP/NPC3[0] , \DP/JREG ,
         \DP/JL1 , \DP/RegA1_out[31] , \DP/RegA1_out[30] , \DP/RegA1_out[29] ,
         \DP/RegA1_out[28] , \DP/RegA1_out[27] , \DP/RegA1_out[26] ,
         \DP/RegA1_out[25] , \DP/RegA1_out[24] , \DP/RegA1_out[23] ,
         \DP/RegA1_out[22] , \DP/RegA1_out[21] , \DP/RegA1_out[20] ,
         \DP/RegA1_out[19] , \DP/RegA1_out[18] , \DP/RegA1_out[17] ,
         \DP/RegA1_out[16] , \DP/RegA1_out[15] , \DP/RegA1_out[14] ,
         \DP/RegA1_out[13] , \DP/RegA1_out[12] , \DP/RegA1_out[11] ,
         \DP/RegA1_out[10] , \DP/RegA1_out[9] , \DP/RegA1_out[8] ,
         \DP/RegA1_out[7] , \DP/RegA1_out[6] , \DP/RegA1_out[5] ,
         \DP/RegA1_out[4] , \DP/RegA1_out[3] , \DP/RegA1_out[2] ,
         \DP/RegA1_out[1] , \DP/RegA1_out[0] , \DP/FwdC[1] , \DP/B[15] ,
         \DP/B[14] , \DP/B[13] , \DP/B[12] , \DP/B[11] , \DP/B[10] , \DP/B[9] ,
         \DP/B[8] , \DP/B[7] , \DP/B[6] , \DP/B[5] , \DP/B[4] , \DP/B[3] ,
         \DP/B[2] , \DP/B[1] , \DP/B[0] , \DP/FwdB[1] , \DP/A[31] , \DP/A[30] ,
         \DP/A[29] , \DP/A[28] , \DP/A[27] , \DP/A[26] , \DP/A[25] ,
         \DP/A[24] , \DP/A[15] , \DP/A[14] , \DP/A[13] , \DP/A[12] ,
         \DP/A[11] , \DP/A[10] , \DP/A[9] , \DP/A[8] , \DP/A[7] , \DP/A[6] ,
         \DP/A[5] , \DP/A[4] , \DP/A[3] , \DP/A[2] , \DP/A[1] , \DP/A[0] ,
         \DP/RegALU1_out[12] , \DP/RegALU1_out[13] , \DP/RegALU1_out[14] ,
         \DP/RegALU1_out[15] , \DP/RegALU1_out[16] , \DP/RegALU1_out[17] ,
         \DP/RegALU1_out[18] , \DP/RegALU1_out[19] , \DP/RegALU1_out[20] ,
         \DP/RegALU1_out[21] , \DP/RegALU1_out[22] , \DP/RegALU1_out[23] ,
         \DP/RegALU1_out[24] , \DP/RegALU1_out[25] , \DP/RegALU1_out[26] ,
         \DP/RegALU1_out[27] , \DP/RegALU1_out[28] , \DP/RegALU1_out[29] ,
         \DP/RegALU1_out[30] , \DP/RegALU1_out[31] , \DP/RD1[0] , \DP/RD1[1] ,
         \DP/RD1[2] , \DP/RD1[3] , \DP/RD1[4] , \DP/RegIMM_out[31] ,
         \DP/RegIMM_out[30] , \DP/RegIMM_out[29] , \DP/RegIMM_out[28] ,
         \DP/RegIMM_out[27] , \DP/RegIMM_out[26] , \DP/RegIMM_out[25] ,
         \DP/RegIMM_out[24] , \DP/RegIMM_out[23] , \DP/RegIMM_out[22] ,
         \DP/RegIMM_out[21] , \DP/RegIMM_out[20] , \DP/RegIMM_out[19] ,
         \DP/RegIMM_out[18] , \DP/RegIMM_out[17] , \DP/RegIMM_out[16] ,
         \DP/RegIMM_out[15] , \DP/RegIMM_out[14] , \DP/RegIMM_out[13] ,
         \DP/RegIMM_out[12] , \DP/RegIMM_out[11] , \DP/RegIMM_out[10] ,
         \DP/RegIMM_out[9] , \DP/RegIMM_out[8] , \DP/RegIMM_out[7] ,
         \DP/RegIMM_out[6] , \DP/RegIMM_out[5] , \DP/RegIMM_out[4] ,
         \DP/RegIMM_out[3] , \DP/RegIMM_out[2] , \DP/RegIMM_out[1] ,
         \DP/RegIMM_out[0] , \DP/RegB_out[0] , \DP/RegB_out[1] ,
         \DP/RegB_out[2] , \DP/RegB_out[3] , \DP/RegB_out[4] ,
         \DP/RegB_out[5] , \DP/RegB_out[6] , \DP/RegB_out[7] ,
         \DP/RegB_out[8] , \DP/RegB_out[9] , \DP/RegB_out[10] ,
         \DP/RegB_out[11] , \DP/RegB_out[12] , \DP/RegB_out[13] ,
         \DP/RegB_out[14] , \DP/RegB_out[15] , \DP/RegB_out[16] ,
         \DP/RegB_out[17] , \DP/RegB_out[18] , \DP/RegB_out[19] ,
         \DP/RegB_out[20] , \DP/RegB_out[21] , \DP/RegB_out[22] ,
         \DP/RegB_out[23] , \DP/RegB_out[24] , \DP/RegB_out[25] ,
         \DP/RegB_out[26] , \DP/RegB_out[27] , \DP/RegB_out[28] ,
         \DP/RegB_out[29] , \DP/RegB_out[30] , \DP/RegB_out[31] ,
         \DP/RegA_out[0] , \DP/RegA_out[1] , \DP/RegA_out[2] ,
         \DP/RegA_out[3] , \DP/RegA_out[4] , \DP/RegA_out[5] ,
         \DP/RegA_out[6] , \DP/RegA_out[7] , \DP/RegA_out[8] ,
         \DP/RegA_out[9] , \DP/RegA_out[10] , \DP/RegA_out[11] ,
         \DP/RegA_out[12] , \DP/RegA_out[13] , \DP/RegA_out[14] ,
         \DP/RegA_out[15] , \DP/RegA_out[16] , \DP/RegA_out[17] ,
         \DP/RegA_out[18] , \DP/RegA_out[19] , \DP/RegA_out[20] ,
         \DP/RegA_out[21] , \DP/RegA_out[22] , \DP/RegA_out[23] ,
         \DP/RegA_out[24] , \DP/RegA_out[25] , \DP/RegA_out[26] ,
         \DP/RegA_out[27] , \DP/RegA_out[28] , \DP/RegA_out[29] ,
         \DP/RegA_out[30] , \DP/RegA_out[31] , \DP/NPC2[0] , \DP/NPC2[1] ,
         \DP/NPC2[2] , \DP/NPC2[3] , \DP/NPC2[4] , \DP/NPC2[5] , \DP/NPC2[6] ,
         \DP/NPC2[7] , \DP/NPC2[8] , \DP/NPC2[9] , \DP/NPC2[10] ,
         \DP/NPC2[11] , \DP/NPC2[12] , \DP/NPC2[13] , \DP/NPC2[14] ,
         \DP/NPC2[15] , \DP/NPC2[16] , \DP/NPC2[17] , \DP/NPC2[18] ,
         \DP/NPC2[19] , \DP/NPC2[20] , \DP/NPC2[21] , \DP/NPC2[22] ,
         \DP/NPC2[23] , \DP/NPC2[24] , \DP/NPC2[25] , \DP/NPC2[26] ,
         \DP/NPC2[27] , \DP/NPC2[28] , \DP/NPC2[29] , \DP/NPC2[30] ,
         \DP/NPC2[31] , \DP/RegB_in[31] , \DP/RegB_in[30] , \DP/RegB_in[29] ,
         \DP/RegB_in[28] , \DP/RegB_in[27] , \DP/RegB_in[26] ,
         \DP/RegB_in[25] , \DP/RegB_in[24] , \DP/RegB_in[23] ,
         \DP/RegB_in[22] , \DP/RegB_in[21] , \DP/RegB_in[20] ,
         \DP/RegB_in[19] , \DP/RegB_in[18] , \DP/RegB_in[17] ,
         \DP/RegB_in[16] , \DP/RegB_in[15] , \DP/RegB_in[14] ,
         \DP/RegB_in[13] , \DP/RegB_in[12] , \DP/RegB_in[11] ,
         \DP/RegB_in[10] , \DP/RegB_in[9] , \DP/RegB_in[8] , \DP/RegB_in[7] ,
         \DP/RegB_in[6] , \DP/RegB_in[5] , \DP/RegB_in[4] , \DP/RegB_in[3] ,
         \DP/RegB_in[2] , \DP/RegB_in[1] , \DP/RegB_in[0] , \DP/RegA_in[31] ,
         \DP/RegA_in[30] , \DP/RegA_in[29] , \DP/RegA_in[28] ,
         \DP/RegA_in[27] , \DP/RegA_in[26] , \DP/RegA_in[25] ,
         \DP/RegA_in[24] , \DP/RegA_in[23] , \DP/RegA_in[22] ,
         \DP/RegA_in[21] , \DP/RegA_in[20] , \DP/RegA_in[19] ,
         \DP/RegA_in[18] , \DP/RegA_in[17] , \DP/RegA_in[16] ,
         \DP/RegA_in[15] , \DP/RegA_in[14] , \DP/RegA_in[13] ,
         \DP/RegA_in[12] , \DP/RegA_in[11] , \DP/RegA_in[10] , \DP/RegA_in[9] ,
         \DP/RegA_in[8] , \DP/RegA_in[7] , \DP/RegA_in[6] , \DP/RegA_in[5] ,
         \DP/RegA_in[4] , \DP/RegA_in[3] , \DP/RegA_in[2] , \DP/RegA_in[1] ,
         \DP/RegA_in[0] , \DP/RF_ADDR[4] , \DP/RF_ADDR[3] , \DP/RF_ADDR[2] ,
         \DP/RF_ADDR[1] , \DP/RF_ADDR[0] , \DP/RD3[4] , \DP/RD3[3] ,
         \DP/RD3[2] , \DP/RD3[1] , \DP/RD3[0] , \DP/RF_DATA[31] ,
         \DP/RF_DATA[30] , \DP/RF_DATA[29] , \DP/RF_DATA[28] ,
         \DP/RF_DATA[27] , \DP/RF_DATA[26] , \DP/RF_DATA[25] ,
         \DP/RF_DATA[24] , \DP/RF_DATA[23] , \DP/RF_DATA[22] ,
         \DP/RF_DATA[21] , \DP/RF_DATA[20] , \DP/RF_DATA[19] ,
         \DP/RF_DATA[18] , \DP/RF_DATA[17] , \DP/RF_DATA[16] ,
         \DP/RF_DATA[15] , \DP/RF_DATA[14] , \DP/RF_DATA[13] ,
         \DP/RF_DATA[12] , \DP/RF_DATA[11] , \DP/RF_DATA[10] , \DP/RF_DATA[9] ,
         \DP/RF_DATA[8] , \DP/RF_DATA[7] , \DP/RF_DATA[6] , \DP/RF_DATA[5] ,
         \DP/RF_DATA[4] , \DP/RF_DATA[3] , \DP/RF_DATA[2] , \DP/RF_DATA[1] ,
         \DP/RF_DATA[0] , \DP/JL2 , \DP/NPC_out[31] , \DP/NPC_out[30] ,
         \DP/NPC_out[29] , \DP/NPC_out[28] , \DP/NPC_out[27] ,
         \DP/NPC_out[26] , \DP/NPC_out[25] , \DP/NPC_out[24] ,
         \DP/NPC_out[23] , \DP/NPC_out[22] , \DP/NPC_out[21] ,
         \DP/NPC_out[20] , \DP/NPC_out[19] , \DP/NPC_out[18] ,
         \DP/NPC_out[17] , \DP/NPC_out[16] , \DP/NPC_out[15] ,
         \DP/NPC_out[14] , \DP/NPC_out[13] , \DP/NPC_out[12] ,
         \DP/NPC_out[11] , \DP/NPC_out[10] , \DP/NPC_out[9] , \DP/NPC_out[8] ,
         \DP/NPC_out[7] , \DP/NPC_out[6] , \DP/NPC_out[5] , \DP/NPC_out[4] ,
         \DP/NPC_out[3] , \DP/NPC_out[2] , \DP/NPC_out[1] , \DP/NPC_out[0] ,
         \DP/NPC1[31] , \DP/NPC1[30] , \DP/NPC1[29] , \DP/NPC1[28] ,
         \DP/NPC1[27] , \DP/NPC1[26] , \DP/NPC1[25] , \DP/NPC1[24] ,
         \DP/NPC1[23] , \DP/NPC1[22] , \DP/NPC1[21] , \DP/NPC1[20] ,
         \DP/NPC1[19] , \DP/NPC1[18] , \DP/NPC1[17] , \DP/NPC1[16] ,
         \DP/NPC1[15] , \DP/NPC1[14] , \DP/NPC1[13] , \DP/NPC1[12] ,
         \DP/NPC1[11] , \DP/NPC1[10] , \DP/NPC1[9] , \DP/NPC1[8] ,
         \DP/NPC1[7] , \DP/NPC1[6] , \DP/NPC1[5] , \DP/NPC1[4] , \DP/NPC1[3] ,
         \DP/NPC1[2] , \DP/NPC1[1] , \DP/NPC1[0] , \DP/OUTCOME , \IR/N34 ,
         \IR/N33 , \IR/N32 , \IR/N31 , \IR/N30 , \IR/N29 , \IR/N28 , \IR/N27 ,
         \IR/N26 , \IR/N25 , \IR/N24 , \IR/N23 , \IR/N22 , \IR/N21 , \IR/N20 ,
         \IR/N19 , \IR/N18 , \IR/N17 , \IR/N16 , \IR/N15 , \IR/N14 , \IR/N13 ,
         \IR/N12 , \IR/N11 , \IR/N10 , \IR/N9 , \IR/N8 , \IR/N7 , \IR/N6 ,
         \IR/N5 , \IR/N4 , \IR/N3 , \DP/RegRD1/N7 , \DP/RegRD1/N6 ,
         \DP/RegRD1/N5 , \DP/RegRD1/N4 , \DP/RegRD1/N3 , \DP/ALU0/N91 ,
         \DP/ALU0/N89 , \DP/ALU0/N88 , \DP/ALU0/N85 , \DP/ALU0/N84 ,
         \DP/ALU0/N83 , \DP/ALU0/N82 , \DP/ALU0/N81 , \DP/ALU0/N80 ,
         \DP/ALU0/N79 , \DP/ALU0/N78 , \DP/ALU0/N77 , \DP/ALU0/N76 ,
         \DP/ALU0/N75 , \DP/ALU0/N74 , \DP/ALU0/N73 , \DP/ALU0/N72 ,
         \DP/ALU0/N71 , \DP/ALU0/N70 , \DP/ALU0/N69 , \DP/ALU0/N68 ,
         \DP/ALU0/N67 , \DP/ALU0/N66 , \DP/ALU0/N65 , \DP/ALU0/N64 ,
         \DP/ALU0/N63 , \DP/ALU0/N62 , \DP/ALU0/N61 , \DP/ALU0/N60 ,
         \DP/ALU0/N59 , \DP/ALU0/N58 , \DP/ALU0/N57 , \DP/ALU0/N56 ,
         \DP/ALU0/N55 , \DP/ALU0/N54 , \DP/ALU0/N53 , \DP/ALU0/N52 ,
         \DP/ALU0/N51 , \DP/ALU0/N50 , \DP/ALU0/N49 , \DP/ALU0/N48 ,
         \DP/ALU0/N47 , \DP/ALU0/N46 , \DP/ALU0/N45 , \DP/ALU0/N44 ,
         \DP/ALU0/N43 , \DP/ALU0/N42 , \DP/ALU0/N41 , \DP/ALU0/N40 ,
         \DP/ALU0/N39 , \DP/ALU0/N38 , \DP/ALU0/N37 , \DP/ALU0/N36 ,
         \DP/ALU0/N35 , \DP/ALU0/N34 , \DP/ALU0/N33 , \DP/ALU0/N32 ,
         \DP/ALU0/N31 , \DP/ALU0/N30 , \DP/ALU0/N29 , \DP/ALU0/N28 ,
         \DP/ALU0/N27 , \DP/ALU0/N25 , \DP/ALU0/N23 , \DP/ALU0/N22 ,
         \DP/ALU0/N21 , \DP/ALU0/S_B_LHI[15] , \DP/ALU0/S_B_LHI[14] ,
         \DP/ALU0/S_B_LHI[13] , \DP/ALU0/S_B_LHI[12] , \DP/ALU0/S_B_LHI[11] ,
         \DP/ALU0/S_B_LHI[10] , \DP/ALU0/S_B_LHI[9] , \DP/ALU0/S_B_LHI[8] ,
         \DP/ALU0/S_B_LHI[7] , \DP/ALU0/S_B_LHI[6] , \DP/ALU0/S_B_LHI[5] ,
         \DP/ALU0/S_B_LHI[4] , \DP/ALU0/S_B_LHI[3] , \DP/ALU0/S_B_LHI[2] ,
         \DP/ALU0/S_B_LHI[1] , \DP/ALU0/S_B_LHI[0] , \DP/ALU0/S_B_MULT[5] ,
         \DP/ALU0/S_B_MULT[4] , \DP/ALU0/S_B_MULT[3] , \DP/ALU0/S_B_MULT[2] ,
         \DP/ALU0/S_B_MULT[1] , \DP/ALU0/S_B_MULT[0] , \DP/ALU0/s_A_MULT[13] ,
         \DP/ALU0/s_A_MULT[12] , \DP/ALU0/s_A_MULT[11] ,
         \DP/ALU0/s_A_MULT[10] , \DP/ALU0/s_A_MULT[9] , \DP/ALU0/s_A_MULT[4] ,
         \DP/ALU0/s_A_MULT[3] , \DP/ALU0/s_A_MULT[2] , \DP/ALU0/s_A_MULT[1] ,
         \DP/ALU0/s_SHIFT[1] , \DP/ALU0/s_SHIFT[0] , \DP/ALU0/S_B_SHIFT[4] ,
         \DP/ALU0/S_B_SHIFT[3] , \DP/ALU0/S_B_SHIFT[2] ,
         \DP/ALU0/S_B_SHIFT[1] , \DP/ALU0/S_B_SHIFT[0] ,
         \DP/ALU0/s_A_SHIFT[31] , \DP/ALU0/s_A_SHIFT[30] ,
         \DP/ALU0/s_A_SHIFT[29] , \DP/ALU0/s_A_SHIFT[28] ,
         \DP/ALU0/s_A_SHIFT[27] , \DP/ALU0/s_A_SHIFT[26] ,
         \DP/ALU0/s_A_SHIFT[25] , \DP/ALU0/s_A_SHIFT[24] ,
         \DP/ALU0/s_A_SHIFT[15] , \DP/ALU0/s_A_SHIFT[14] ,
         \DP/ALU0/s_A_SHIFT[13] , \DP/ALU0/s_A_SHIFT[12] ,
         \DP/ALU0/s_A_SHIFT[11] , \DP/ALU0/s_A_SHIFT[10] ,
         \DP/ALU0/s_A_SHIFT[9] , \DP/ALU0/s_A_SHIFT[8] ,
         \DP/ALU0/s_A_SHIFT[7] , \DP/ALU0/s_A_SHIFT[6] ,
         \DP/ALU0/s_A_SHIFT[5] , \DP/ALU0/s_A_SHIFT[4] ,
         \DP/ALU0/s_A_SHIFT[3] , \DP/ALU0/s_A_SHIFT[2] ,
         \DP/ALU0/s_A_SHIFT[1] , \DP/ALU0/s_A_SHIFT[0] , \DP/ALU0/s_LOGIC[3] ,
         \DP/ALU0/s_LOGIC[2] , \DP/ALU0/S_B_LOGIC[15] ,
         \DP/ALU0/S_B_LOGIC[14] , \DP/ALU0/S_B_LOGIC[13] ,
         \DP/ALU0/S_B_LOGIC[12] , \DP/ALU0/S_B_LOGIC[11] ,
         \DP/ALU0/S_B_LOGIC[10] , \DP/ALU0/S_B_LOGIC[9] ,
         \DP/ALU0/S_B_LOGIC[8] , \DP/ALU0/S_B_LOGIC[7] ,
         \DP/ALU0/S_B_LOGIC[6] , \DP/ALU0/S_B_LOGIC[5] ,
         \DP/ALU0/S_B_LOGIC[4] , \DP/ALU0/S_B_LOGIC[3] ,
         \DP/ALU0/S_B_LOGIC[2] , \DP/ALU0/S_B_LOGIC[1] ,
         \DP/ALU0/S_B_LOGIC[0] , \DP/ALU0/s_A_LOGIC[15] ,
         \DP/ALU0/s_A_LOGIC[14] , \DP/ALU0/s_A_LOGIC[13] ,
         \DP/ALU0/s_A_LOGIC[12] , \DP/ALU0/s_A_LOGIC[11] ,
         \DP/ALU0/s_A_LOGIC[10] , \DP/ALU0/s_A_LOGIC[9] ,
         \DP/ALU0/s_A_LOGIC[8] , \DP/ALU0/s_A_LOGIC[7] ,
         \DP/ALU0/s_A_LOGIC[6] , \DP/ALU0/s_A_LOGIC[5] ,
         \DP/ALU0/s_A_LOGIC[4] , \DP/ALU0/s_A_LOGIC[3] ,
         \DP/ALU0/s_A_LOGIC[2] , \DP/ALU0/s_A_LOGIC[1] ,
         \DP/ALU0/s_A_LOGIC[0] , \DP/ALU0/S_B_ADDER[31] ,
         \DP/ALU0/S_B_ADDER[30] , \DP/ALU0/S_B_ADDER[29] ,
         \DP/ALU0/S_B_ADDER[28] , \DP/ALU0/S_B_ADDER[27] ,
         \DP/ALU0/S_B_ADDER[26] , \DP/ALU0/S_B_ADDER[25] ,
         \DP/ALU0/S_B_ADDER[24] , \DP/ALU0/S_B_ADDER[23] ,
         \DP/ALU0/S_B_ADDER[22] , \DP/ALU0/S_B_ADDER[21] ,
         \DP/ALU0/S_B_ADDER[20] , \DP/ALU0/S_B_ADDER[19] ,
         \DP/ALU0/S_B_ADDER[18] , \DP/ALU0/S_B_ADDER[17] ,
         \DP/ALU0/S_B_ADDER[16] , \DP/ALU0/S_B_ADDER[15] ,
         \DP/ALU0/S_B_ADDER[14] , \DP/ALU0/S_B_ADDER[13] ,
         \DP/ALU0/S_B_ADDER[12] , \DP/ALU0/S_B_ADDER[11] ,
         \DP/ALU0/S_B_ADDER[10] , \DP/ALU0/S_B_ADDER[9] ,
         \DP/ALU0/S_B_ADDER[8] , \DP/ALU0/S_B_ADDER[7] ,
         \DP/ALU0/S_B_ADDER[6] , \DP/ALU0/S_B_ADDER[5] ,
         \DP/ALU0/S_B_ADDER[4] , \DP/ALU0/S_B_ADDER[3] ,
         \DP/ALU0/S_B_ADDER[2] , \DP/ALU0/S_B_ADDER[1] ,
         \DP/ALU0/S_B_ADDER[0] , \DP/ALU0/s_A_ADDER[31] ,
         \DP/ALU0/s_A_ADDER[30] , \DP/ALU0/s_A_ADDER[29] ,
         \DP/ALU0/s_A_ADDER[28] , \DP/ALU0/s_A_ADDER[27] ,
         \DP/ALU0/s_A_ADDER[26] , \DP/ALU0/s_A_ADDER[25] ,
         \DP/ALU0/s_A_ADDER[24] , \DP/ALU0/s_A_ADDER[23] ,
         \DP/ALU0/s_A_ADDER[22] , \DP/ALU0/s_A_ADDER[21] ,
         \DP/ALU0/s_A_ADDER[20] , \DP/ALU0/s_A_ADDER[19] ,
         \DP/ALU0/s_A_ADDER[18] , \DP/ALU0/s_A_ADDER[17] ,
         \DP/ALU0/s_A_ADDER[16] , \DP/ALU0/s_A_ADDER[15] ,
         \DP/ALU0/s_A_ADDER[14] , \DP/ALU0/s_A_ADDER[13] ,
         \DP/ALU0/s_A_ADDER[12] , \DP/ALU0/s_A_ADDER[11] ,
         \DP/ALU0/s_A_ADDER[10] , \DP/ALU0/s_A_ADDER[9] ,
         \DP/ALU0/s_A_ADDER[8] , \DP/ALU0/s_A_ADDER[7] ,
         \DP/ALU0/s_A_ADDER[6] , \DP/ALU0/s_A_ADDER[5] ,
         \DP/ALU0/s_A_ADDER[4] , \DP/ALU0/s_A_ADDER[3] ,
         \DP/ALU0/s_A_ADDER[2] , \DP/ALU0/s_A_ADDER[1] ,
         \DP/ALU0/s_A_ADDER[0] , \DP/ALU0/s_SIGN , \DP/FFDBRANCH/net2330 ,
         \DP/FFDBRANCH/N3 , \DP/FFDBRANCH/N2 , \DP/RegNPC/net2366 ,
         \DP/RegNPC1/net2366 , \DP/RegNPC1/N34 , \DP/RegNPC1/N33 ,
         \DP/RegNPC1/N32 , \DP/RegNPC1/N31 , \DP/RegNPC1/N30 ,
         \DP/RegNPC1/N29 , \DP/RegNPC1/N28 , \DP/RegNPC1/N27 ,
         \DP/RegNPC1/N26 , \DP/RegNPC1/N25 , \DP/RegNPC1/N24 ,
         \DP/RegNPC1/N23 , \DP/RegNPC1/N22 , \DP/RegNPC1/N21 ,
         \DP/RegNPC1/N20 , \DP/RegNPC1/N19 , \DP/RegNPC1/N18 ,
         \DP/RegNPC1/N17 , \DP/RegNPC1/N16 , \DP/RegNPC1/N15 ,
         \DP/RegNPC1/N14 , \DP/RegNPC1/N13 , \DP/RegNPC1/N12 ,
         \DP/RegNPC1/N11 , \DP/RegNPC1/N10 , \DP/RegNPC1/N9 , \DP/RegNPC1/N8 ,
         \DP/RegNPC1/N7 , \DP/RegNPC1/N6 , \DP/RegNPC1/N5 , \DP/RegNPC1/N4 ,
         \DP/RegNPC1/N3 , \DP/RegNPC1/N2 , \DP/RegA/net2366 , \DP/RegA/N34 ,
         \DP/RegA/N33 , \DP/RegA/N32 , \DP/RegA/N31 , \DP/RegA/N30 ,
         \DP/RegA/N29 , \DP/RegA/N28 , \DP/RegA/N27 , \DP/RegA/N26 ,
         \DP/RegA/N25 , \DP/RegA/N24 , \DP/RegA/N23 , \DP/RegA/N22 ,
         \DP/RegA/N21 , \DP/RegA/N20 , \DP/RegA/N19 , \DP/RegA/N18 ,
         \DP/RegA/N17 , \DP/RegA/N16 , \DP/RegA/N15 , \DP/RegA/N14 ,
         \DP/RegA/N13 , \DP/RegA/N12 , \DP/RegA/N11 , \DP/RegA/N10 ,
         \DP/RegA/N9 , \DP/RegA/N8 , \DP/RegA/N7 , \DP/RegA/N6 , \DP/RegA/N5 ,
         \DP/RegA/N4 , \DP/RegA/N3 , \DP/RegA/N2 , \DP/RegB/net2366 ,
         \DP/RegB/N34 , \DP/RegB/N33 , \DP/RegB/N32 , \DP/RegB/N31 ,
         \DP/RegB/N30 , \DP/RegB/N29 , \DP/RegB/N28 , \DP/RegB/N27 ,
         \DP/RegB/N26 , \DP/RegB/N25 , \DP/RegB/N24 , \DP/RegB/N23 ,
         \DP/RegB/N22 , \DP/RegB/N21 , \DP/RegB/N20 , \DP/RegB/N19 ,
         \DP/RegB/N18 , \DP/RegB/N17 , \DP/RegB/N16 , \DP/RegB/N15 ,
         \DP/RegB/N14 , \DP/RegB/N13 , \DP/RegB/N12 , \DP/RegB/N11 ,
         \DP/RegB/N10 , \DP/RegB/N9 , \DP/RegB/N8 , \DP/RegB/N7 , \DP/RegB/N6 ,
         \DP/RegB/N5 , \DP/RegB/N4 , \DP/RegB/N3 , \DP/RegB/N2 ,
         \DP/RegIMM/N34 , \DP/RegIMM/N27 , \DP/RegIMM/N26 , \DP/RegIMM/N25 ,
         \DP/RegIMM/N24 , \DP/RegIMM/N23 , \DP/RegIMM/N22 , \DP/RegIMM/N21 ,
         \DP/RegIMM/N20 , \DP/RegIMM/N19 , \DP/RegIMM/N13 , \DP/RegIMM/N12 ,
         \DP/RegIMM/N11 , \DP/RegIMM/N10 , \DP/RegIMM/N9 , \DP/RegIMM/N8 ,
         \DP/RegIMM/N7 , \DP/RegIMM/N6 , \DP/RegIMM/N5 , \DP/RegIMM/N4 ,
         \DP/RegIMM/N3 , \DP/RegA1/net2366 , \DP/RegA1/N34 , \DP/RegA1/N33 ,
         \DP/RegA1/N32 , \DP/RegA1/N31 , \DP/RegA1/N30 , \DP/RegA1/N29 ,
         \DP/RegA1/N28 , \DP/RegA1/N27 , \DP/RegA1/N26 , \DP/RegA1/N25 ,
         \DP/RegA1/N24 , \DP/RegA1/N23 , \DP/RegA1/N22 , \DP/RegA1/N21 ,
         \DP/RegA1/N20 , \DP/RegA1/N19 , \DP/RegA1/N18 , \DP/RegA1/N17 ,
         \DP/RegA1/N16 , \DP/RegA1/N15 , \DP/RegA1/N14 , \DP/RegA1/N13 ,
         \DP/RegA1/N12 , \DP/RegA1/N11 , \DP/RegA1/N10 , \DP/RegA1/N9 ,
         \DP/RegA1/N8 , \DP/RegA1/N7 , \DP/RegA1/N6 , \DP/RegA1/N5 ,
         \DP/RegA1/N4 , \DP/RegA1/N3 , \DP/RegA1/N2 , \DP/FFDJL1/N3 ,
         \DP/FFDJREG/N3 , \DP/RegNPC2/net2366 , \DP/RegNPC2/N34 ,
         \DP/RegNPC2/N33 , \DP/RegNPC2/N32 , \DP/RegNPC2/N31 ,
         \DP/RegNPC2/N30 , \DP/RegNPC2/N29 , \DP/RegNPC2/N28 ,
         \DP/RegNPC2/N27 , \DP/RegNPC2/N26 , \DP/RegNPC2/N25 ,
         \DP/RegNPC2/N24 , \DP/RegNPC2/N23 , \DP/RegNPC2/N22 ,
         \DP/RegNPC2/N21 , \DP/RegNPC2/N20 , \DP/RegNPC2/N19 ,
         \DP/RegNPC2/N18 , \DP/RegNPC2/N17 , \DP/RegNPC2/N16 ,
         \DP/RegNPC2/N15 , \DP/RegNPC2/N14 , \DP/RegNPC2/N13 ,
         \DP/RegNPC2/N12 , \DP/RegNPC2/N11 , \DP/RegNPC2/N10 , \DP/RegNPC2/N9 ,
         \DP/RegNPC2/N8 , \DP/RegNPC2/N7 , \DP/RegNPC2/N6 , \DP/RegNPC2/N5 ,
         \DP/RegNPC2/N4 , \DP/RegNPC2/N3 , \DP/RegNPC2/N2 ,
         \DP/RegALU1/net2366 , \DP/RegALU1/N34 , \DP/RegALU1/N33 ,
         \DP/RegALU1/N32 , \DP/RegALU1/N31 , \DP/RegALU1/N30 ,
         \DP/RegALU1/N29 , \DP/RegALU1/N28 , \DP/RegALU1/N27 ,
         \DP/RegALU1/N26 , \DP/RegALU1/N25 , \DP/RegALU1/N24 ,
         \DP/RegALU1/N23 , \DP/RegALU1/N22 , \DP/RegALU1/N21 ,
         \DP/RegALU1/N20 , \DP/RegALU1/N19 , \DP/RegALU1/N18 ,
         \DP/RegALU1/N17 , \DP/RegALU1/N16 , \DP/RegALU1/N15 ,
         \DP/RegALU1/N14 , \DP/RegALU1/N13 , \DP/RegALU1/N12 ,
         \DP/RegALU1/N11 , \DP/RegALU1/N10 , \DP/RegALU1/N9 , \DP/RegALU1/N8 ,
         \DP/RegALU1/N7 , \DP/RegALU1/N6 , \DP/RegALU1/N5 , \DP/RegALU1/N4 ,
         \DP/RegALU1/N3 , \DP/RegALU1/N2 , \DP/RegME/N34 , \DP/RegME/N33 ,
         \DP/RegME/N32 , \DP/RegME/N31 , \DP/RegME/N30 , \DP/RegME/N29 ,
         \DP/RegME/N28 , \DP/RegME/N27 , \DP/RegME/N26 , \DP/RegME/N25 ,
         \DP/RegME/N24 , \DP/RegME/N23 , \DP/RegME/N22 , \DP/RegME/N21 ,
         \DP/RegME/N20 , \DP/RegME/N19 , \DP/RegME/N18 , \DP/RegME/N17 ,
         \DP/RegME/N16 , \DP/RegME/N15 , \DP/RegME/N14 , \DP/RegME/N13 ,
         \DP/RegME/N12 , \DP/RegME/N11 , \DP/RegME/N10 , \DP/RegME/N9 ,
         \DP/RegME/N8 , \DP/RegME/N7 , \DP/RegME/N6 , \DP/RegME/N5 ,
         \DP/RegME/N4 , \DP/RegME/N3 , \DP/RegRD2/N7 , \DP/RegRD2/N6 ,
         \DP/RegRD2/N5 , \DP/RegRD2/N4 , \DP/RegRD2/N3 , \DP/RegALU2/N34 ,
         \DP/RegALU2/N33 , \DP/RegALU2/N32 , \DP/RegALU2/N31 ,
         \DP/RegALU2/N30 , \DP/RegALU2/N29 , \DP/RegALU2/N28 ,
         \DP/RegALU2/N27 , \DP/RegALU2/N26 , \DP/RegALU2/N25 ,
         \DP/RegALU2/N24 , \DP/RegALU2/N23 , \DP/RegALU2/N22 ,
         \DP/RegALU2/N21 , \DP/RegALU2/N20 , \DP/RegALU2/N19 ,
         \DP/RegALU2/N18 , \DP/RegALU2/N17 , \DP/RegALU2/N16 ,
         \DP/RegALU2/N15 , \DP/RegALU2/N14 , \DP/RegALU2/N13 ,
         \DP/RegALU2/N12 , \DP/RegALU2/N11 , \DP/RegALU2/N10 , \DP/RegALU2/N9 ,
         \DP/RegALU2/N8 , \DP/RegALU2/N7 , \DP/RegALU2/N6 , \DP/RegALU2/N5 ,
         \DP/RegALU2/N4 , \DP/RegALU2/N3 , \DP/RegLMD/net2366 ,
         \DP/RegLMD/N34 , \DP/RegLMD/N33 , \DP/RegLMD/N32 , \DP/RegLMD/N31 ,
         \DP/RegLMD/N30 , \DP/RegLMD/N29 , \DP/RegLMD/N28 , \DP/RegLMD/N27 ,
         \DP/RegLMD/N26 , \DP/RegLMD/N25 , \DP/RegLMD/N24 , \DP/RegLMD/N23 ,
         \DP/RegLMD/N22 , \DP/RegLMD/N21 , \DP/RegLMD/N20 , \DP/RegLMD/N19 ,
         \DP/RegLMD/N18 , \DP/RegLMD/N17 , \DP/RegLMD/N16 , \DP/RegLMD/N15 ,
         \DP/RegLMD/N14 , \DP/RegLMD/N13 , \DP/RegLMD/N12 , \DP/RegLMD/N11 ,
         \DP/RegLMD/N10 , \DP/RegLMD/N9 , \DP/RegLMD/N8 , \DP/RegLMD/N7 ,
         \DP/RegLMD/N6 , \DP/RegLMD/N5 , \DP/RegLMD/N4 , \DP/RegLMD/N3 ,
         \DP/RegRD3/N7 , \DP/RegRD3/N6 , \DP/RegRD3/N5 , \DP/RegRD3/N4 ,
         \DP/RegRD3/N3 , \DP/FFDJL2/net2330 , \DP/FFDJL2/N3 , \DP/FFDJL2/N2 ,
         \DP/RegNPC3/net2366 , \DP/RegNPC3/N34 , \DP/RegNPC3/N33 ,
         \DP/RegNPC3/N32 , \DP/RegNPC3/N31 , \DP/RegNPC3/N30 ,
         \DP/RegNPC3/N29 , \DP/RegNPC3/N28 , \DP/RegNPC3/N27 ,
         \DP/RegNPC3/N26 , \DP/RegNPC3/N25 , \DP/RegNPC3/N24 ,
         \DP/RegNPC3/N23 , \DP/RegNPC3/N22 , \DP/RegNPC3/N21 ,
         \DP/RegNPC3/N20 , \DP/RegNPC3/N19 , \DP/RegNPC3/N18 ,
         \DP/RegNPC3/N17 , \DP/RegNPC3/N16 , \DP/RegNPC3/N15 ,
         \DP/RegNPC3/N14 , \DP/RegNPC3/N13 , \DP/RegNPC3/N12 ,
         \DP/RegNPC3/N11 , \DP/RegNPC3/N10 , \DP/RegNPC3/N9 , \DP/RegNPC3/N8 ,
         \DP/RegNPC3/N7 , \DP/RegNPC3/N6 , \DP/RegNPC3/N5 , \DP/RegNPC3/N4 ,
         \DP/RegNPC3/N3 , \DP/RegNPC3/N2 , \DP/RegFB/N5 , \DP/RegFB/N4 ,
         \DP/RegFB/N3 , \DP/RegFC/N5 , \DP/RegFC/N4 , \DP/RegFC/N3 ,
         \DP/FFDFD/N3 , \DP/ALU0/MULT/SHIFTERi_0/N19 , n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n66, n94, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n109, n110, n112,
         n113, n115, n116, n118, n119, n121, n122, n124, n125, n127, n128,
         n130, n131, n133, n134, n136, n137, n139, n140, n142, n143, n145,
         n146, n148, n149, n151, n152, n154, n155, n157, n158, n161, n164,
         n167, n170, n173, n175, n176, n178, n179, n182, n183, n186, n189,
         n196, n200, n202, n204, n205, n206, n207, n208, n218, n224, n400,
         n401, n404, n405, n406, n407, n575, n578, n580, n582, n584, n1110,
         n1272, n2339, n2340, n2341, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2469, n2470, n2471,
         n2473, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3582, n3583, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3615,
         n3616, n3618, n3620, n3621, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4242, n4243, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4254, n4255, n4256, n4257, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4351, n4352, n4353, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4373, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4424, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4468, n4469, n4470, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918;
  wire   [31:12] w_PC_OUT;
  wire   [31:0] IR_OUT;
  wire   [4:0] w_ALU_OPCODE;
  wire   [2:0] w_LOAD_SIZE;
  assign \DP/LOAD8[7]  = DRAM_DATA_IN[7];
  assign \DP/LOAD8[6]  = DRAM_DATA_IN[6];
  assign \DP/LOAD8[5]  = DRAM_DATA_IN[5];
  assign \DP/LOAD8[4]  = DRAM_DATA_IN[4];
  assign \DP/LOAD8[3]  = DRAM_DATA_IN[3];
  assign \DP/LOAD8[2]  = DRAM_DATA_IN[2];
  assign \DP/LOAD8[1]  = DRAM_DATA_IN[1];
  assign \DP/LOAD8[0]  = DRAM_DATA_IN[0];
  assign \DP/LOAD16[15]  = DRAM_DATA_IN[15];
  assign \DP/LOAD16[14]  = DRAM_DATA_IN[14];
  assign \DP/LOAD16[13]  = DRAM_DATA_IN[13];
  assign \DP/LOAD16[12]  = DRAM_DATA_IN[12];
  assign \DP/LOAD16[11]  = DRAM_DATA_IN[11];
  assign \DP/LOAD16[10]  = DRAM_DATA_IN[10];
  assign \DP/LOAD16[9]  = DRAM_DATA_IN[9];
  assign \DP/LOAD16[8]  = DRAM_DATA_IN[8];

  DFF_X1 \CU/IF_EN_reg  ( .D(n2460), .CK(CLK), .QN(w_IF_EN) );
  DFF_X1 \IR/DOUT_reg[0]  ( .D(\IR/N3 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[0]), .QN(n2375) );
  DFF_X1 \IR/DOUT_reg[1]  ( .D(\IR/N4 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[1]), .QN(n2382) );
  DFF_X1 \IR/DOUT_reg[2]  ( .D(\IR/N5 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[2]), .QN(n2377) );
  DFF_X1 \IR/DOUT_reg[3]  ( .D(\IR/N6 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[3]), .QN(n2390) );
  DFF_X1 \IR/DOUT_reg[4]  ( .D(\IR/N7 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[4]) );
  DFF_X1 \IR/DOUT_reg[5]  ( .D(\IR/N8 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[5]), .QN(n2364) );
  DFF_X1 \IR/DOUT_reg[6]  ( .D(\IR/N9 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[6]) );
  DFF_X1 \IR/DOUT_reg[7]  ( .D(\IR/N10 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[7]) );
  DFF_X1 \IR/DOUT_reg[8]  ( .D(\IR/N11 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[8]) );
  DFF_X1 \IR/DOUT_reg[9]  ( .D(\IR/N12 ), .CK(n2456), .QN(n2391) );
  DFF_X1 \IR/DOUT_reg[10]  ( .D(\IR/N13 ), .CK(n2456), .Q(IR_OUT[10]) );
  DFF_X1 \IR/DOUT_reg[11]  ( .D(\IR/N14 ), .CK(n2456), .Q(IR_OUT[11]) );
  DFF_X1 \IR/DOUT_reg[12]  ( .D(\IR/N15 ), .CK(n2456), .Q(IR_OUT[12]) );
  DFF_X1 \IR/DOUT_reg[13]  ( .D(\IR/N16 ), .CK(n2456), .Q(IR_OUT[13]) );
  DFF_X1 \IR/DOUT_reg[14]  ( .D(\IR/N17 ), .CK(n2456), .Q(IR_OUT[14]) );
  DFF_X1 \IR/DOUT_reg[15]  ( .D(\IR/N18 ), .CK(n2456), .Q(IR_OUT[15]) );
  DFF_X1 \IR/DOUT_reg[16]  ( .D(\IR/N19 ), .CK(n2456), .Q(IR_OUT[16]) );
  DFF_X1 \IR/DOUT_reg[17]  ( .D(\IR/N20 ), .CK(n2456), .Q(IR_OUT[17]) );
  DFF_X1 \IR/DOUT_reg[18]  ( .D(\IR/N21 ), .CK(n2456), .Q(IR_OUT[18]) );
  DFF_X1 \IR/DOUT_reg[19]  ( .D(\IR/N22 ), .CK(n2456), .Q(IR_OUT[19]) );
  DFF_X1 \IR/DOUT_reg[20]  ( .D(\IR/N23 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[20]) );
  DFF_X1 \IR/DOUT_reg[21]  ( .D(\IR/N24 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[21]) );
  DFF_X1 \IR/DOUT_reg[22]  ( .D(\IR/N25 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[22]) );
  DFF_X1 \IR/DOUT_reg[23]  ( .D(\IR/N26 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[23]) );
  DFF_X1 \IR/DOUT_reg[24]  ( .D(\IR/N27 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[24]) );
  DFF_X1 \IR/DOUT_reg[25]  ( .D(\IR/N28 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[25]) );
  DFF_X1 \IR/DOUT_reg[26]  ( .D(\IR/N29 ), .CK(\DP/RegNPC/net2366 ), .Q(n2372), 
        .QN(n224) );
  DFF_X1 \IR/DOUT_reg[27]  ( .D(\IR/N30 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[27]), .QN(n2388) );
  DFF_X1 \IR/DOUT_reg[28]  ( .D(\IR/N31 ), .CK(\DP/RegNPC/net2366 ), .QN(n2394) );
  DFF_X1 \IR/DOUT_reg[29]  ( .D(\IR/N32 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[29]) );
  DFF_X1 \IR/DOUT_reg[30]  ( .D(\IR/N33 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[30]), .QN(n2371) );
  DFF_X1 \IR/DOUT_reg[31]  ( .D(\IR/N34 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IR_OUT[31]), .QN(n2397) );
  DFF_X1 \CU/JUMP1_reg  ( .D(\CU/N72 ), .CK(CLK), .Q(\CU/JUMP1 ), .QN(n4536)
         );
  DFF_X1 \CU/JUMP2_reg  ( .D(\CU/N73 ), .CK(CLK), .Q(\CU/JUMP2 ), .QN(n4537)
         );
  DFF_X1 \CU/JUMP3_reg  ( .D(\CU/N74 ), .CK(CLK), .Q(\CU/JUMP3 ), .QN(n4538)
         );
  DFF_X1 \CU/cw1_reg[13]  ( .D(\CU/N51 ), .CK(CLK), .QN(n207) );
  DFF_X1 \CU/cw1_reg[14]  ( .D(\CU/N52 ), .CK(CLK), .Q(w_JUMP_EQ) );
  DFF_X1 \CU/cw1_reg[6]  ( .D(\CU/N44 ), .CK(CLK), .Q(\CU/cw1[6] ) );
  DFF_X1 \CU/cw2_reg[6]  ( .D(\CU/N63 ), .CK(CLK), .Q(w_SIGN_LD) );
  DFF_X1 \CU/cw1_reg[3]  ( .D(\CU/N41 ), .CK(CLK), .Q(\CU/cw1[3] ) );
  DFF_X1 \CU/cw1_reg[5]  ( .D(\CU/N43 ), .CK(CLK), .Q(\CU/cw1[5] ) );
  DFF_X1 \CU/cw2_reg[5]  ( .D(\CU/N62 ), .CK(CLK), .Q(w_LOAD_SIZE[2]) );
  DFF_X1 \CU/cw1_reg[4]  ( .D(\CU/N42 ), .CK(CLK), .Q(\CU/cw1[4] ) );
  DFF_X1 \CU/cw1_reg[1]  ( .D(\CU/N39 ), .CK(CLK), .Q(\CU/cw1[1] ) );
  DFF_X1 \CU/cw2_reg[1]  ( .D(\CU/N58 ), .CK(CLK), .Q(\CU/cw2[1] ) );
  DFF_X1 \CU/cw1_reg[15]  ( .D(\CU/N53 ), .CK(CLK), .QN(n208) );
  DFF_X1 \CU/aluOpcode1_reg[2]  ( .D(\CU/N77 ), .CK(CLK), .Q(w_ALU_OPCODE[2]), 
        .QN(n2362) );
  DFF_X1 \CU/aluOpcode1_reg[3]  ( .D(\CU/N78 ), .CK(CLK), .Q(w_ALU_OPCODE[3]), 
        .QN(n2374) );
  DFF_X1 \CU/cw1_reg[2]  ( .D(\CU/N40 ), .CK(CLK), .Q(\CU/cw1[2] ) );
  DFF_X1 \CU/cw2_reg[2]  ( .D(\CU/N59 ), .CK(CLK), .Q(\CU/cw2[2] ) );
  DFF_X1 \CU/cw3_reg[2]  ( .D(\CU/N71 ), .CK(CLK), .Q(w_WB_EN) );
  DFF_X1 \CU/cw1_reg[0]  ( .D(\CU/N40 ), .CK(CLK), .Q(w_RF_WE_EX) );
  DFF_X1 \CU/cw2_reg[0]  ( .D(\CU/N57 ), .CK(CLK), .QN(n2395) );
  DFF_X1 \CU/cw3_reg[0]  ( .D(\CU/N69 ), .CK(CLK), .Q(w_RF_WE) );
  DFF_X1 \CU/aluOpcode1_reg[0]  ( .D(\CU/N75 ), .CK(CLK), .Q(n2363), .QN(n218)
         );
  DFF_X1 \CU/cw1_reg[18]  ( .D(\CU/N56 ), .CK(CLK), .Q(w_EX_EN) );
  DFF_X1 \CU/cw1_reg[11]  ( .D(\CU/N49 ), .CK(CLK), .Q(\CU/cw1[11] ) );
  DFF_X1 \CU/cw2_reg[11]  ( .D(\CU/N68 ), .CK(CLK), .Q(DRAM_EN) );
  DFF_X1 \CU/cw1_reg[9]  ( .D(\CU/N47 ), .CK(CLK), .Q(\CU/cw1[9] ) );
  DFF_X1 \CU/cw1_reg[8]  ( .D(\CU/N46 ), .CK(CLK), .Q(\CU/cw1[8] ) );
  DFF_X1 \CU/cw1_reg[7]  ( .D(\CU/N45 ), .CK(CLK), .Q(\CU/cw1[7] ) );
  DFF_X1 \CU/cw2_reg[7]  ( .D(\CU/N64 ), .CK(CLK), .QN(n204) );
  DFF_X1 \CU/cw1_reg[10]  ( .D(\CU/N48 ), .CK(CLK), .Q(\CU/cw1[10] ) );
  DFF_X1 \CU/cw2_reg[10]  ( .D(\CU/N67 ), .CK(CLK), .Q(DRAM_RW) );
  DFF_X1 \DP/RegRD1/DOUT_reg[0]  ( .D(\DP/RegRD1/N3 ), .CK(n2452), .Q(
        \DP/RD1[0] ) );
  DFF_X1 \DP/RegRD1/DOUT_reg[4]  ( .D(\DP/RegRD1/N7 ), .CK(n2452), .Q(
        \DP/RD1[4] ) );
  DLL_X1 \DP/ALU0/s_SHIFT_reg[0]  ( .D(n2339), .GN(n2444), .Q(
        \DP/ALU0/s_SHIFT[0] ) );
  DLL_X1 \DP/ALU0/s_SHIFT_reg[1]  ( .D(n2341), .GN(n2444), .Q(
        \DP/ALU0/s_SHIFT[1] ) );
  DLL_X1 \DP/ALU0/s_LOGIC_reg[2]  ( .D(\DP/ALU0/N88 ), .GN(n2447), .Q(
        \DP/ALU0/s_LOGIC[2] ) );
  DLL_X1 \DP/ALU0/s_LOGIC_reg[3]  ( .D(\DP/ALU0/N89 ), .GN(n2447), .Q(
        \DP/ALU0/s_LOGIC[3] ) );
  DLH_X1 \DP/ALU0/s_ADD_SUB_reg  ( .G(\DP/ALU0/N21 ), .D(n1272), .Q(n57) );
  DFF_X1 \DP/RegIMM/DOUT_reg[0]  ( .D(\DP/RegIMM/N3 ), .CK(n2453), .Q(
        \DP/RegIMM_out[0] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[1]  ( .D(\DP/RegIMM/N4 ), .CK(n2452), .Q(
        \DP/RegIMM_out[1] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[2]  ( .D(\DP/RegIMM/N5 ), .CK(n2452), .Q(
        \DP/RegIMM_out[2] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[3]  ( .D(\DP/RegIMM/N6 ), .CK(n2453), .Q(
        \DP/RegIMM_out[3] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[4]  ( .D(\DP/RegIMM/N7 ), .CK(n2453), .Q(
        \DP/RegIMM_out[4] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[5]  ( .D(\DP/RegIMM/N8 ), .CK(n2453), .Q(
        \DP/RegIMM_out[5] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[6]  ( .D(\DP/RegIMM/N9 ), .CK(n2453), .Q(
        \DP/RegIMM_out[6] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[7]  ( .D(\DP/RegIMM/N10 ), .CK(n2453), .Q(
        \DP/RegIMM_out[7] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[8]  ( .D(\DP/RegIMM/N11 ), .CK(n2453), .Q(
        \DP/RegIMM_out[8] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[9]  ( .D(\DP/RegIMM/N12 ), .CK(n2453), .Q(
        \DP/RegIMM_out[9] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[10]  ( .D(\DP/RegIMM/N13 ), .CK(n2453), .Q(
        \DP/RegIMM_out[10] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[11]  ( .D(n584), .CK(n2453), .QN(
        \DP/RegIMM_out[11] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[12]  ( .D(n582), .CK(n2453), .QN(
        \DP/RegIMM_out[12] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[13]  ( .D(n580), .CK(n2453), .QN(
        \DP/RegIMM_out[13] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[14]  ( .D(n578), .CK(n2455), .QN(
        \DP/RegIMM_out[14] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[15]  ( .D(n575), .CK(n2454), .QN(
        \DP/RegIMM_out[15] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[16]  ( .D(\DP/RegIMM/N19 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegIMM_out[16] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[17]  ( .D(\DP/RegIMM/N20 ), .CK(n2452), .Q(
        \DP/RegIMM_out[17] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[18]  ( .D(\DP/RegIMM/N21 ), .CK(n2454), .Q(
        \DP/RegIMM_out[18] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[19]  ( .D(\DP/RegIMM/N22 ), .CK(n2453), .Q(
        \DP/RegIMM_out[19] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[20]  ( .D(\DP/RegIMM/N23 ), .CK(n2454), .Q(
        \DP/RegIMM_out[20] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[21]  ( .D(\DP/RegIMM/N24 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegIMM_out[21] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[22]  ( .D(\DP/RegIMM/N25 ), .CK(n2453), .Q(
        \DP/RegIMM_out[22] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[23]  ( .D(\DP/RegIMM/N26 ), .CK(n2452), .Q(
        \DP/RegIMM_out[23] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[24]  ( .D(\DP/RegIMM/N27 ), .CK(n2455), .Q(
        \DP/RegIMM_out[24] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[25]  ( .D(\DP/RegIMM/N34 ), .CK(n2452), .Q(
        \DP/RegIMM_out[25] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[26]  ( .D(\DP/RegIMM/N34 ), .CK(n2455), .Q(
        \DP/RegIMM_out[26] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[27]  ( .D(\DP/RegIMM/N34 ), .CK(n2454), .Q(
        \DP/RegIMM_out[27] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[28]  ( .D(\DP/RegIMM/N34 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegIMM_out[28] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[29]  ( .D(\DP/RegIMM/N34 ), .CK(n2453), .Q(
        \DP/RegIMM_out[29] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[30]  ( .D(\DP/RegIMM/N34 ), .CK(n2453), .Q(
        \DP/RegIMM_out[30] ) );
  DFF_X1 \DP/RegIMM/DOUT_reg[31]  ( .D(\DP/RegIMM/N34 ), .CK(n2455), .Q(
        \DP/RegIMM_out[31] ) );
  DFF_X1 \DP/FFDJL1/Q_reg  ( .D(\DP/FFDJL1/N3 ), .CK(\DP/FFDJL2/net2330 ), .Q(
        \DP/JL1 ) );
  DFF_X1 \DP/FFDJREG/Q_reg  ( .D(\DP/FFDJREG/N3 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/JREG ) );
  DFF_X1 \DP/RegRD2/DOUT_reg[0]  ( .D(\DP/RegRD2/N3 ), .CK(n2452), .Q(
        \DP/RD2[0] ) );
  DFF_X1 \DP/RegRD2/DOUT_reg[1]  ( .D(\DP/RegRD2/N4 ), .CK(n2452), .Q(
        \DP/RD2[1] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[0]  ( .D(\DP/RegLMD/N3 ), .CK(\DP/RegLMD/net2366 ), .Q(\DP/RegLMD_out[0] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[1]  ( .D(\DP/RegLMD/N4 ), .CK(\DP/RegLMD/net2366 ), .Q(\DP/RegLMD_out[1] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[2]  ( .D(\DP/RegLMD/N5 ), .CK(\DP/RegLMD/net2366 ), .Q(\DP/RegLMD_out[2] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[3]  ( .D(\DP/RegLMD/N6 ), .CK(\DP/RegLMD/net2366 ), .Q(\DP/RegLMD_out[3] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[4]  ( .D(\DP/RegLMD/N7 ), .CK(\DP/RegLMD/net2366 ), .Q(\DP/RegLMD_out[4] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[5]  ( .D(\DP/RegLMD/N8 ), .CK(\DP/RegLMD/net2366 ), .Q(\DP/RegLMD_out[5] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[6]  ( .D(\DP/RegLMD/N9 ), .CK(\DP/RegLMD/net2366 ), .Q(\DP/RegLMD_out[6] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[7]  ( .D(\DP/RegLMD/N10 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegLMD_out[7] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[8]  ( .D(\DP/RegLMD/N11 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegLMD_out[8] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[9]  ( .D(\DP/RegLMD/N12 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegLMD_out[9] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[10]  ( .D(\DP/RegLMD/N13 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegLMD_out[10] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[11]  ( .D(\DP/RegLMD/N14 ), .CK(n2455), .Q(
        \DP/RegLMD_out[11] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[12]  ( .D(\DP/RegLMD/N15 ), .CK(n2455), .Q(
        \DP/RegLMD_out[12] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[13]  ( .D(\DP/RegLMD/N16 ), .CK(n2455), .Q(
        \DP/RegLMD_out[13] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[14]  ( .D(\DP/RegLMD/N17 ), .CK(n2455), .Q(
        \DP/RegLMD_out[14] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[15]  ( .D(\DP/RegLMD/N18 ), .CK(n2455), .Q(
        \DP/RegLMD_out[15] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[16]  ( .D(\DP/RegLMD/N19 ), .CK(n2455), .Q(
        \DP/RegLMD_out[16] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[17]  ( .D(\DP/RegLMD/N20 ), .CK(n2455), .Q(
        \DP/RegLMD_out[17] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[18]  ( .D(\DP/RegLMD/N21 ), .CK(n2455), .Q(
        \DP/RegLMD_out[18] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[19]  ( .D(\DP/RegLMD/N22 ), .CK(n2455), .Q(
        \DP/RegLMD_out[19] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[20]  ( .D(\DP/RegLMD/N23 ), .CK(n2455), .Q(
        \DP/RegLMD_out[20] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[21]  ( .D(\DP/RegLMD/N24 ), .CK(n2455), .Q(
        \DP/RegLMD_out[21] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[22]  ( .D(\DP/RegLMD/N25 ), .CK(n2454), .Q(
        \DP/RegLMD_out[22] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[23]  ( .D(\DP/RegLMD/N26 ), .CK(n2454), .Q(
        \DP/RegLMD_out[23] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[24]  ( .D(\DP/RegLMD/N27 ), .CK(n2454), .Q(
        \DP/RegLMD_out[24] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[25]  ( .D(\DP/RegLMD/N28 ), .CK(n2454), .Q(
        \DP/RegLMD_out[25] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[26]  ( .D(\DP/RegLMD/N29 ), .CK(n2454), .Q(
        \DP/RegLMD_out[26] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[27]  ( .D(\DP/RegLMD/N30 ), .CK(n2454), .Q(
        \DP/RegLMD_out[27] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[28]  ( .D(\DP/RegLMD/N31 ), .CK(n2454), .Q(
        \DP/RegLMD_out[28] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[29]  ( .D(\DP/RegLMD/N32 ), .CK(n2454), .Q(
        \DP/RegLMD_out[29] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[30]  ( .D(\DP/RegLMD/N33 ), .CK(n2454), .Q(
        \DP/RegLMD_out[30] ) );
  DFF_X1 \DP/RegLMD/DOUT_reg[31]  ( .D(\DP/RegLMD/N34 ), .CK(n2454), .Q(
        \DP/RegLMD_out[31] ) );
  DFF_X1 \DP/RegRD3/DOUT_reg[0]  ( .D(\DP/RegRD3/N3 ), .CK(n2452), .Q(
        \DP/RD3[0] ) );
  DFF_X1 \DP/RegRD3/DOUT_reg[1]  ( .D(\DP/RegRD3/N4 ), .CK(n2454), .Q(
        \DP/RD3[1] ) );
  DFF_X1 \DP/RegRD3/DOUT_reg[2]  ( .D(\DP/RegRD3/N5 ), .CK(n2453), .Q(
        \DP/RD3[2] ) );
  DFF_X1 \DP/RegRD3/DOUT_reg[3]  ( .D(\DP/RegRD3/N6 ), .CK(n2452), .Q(
        \DP/RD3[3] ) );
  DFF_X1 \DP/RegRD3/DOUT_reg[4]  ( .D(\DP/RegRD3/N7 ), .CK(n2452), .Q(
        \DP/RD3[4] ) );
  DFF_X1 \DP/RegFB/DOUT_reg[0]  ( .D(\DP/RegFB/N3 ), .CK(\DP/RegNPC1/net2366 ), 
        .Q(n2368), .QN(n404) );
  DFF_X1 \DP/RegFB/DOUT_reg[1]  ( .D(\DP/RegFB/N4 ), .CK(\DP/RegNPC1/net2366 ), 
        .Q(\DP/FwdB[1] ), .QN(n2404) );
  DFF_X1 \DP/RegA1/DOUT_reg[18]  ( .D(\DP/RegA1/N21 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[18] ) );
  DFF_X1 \DP/FFDBRANCH/Q_reg  ( .D(\DP/FFDBRANCH/N3 ), .CK(
        \DP/FFDBRANCH/net2330 ), .Q(\DP/OUTCOME ), .QN(n2405) );
  DFF_X1 \PC/DOUT_reg[6]  ( .D(\PC/N9 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IROM_ADDR[6]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[6]  ( .D(\PC/N9 ), .CK(\DP/RegNPC/net2366 ), .Q(
        \DP/NPC1[6] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[6]  ( .D(\DP/RegNPC1/N9 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[6] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[6]  ( .D(\DP/RegNPC2/N9 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[6] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[6]  ( .D(\DP/RegNPC3/N9 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[6] ) );
  DFF_X1 \DP/RegB/DOUT_reg[0]  ( .D(\DP/RegB/N3 ), .CK(\DP/RegB/net2366 ), .Q(
        \DP/RegB_out[0] ) );
  DFF_X1 \DP/RegME/DOUT_reg[0]  ( .D(\DP/RegME/N3 ), .CK(n2452), .Q(
        \DP/RegME_out[0] ) );
  DFF_X1 \DP/RegB/DOUT_reg[1]  ( .D(\DP/RegB/N4 ), .CK(\DP/RegB/net2366 ), .Q(
        \DP/RegB_out[1] ) );
  DFF_X1 \DP/RegME/DOUT_reg[1]  ( .D(\DP/RegME/N4 ), .CK(n2453), .Q(
        \DP/RegME_out[1] ) );
  DFF_X1 \DP/RegB/DOUT_reg[2]  ( .D(\DP/RegB/N5 ), .CK(\DP/RegB/net2366 ), .Q(
        \DP/RegB_out[2] ) );
  DFF_X1 \DP/RegME/DOUT_reg[2]  ( .D(\DP/RegME/N5 ), .CK(n2454), .Q(
        \DP/RegME_out[2] ) );
  DFF_X1 \DP/RegB/DOUT_reg[3]  ( .D(\DP/RegB/N6 ), .CK(\DP/RegB/net2366 ), .Q(
        \DP/RegB_out[3] ) );
  DFF_X1 \DP/RegME/DOUT_reg[3]  ( .D(\DP/RegME/N6 ), .CK(n2452), .Q(
        \DP/RegME_out[3] ) );
  DFF_X1 \DP/RegB/DOUT_reg[4]  ( .D(\DP/RegB/N7 ), .CK(\DP/RegB/net2366 ), .Q(
        \DP/RegB_out[4] ) );
  DFF_X1 \DP/RegME/DOUT_reg[4]  ( .D(\DP/RegME/N7 ), .CK(n2453), .Q(
        \DP/RegME_out[4] ) );
  DFF_X1 \DP/RegB/DOUT_reg[5]  ( .D(\DP/RegB/N8 ), .CK(\DP/RegB/net2366 ), .Q(
        \DP/RegB_out[5] ) );
  DFF_X1 \DP/RegME/DOUT_reg[5]  ( .D(\DP/RegME/N8 ), .CK(n2455), .Q(
        \DP/RegME_out[5] ) );
  DFF_X1 \DP/RegB/DOUT_reg[6]  ( .D(\DP/RegB/N9 ), .CK(\DP/RegB/net2366 ), .Q(
        \DP/RegB_out[6] ) );
  DFF_X1 \DP/RegME/DOUT_reg[6]  ( .D(\DP/RegME/N9 ), .CK(n2454), .Q(
        \DP/RegME_out[6] ) );
  DFF_X1 \DP/RegB/DOUT_reg[7]  ( .D(\DP/RegB/N10 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[7] ) );
  DFF_X1 \DP/RegME/DOUT_reg[7]  ( .D(\DP/RegME/N10 ), .CK(n2452), .Q(
        \DP/RegME_out[7] ) );
  DFF_X1 \DP/RegB/DOUT_reg[8]  ( .D(\DP/RegB/N11 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[8] ) );
  DFF_X1 \DP/RegME/DOUT_reg[8]  ( .D(\DP/RegME/N11 ), .CK(n2453), .Q(
        \DP/RegME_out[8] ) );
  DFF_X1 \DP/RegB/DOUT_reg[9]  ( .D(\DP/RegB/N12 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[9] ) );
  DFF_X1 \DP/RegME/DOUT_reg[9]  ( .D(\DP/RegME/N12 ), .CK(n2455), .Q(
        \DP/RegME_out[9] ) );
  DFF_X1 \DP/RegB/DOUT_reg[10]  ( .D(\DP/RegB/N13 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[10] ) );
  DFF_X1 \DP/RegME/DOUT_reg[10]  ( .D(\DP/RegME/N13 ), .CK(n2454), .Q(
        \DP/RegME_out[10] ) );
  DFF_X1 \DP/RegB/DOUT_reg[11]  ( .D(\DP/RegB/N14 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[11] ) );
  DFF_X1 \DP/RegME/DOUT_reg[11]  ( .D(\DP/RegME/N14 ), .CK(n2452), .Q(
        \DP/RegME_out[11] ) );
  DFF_X1 \DP/RegB/DOUT_reg[12]  ( .D(\DP/RegB/N15 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[12] ) );
  DFF_X1 \DP/RegME/DOUT_reg[12]  ( .D(\DP/RegME/N15 ), .CK(n2453), .Q(
        \DP/RegME_out[12] ) );
  DFF_X1 \DP/RegB/DOUT_reg[13]  ( .D(\DP/RegB/N16 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[13] ) );
  DFF_X1 \DP/RegME/DOUT_reg[13]  ( .D(\DP/RegME/N16 ), .CK(n2455), .Q(
        \DP/RegME_out[13] ) );
  DFF_X1 \DP/RegB/DOUT_reg[14]  ( .D(\DP/RegB/N17 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[14] ) );
  DFF_X1 \DP/RegME/DOUT_reg[14]  ( .D(\DP/RegME/N17 ), .CK(n2455), .Q(
        \DP/RegME_out[14] ) );
  DFF_X1 \DP/RegB/DOUT_reg[15]  ( .D(\DP/RegB/N18 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[15] ) );
  DFF_X1 \DP/RegME/DOUT_reg[15]  ( .D(\DP/RegME/N18 ), .CK(n2453), .Q(
        \DP/RegME_out[15] ) );
  DFF_X1 \DP/RegB/DOUT_reg[16]  ( .D(\DP/RegB/N19 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[16] ) );
  DFF_X1 \DP/RegME/DOUT_reg[16]  ( .D(\DP/RegME/N19 ), .CK(n2455), .Q(
        \DP/RegME_out[16] ) );
  DFF_X1 \DP/RegB/DOUT_reg[17]  ( .D(\DP/RegB/N20 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[17] ) );
  DFF_X1 \DP/RegME/DOUT_reg[17]  ( .D(\DP/RegME/N20 ), .CK(n2454), .Q(
        \DP/RegME_out[17] ) );
  DFF_X1 \DP/RegB/DOUT_reg[18]  ( .D(\DP/RegB/N21 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[18] ) );
  DFF_X1 \DP/RegME/DOUT_reg[18]  ( .D(\DP/RegME/N21 ), .CK(n2452), .Q(
        \DP/RegME_out[18] ) );
  DFF_X1 \DP/RegB/DOUT_reg[19]  ( .D(\DP/RegB/N22 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[19] ) );
  DFF_X1 \DP/RegME/DOUT_reg[19]  ( .D(\DP/RegME/N22 ), .CK(n2454), .Q(
        \DP/RegME_out[19] ) );
  DFF_X1 \DP/RegB/DOUT_reg[20]  ( .D(\DP/RegB/N23 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[20] ) );
  DFF_X1 \DP/RegME/DOUT_reg[20]  ( .D(\DP/RegME/N23 ), .CK(n2454), .Q(
        \DP/RegME_out[20] ) );
  DFF_X1 \DP/RegB/DOUT_reg[21]  ( .D(\DP/RegB/N24 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[21] ) );
  DFF_X1 \DP/RegME/DOUT_reg[21]  ( .D(\DP/RegME/N24 ), .CK(n2453), .Q(
        \DP/RegME_out[21] ) );
  DFF_X1 \DP/RegB/DOUT_reg[22]  ( .D(\DP/RegB/N25 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[22] ) );
  DFF_X1 \DP/RegME/DOUT_reg[22]  ( .D(\DP/RegME/N25 ), .CK(n2455), .Q(
        \DP/RegME_out[22] ) );
  DFF_X1 \DP/RegB/DOUT_reg[23]  ( .D(\DP/RegB/N26 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[23] ) );
  DFF_X1 \DP/RegME/DOUT_reg[23]  ( .D(\DP/RegME/N26 ), .CK(n2454), .Q(
        \DP/RegME_out[23] ) );
  DFF_X1 \DP/RegB/DOUT_reg[24]  ( .D(\DP/RegB/N27 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[24] ) );
  DFF_X1 \DP/RegME/DOUT_reg[24]  ( .D(\DP/RegME/N27 ), .CK(n2453), .Q(
        \DP/RegME_out[24] ) );
  DFF_X1 \DP/RegB/DOUT_reg[25]  ( .D(\DP/RegB/N28 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[25] ) );
  DFF_X1 \DP/RegME/DOUT_reg[25]  ( .D(\DP/RegME/N28 ), .CK(n2454), .Q(
        \DP/RegME_out[25] ) );
  DFF_X1 \DP/RegB/DOUT_reg[26]  ( .D(\DP/RegB/N29 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[26] ) );
  DFF_X1 \DP/RegME/DOUT_reg[26]  ( .D(\DP/RegME/N29 ), .CK(n2452), .Q(
        \DP/RegME_out[26] ) );
  DFF_X1 \DP/RegB/DOUT_reg[27]  ( .D(\DP/RegB/N30 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[27] ) );
  DFF_X1 \DP/RegME/DOUT_reg[27]  ( .D(\DP/RegME/N30 ), .CK(n2455), .Q(
        \DP/RegME_out[27] ) );
  DFF_X1 \DP/RegB/DOUT_reg[28]  ( .D(\DP/RegB/N31 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[28] ) );
  DFF_X1 \DP/RegME/DOUT_reg[28]  ( .D(\DP/RegME/N31 ), .CK(n2452), .Q(
        \DP/RegME_out[28] ) );
  DFF_X1 \DP/RegB/DOUT_reg[29]  ( .D(\DP/RegB/N32 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[29] ) );
  DFF_X1 \DP/RegME/DOUT_reg[29]  ( .D(\DP/RegME/N32 ), .CK(\DP/RegLMD/net2366 ), .Q(\DP/RegME_out[29] ) );
  DFF_X1 \DP/RegB/DOUT_reg[30]  ( .D(\DP/RegB/N33 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[30] ) );
  DFF_X1 \DP/RegME/DOUT_reg[30]  ( .D(\DP/RegME/N33 ), .CK(n2455), .Q(
        \DP/RegME_out[30] ) );
  DFF_X1 \DP/RegB/DOUT_reg[31]  ( .D(\DP/RegB/N34 ), .CK(\DP/RegB/net2366 ), 
        .Q(\DP/RegB_out[31] ) );
  DFF_X1 \DP/RegME/DOUT_reg[31]  ( .D(\DP/RegME/N34 ), .CK(n2454), .Q(
        \DP/RegME_out[31] ) );
  DFF_X1 \DP/RegA/DOUT_reg[0]  ( .D(\DP/RegA/N3 ), .CK(\DP/RegA/net2366 ), .Q(
        \DP/RegA_out[0] ) );
  DFF_X1 \DP/RegA/DOUT_reg[1]  ( .D(\DP/RegA/N4 ), .CK(\DP/RegA/net2366 ), .Q(
        \DP/RegA_out[1] ) );
  DFF_X1 \DP/RegA/DOUT_reg[2]  ( .D(\DP/RegA/N5 ), .CK(\DP/RegA/net2366 ), .Q(
        \DP/RegA_out[2] ) );
  DFF_X1 \DP/RegA/DOUT_reg[3]  ( .D(\DP/RegA/N6 ), .CK(\DP/RegA/net2366 ), .Q(
        \DP/RegA_out[3] ) );
  DFF_X1 \DP/RegA/DOUT_reg[4]  ( .D(\DP/RegA/N7 ), .CK(\DP/RegA/net2366 ), .Q(
        \DP/RegA_out[4] ) );
  DFF_X1 \DP/RegA/DOUT_reg[5]  ( .D(\DP/RegA/N8 ), .CK(\DP/RegA/net2366 ), .Q(
        \DP/RegA_out[5] ) );
  DFF_X1 \DP/RegA/DOUT_reg[6]  ( .D(\DP/RegA/N9 ), .CK(\DP/RegA/net2366 ), .Q(
        \DP/RegA_out[6] ) );
  DFF_X1 \DP/RegA/DOUT_reg[7]  ( .D(\DP/RegA/N10 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[7] ) );
  DFF_X1 \DP/RegA/DOUT_reg[8]  ( .D(\DP/RegA/N11 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[8] ) );
  DFF_X1 \DP/RegA/DOUT_reg[9]  ( .D(\DP/RegA/N12 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[9] ) );
  DFF_X1 \DP/RegA/DOUT_reg[10]  ( .D(\DP/RegA/N13 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[10] ) );
  DFF_X1 \DP/RegA/DOUT_reg[11]  ( .D(\DP/RegA/N14 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[11] ) );
  DFF_X1 \DP/RegA/DOUT_reg[12]  ( .D(\DP/RegA/N15 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[12] ) );
  DFF_X1 \DP/RegA/DOUT_reg[13]  ( .D(\DP/RegA/N16 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[13] ) );
  DFF_X1 \DP/RegA/DOUT_reg[14]  ( .D(\DP/RegA/N17 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[14] ) );
  DFF_X1 \DP/RegA/DOUT_reg[15]  ( .D(\DP/RegA/N18 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[15] ) );
  DFF_X1 \DP/RegA/DOUT_reg[16]  ( .D(\DP/RegA/N19 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[16] ) );
  DFF_X1 \DP/RegA/DOUT_reg[17]  ( .D(\DP/RegA/N20 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[17] ) );
  DFF_X1 \DP/RegA/DOUT_reg[18]  ( .D(\DP/RegA/N21 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[18] ) );
  DFF_X1 \DP/RegA/DOUT_reg[19]  ( .D(\DP/RegA/N22 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[19] ) );
  DFF_X1 \DP/RegA/DOUT_reg[20]  ( .D(\DP/RegA/N23 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[20] ) );
  DFF_X1 \DP/RegA/DOUT_reg[21]  ( .D(\DP/RegA/N24 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[21] ) );
  DFF_X1 \DP/RegA/DOUT_reg[22]  ( .D(\DP/RegA/N25 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[22] ) );
  DFF_X1 \DP/RegA/DOUT_reg[23]  ( .D(\DP/RegA/N26 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[23] ) );
  DFF_X1 \DP/RegA/DOUT_reg[24]  ( .D(\DP/RegA/N27 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[24] ) );
  DFF_X1 \DP/RegA/DOUT_reg[25]  ( .D(\DP/RegA/N28 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[25] ) );
  DFF_X1 \DP/RegA/DOUT_reg[26]  ( .D(\DP/RegA/N29 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[26] ) );
  DFF_X1 \DP/RegA/DOUT_reg[27]  ( .D(\DP/RegA/N30 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[27] ) );
  DFF_X1 \DP/RegA/DOUT_reg[28]  ( .D(\DP/RegA/N31 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[28] ) );
  DFF_X1 \DP/RegA/DOUT_reg[29]  ( .D(\DP/RegA/N32 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[29] ) );
  DFF_X1 \DP/RegA/DOUT_reg[30]  ( .D(\DP/RegA/N33 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[30] ) );
  DFF_X1 \DP/RegA/DOUT_reg[31]  ( .D(\DP/RegA/N34 ), .CK(\DP/RegA/net2366 ), 
        .Q(\DP/RegA_out[31] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[31]  ( .D(\DP/RegA1/N34 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[31] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[31]  ( .D(\DP/RegNPC1/N34 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[31] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[31]  ( .D(\DP/A[31] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[31] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[31]  ( .D(n106), .GN(n2447), .Q(n56) );
  DLH_X1 \DP/ALU0/s_SIGN_reg  ( .G(\DP/ALU0/N91 ), .D(n105), .Q(
        \DP/ALU0/s_SIGN ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[0]  ( .D(\DP/RegALU1/N3 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[0]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[0]  ( .D(\DP/RegALU2/N3 ), .CK(n2454), .Q(
        \DP/RegALU2_out[0] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[0]  ( .D(\DP/RegA1/N3 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[0] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[0]  ( .G(n2340), .D(\DP/B[0] ), .Q(
        \DP/ALU0/S_B_LHI[0] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[0]  ( .G(n2440), .D(\DP/B[0] ), .Q(
        \DP/ALU0/S_B_MULT[0] ) );
  DLL_X1 \DP/ALU0/S_B_SHIFT_reg[0]  ( .D(\DP/B[0] ), .GN(n2444), .Q(
        \DP/ALU0/S_B_SHIFT[0] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[0]  ( .D(\DP/B[0] ), .GN(n2447), .Q(
        \DP/ALU0/S_B_LOGIC[0] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[0]  ( .G(n2457), .D(\DP/ALU0/N54 ), .Q(
        \DP/ALU0/S_B_ADDER[0] ) );
  DFF_X1 \PC/DOUT_reg[0]  ( .D(\PC/N3 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IROM_ADDR[0]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[0]  ( .D(\PC/N3 ), .CK(\DP/RegNPC/net2366 ), .Q(
        \DP/NPC1[0] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[0]  ( .D(\DP/RegNPC1/N3 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[0] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[0]  ( .G(n2440), .D(\DP/A[0] ), .Q(
        \DP/ALU0/MULT/SHIFTERi_0/N19 ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[0]  ( .D(\DP/A[0] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[0] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[0]  ( .D(\DP/A[0] ), .GN(n2447), .Q(
        \DP/ALU0/s_A_LOGIC[0] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[0]  ( .G(n2457), .D(\DP/ALU0/N22 ), .Q(
        \DP/ALU0/s_A_ADDER[0] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[5]  ( .D(\DP/RegALU1/N8 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[5]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[5]  ( .D(\DP/RegALU2/N8 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegALU2_out[5] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[5]  ( .G(n2340), .D(\DP/B[5] ), .Q(
        \DP/ALU0/S_B_LHI[5] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[5]  ( .G(n2440), .D(\DP/B[5] ), .Q(
        \DP/ALU0/S_B_MULT[5] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[5]  ( .D(\DP/B[5] ), .GN(n2447), .Q(
        \DP/ALU0/S_B_LOGIC[5] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[5]  ( .G(n2457), .D(\DP/ALU0/N59 ), .Q(
        \DP/ALU0/S_B_ADDER[5] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[5]  ( .D(\DP/RegA1/N8 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[5] ) );
  DFF_X1 \PC/DOUT_reg[5]  ( .D(\PC/N8 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IROM_ADDR[5]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[5]  ( .D(\PC/N8 ), .CK(\DP/RegNPC/net2366 ), .Q(
        \DP/NPC1[5] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[5]  ( .D(\DP/RegNPC1/N8 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[5] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[5]  ( .G(n2441), .D(n186), .Q(n55) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[5]  ( .D(\DP/A[5] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[5] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[5]  ( .D(\DP/A[5] ), .GN(n2447), .Q(
        \DP/ALU0/s_A_LOGIC[5] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[5]  ( .G(n2457), .D(\DP/ALU0/N27 ), .Q(
        \DP/ALU0/s_A_ADDER[5] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[8]  ( .D(\DP/RegALU1/N11 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[8]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[8]  ( .D(\DP/RegALU2/N11 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegALU2_out[8] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[8]  ( .G(n2340), .D(\DP/B[8] ), .Q(
        \DP/ALU0/S_B_LHI[8] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[8]  ( .G(n2440), .D(n176), .Q(n54) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[8]  ( .D(\DP/B[8] ), .GN(n2447), .Q(
        \DP/ALU0/S_B_LOGIC[8] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[8]  ( .D(\DP/RegA1/N11 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[8] ) );
  DFF_X1 \PC/DOUT_reg[8]  ( .D(\PC/N11 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IROM_ADDR[8]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[8]  ( .D(\PC/N11 ), .CK(\DP/RegNPC/net2366 ), .Q(
        \DP/NPC1[8] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[8]  ( .D(\DP/RegNPC1/N11 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[8] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[8]  ( .G(n2441), .D(n175), .Q(n53) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[8]  ( .D(\DP/A[8] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[8] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[8]  ( .D(\DP/A[8] ), .GN(n2447), .Q(
        \DP/ALU0/s_A_LOGIC[8] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[8]  ( .G(n2457), .D(\DP/ALU0/N30 ), .Q(
        \DP/ALU0/s_A_ADDER[8] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[9]  ( .D(\DP/RegALU1/N12 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[9]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[9]  ( .D(\DP/RegALU2/N12 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegALU2_out[9] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[9]  ( .G(n2340), .D(\DP/B[9] ), .Q(
        \DP/ALU0/S_B_LHI[9] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[9]  ( .G(n2440), .D(n173), .Q(n52) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[9]  ( .D(\DP/B[9] ), .GN(n2447), .Q(
        \DP/ALU0/S_B_LOGIC[9] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[9]  ( .D(\DP/RegA1/N12 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[9] ) );
  DFF_X1 \PC/DOUT_reg[9]  ( .D(\PC/N12 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IROM_ADDR[9]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[9]  ( .D(\PC/N12 ), .CK(\DP/RegNPC/net2366 ), .Q(
        \DP/NPC1[9] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[9]  ( .D(\DP/RegNPC1/N12 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[9] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[9]  ( .G(n2441), .D(\DP/A[9] ), .Q(
        \DP/ALU0/s_A_MULT[9] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[9]  ( .D(\DP/A[9] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[9] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[9]  ( .D(\DP/A[9] ), .GN(n2447), .Q(
        \DP/ALU0/s_A_LOGIC[9] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[9]  ( .G(n2457), .D(\DP/ALU0/N31 ), .Q(
        \DP/ALU0/s_A_ADDER[9] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[11]  ( .D(\DP/RegALU1/N14 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[11]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[11]  ( .D(\DP/RegALU2/N14 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegALU2_out[11] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[11]  ( .G(n2340), .D(\DP/B[11] ), .Q(
        \DP/ALU0/S_B_LHI[11] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[11]  ( .G(n2440), .D(n167), .Q(n51) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[11]  ( .D(\DP/B[11] ), .GN(n2447), .Q(
        \DP/ALU0/S_B_LOGIC[11] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[11]  ( .D(\DP/RegA1/N14 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[11] ) );
  DFF_X1 \PC/DOUT_reg[11]  ( .D(\PC/N14 ), .CK(n2456), .Q(IROM_ADDR[11]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[11]  ( .D(\PC/N14 ), .CK(\DP/RegNPC/net2366 ), 
        .Q(\DP/NPC1[11] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[11]  ( .D(\DP/RegNPC1/N14 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[11] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[11]  ( .G(n2440), .D(\DP/A[11] ), .Q(
        \DP/ALU0/s_A_MULT[11] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[11]  ( .D(\DP/A[11] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[11] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[11]  ( .D(\DP/A[11] ), .GN(n2447), .Q(
        \DP/ALU0/s_A_LOGIC[11] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[11]  ( .G(n2457), .D(\DP/ALU0/N33 ), .Q(
        \DP/ALU0/s_A_ADDER[11] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[14]  ( .D(\DP/RegALU1/N17 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[14] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[14]  ( .D(\DP/RegALU2/N17 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegALU2_out[14] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[14]  ( .G(n2340), .D(\DP/B[14] ), .Q(
        \DP/ALU0/S_B_LHI[14] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[14]  ( .G(n2440), .D(n158), .Q(n50) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[14]  ( .D(\DP/B[14] ), .GN(n2447), .Q(
        \DP/ALU0/S_B_LOGIC[14] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[14]  ( .D(\DP/RegA1/N17 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[14] ) );
  DFF_X1 \PC/DOUT_reg[14]  ( .D(\PC/N17 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[14]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[14]  ( .D(\PC/N17 ), .CK(\DP/RegNPC/net2366 ), 
        .Q(\DP/NPC1[14] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[14]  ( .D(\DP/RegNPC1/N17 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[14] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[14]  ( .G(n2441), .D(n157), .Q(n49) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[14]  ( .D(\DP/A[14] ), .GN(n4740), .Q(
        \DP/ALU0/s_A_SHIFT[14] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[14]  ( .D(\DP/A[14] ), .GN(n2447), .Q(
        \DP/ALU0/s_A_LOGIC[14] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[14]  ( .G(n2457), .D(\DP/ALU0/N36 ), .Q(
        \DP/ALU0/s_A_ADDER[14] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[15]  ( .D(\DP/RegALU1/N18 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[15] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[15]  ( .D(\DP/RegALU2/N18 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegALU2_out[15] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[15]  ( .G(n2340), .D(\DP/B[15] ), .Q(
        \DP/ALU0/S_B_LHI[15] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[15]  ( .G(n2440), .D(n155), .Q(n48) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[15]  ( .D(\DP/B[15] ), .GN(n2447), .Q(
        \DP/ALU0/S_B_LOGIC[15] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[15]  ( .D(\DP/RegA1/N18 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[15] ) );
  DFF_X1 \PC/DOUT_reg[15]  ( .D(\PC/N18 ), .CK(n2456), .Q(w_PC_OUT[15]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[15]  ( .D(\PC/N18 ), .CK(\DP/RegNPC/net2366 ), 
        .Q(\DP/NPC1[15] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[15]  ( .D(\DP/RegNPC1/N18 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[15] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[15]  ( .G(n2441), .D(n154), .Q(n47) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[15]  ( .D(\DP/A[15] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[15] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[15]  ( .D(\DP/A[15] ), .GN(n2447), .Q(
        \DP/ALU0/s_A_LOGIC[15] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[15]  ( .G(n2457), .D(\DP/ALU0/N37 ), .Q(
        \DP/ALU0/s_A_ADDER[15] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[19]  ( .D(\DP/RegALU1/N22 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[19] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[19]  ( .D(\DP/RegALU2/N22 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegALU2_out[19] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[19]  ( .D(n143), .GN(n2447), .Q(n46) );
  DFF_X1 \DP/RegA1/DOUT_reg[19]  ( .D(\DP/RegA1/N22 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[19] ) );
  DFF_X1 \PC/DOUT_reg[19]  ( .D(\PC/N22 ), .CK(n2456), .Q(w_PC_OUT[19]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[19]  ( .D(\PC/N22 ), .CK(\DP/RegNPC/net2366 ), 
        .Q(\DP/NPC1[19] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[19]  ( .D(\DP/RegNPC1/N22 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[19] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[19]  ( .D(n142), .GN(n4740), .Q(n45) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[19]  ( .D(n142), .GN(n2446), .Q(n44) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[19]  ( .G(n2457), .D(\DP/ALU0/N41 ), .Q(
        \DP/ALU0/s_A_ADDER[19] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[23]  ( .D(\DP/RegALU2/N26 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegALU2_out[23] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[23]  ( .D(n131), .GN(n2446), .Q(n43) );
  DFF_X1 \DP/RegA1/DOUT_reg[23]  ( .D(\DP/RegA1/N26 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[23] ) );
  DFF_X1 \PC/DOUT_reg[23]  ( .D(\PC/N26 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[23]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[23]  ( .D(\PC/N26 ), .CK(n2456), .Q(\DP/NPC1[23] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[23]  ( .D(\DP/RegNPC1/N26 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[23] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[23]  ( .D(n130), .GN(n2444), .Q(n42) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[23]  ( .D(n130), .GN(n2447), .Q(n41) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[23]  ( .G(n2457), .D(\DP/ALU0/N45 ), .Q(
        \DP/ALU0/s_A_ADDER[23] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[26]  ( .D(\DP/RegALU1/N29 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[26] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[26]  ( .D(\DP/RegALU2/N29 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegALU2_out[26] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[26]  ( .D(n122), .GN(n2446), .Q(n40) );
  DFF_X1 \DP/RegA1/DOUT_reg[26]  ( .D(\DP/RegA1/N29 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[26] ) );
  DFF_X1 \PC/DOUT_reg[26]  ( .D(\PC/N29 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[26]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[26]  ( .D(\PC/N29 ), .CK(n2456), .Q(\DP/NPC1[26] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[26]  ( .D(\DP/RegNPC1/N29 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[26] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[26]  ( .D(\DP/A[26] ), .GN(n4740), .Q(
        \DP/ALU0/s_A_SHIFT[26] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[26]  ( .D(n121), .GN(n2447), .Q(n39) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[26]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N48 ), 
        .Q(\DP/ALU0/s_A_ADDER[26] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[27]  ( .D(\DP/RegALU1/N30 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[27] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[27]  ( .D(\DP/RegALU2/N30 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegALU2_out[27] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[27]  ( .D(n119), .GN(n2447), .Q(n38) );
  DFF_X1 \DP/RegA1/DOUT_reg[27]  ( .D(\DP/RegA1/N30 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[27] ) );
  DFF_X1 \PC/DOUT_reg[27]  ( .D(\PC/N30 ), .CK(n2456), .Q(w_PC_OUT[27]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[27]  ( .D(\PC/N30 ), .CK(\DP/RegNPC/net2366 ), 
        .Q(\DP/NPC1[27] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[27]  ( .D(\DP/RegNPC1/N30 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[27] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[27]  ( .D(\DP/A[27] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[27] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[27]  ( .D(n118), .GN(n2446), .Q(n37) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[27]  ( .G(n2457), .D(\DP/ALU0/N49 ), .Q(
        \DP/ALU0/s_A_ADDER[27] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[29]  ( .D(\DP/RegALU1/N32 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[29] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[29]  ( .D(\DP/RegALU2/N32 ), .CK(
        \DP/RegLMD/net2366 ), .Q(\DP/RegALU2_out[29] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[29]  ( .D(n113), .GN(n2446), .Q(n36) );
  DFF_X1 \DP/RegA1/DOUT_reg[29]  ( .D(\DP/RegA1/N32 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[29] ) );
  DFF_X1 \PC/DOUT_reg[29]  ( .D(\PC/N32 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[29]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[29]  ( .D(\PC/N32 ), .CK(n2456), .Q(\DP/NPC1[29] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[29]  ( .D(\DP/RegNPC1/N32 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[29] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[29]  ( .D(\DP/A[29] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[29] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[29]  ( .D(n112), .GN(n2447), .Q(n35) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[29]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N51 ), 
        .Q(\DP/ALU0/s_A_ADDER[29] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[30]  ( .D(\DP/RegALU1/N33 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[30] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[30]  ( .D(\DP/RegALU2/N33 ), .CK(n2455), .Q(
        \DP/RegALU2_out[30] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[30]  ( .D(n110), .GN(n2446), .Q(n34) );
  DFF_X1 \DP/RegA1/DOUT_reg[30]  ( .D(\DP/RegA1/N33 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[30] ) );
  DFF_X1 \PC/DOUT_reg[30]  ( .D(\PC/N33 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[30]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[30]  ( .D(\PC/N33 ), .CK(n2456), .Q(\DP/NPC1[30] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[30]  ( .D(\DP/RegNPC1/N33 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[30] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[30]  ( .D(\DP/A[30] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[30] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[28]  ( .D(\DP/RegALU1/N31 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[28] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[28]  ( .D(\DP/RegALU2/N31 ), .CK(n2454), .Q(
        \DP/RegALU2_out[28] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[28]  ( .D(n116), .GN(n2447), .Q(n33) );
  DFF_X1 \DP/RegA1/DOUT_reg[28]  ( .D(\DP/RegA1/N31 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[28] ) );
  DFF_X1 \DP/RegNPC/DOUT_reg[28]  ( .D(\PC/N31 ), .CK(n2456), .Q(\DP/NPC1[28] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[28]  ( .D(\DP/RegNPC1/N31 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[28] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[28]  ( .D(\DP/A[28] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[28] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[25]  ( .D(\DP/RegALU1/N28 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[25] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[25]  ( .D(\DP/RegALU2/N28 ), .CK(n2452), .Q(
        \DP/RegALU2_out[25] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[25]  ( .D(n125), .GN(n2447), .Q(n32) );
  DFF_X1 \DP/RegA1/DOUT_reg[25]  ( .D(\DP/RegA1/N28 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[25] ) );
  DFF_X1 \PC/DOUT_reg[25]  ( .D(\PC/N28 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[25]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[25]  ( .D(\PC/N28 ), .CK(\DP/RegNPC/net2366 ), 
        .Q(\DP/NPC1[25] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[25]  ( .D(\DP/RegNPC1/N28 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[25] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[25]  ( .D(\DP/A[25] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[25] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[6]  ( .D(\DP/RegALU1/N9 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[6]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[6]  ( .D(\DP/RegALU2/N9 ), .CK(n2453), .Q(
        \DP/RegALU2_out[6] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[6]  ( .G(n2340), .D(\DP/B[6] ), .Q(
        \DP/ALU0/S_B_LHI[6] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[6]  ( .G(n2440), .D(n183), .Q(n31) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[6]  ( .D(\DP/B[6] ), .GN(n2446), .Q(
        \DP/ALU0/S_B_LOGIC[6] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[6]  ( .G(n2441), .D(n182), .Q(n30) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[6]  ( .D(\DP/A[6] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[6] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[6]  ( .D(\DP/A[6] ), .GN(n2446), .Q(
        \DP/ALU0/s_A_LOGIC[6] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[6]  ( .G(n2457), .D(\DP/ALU0/N28 ), .Q(
        \DP/ALU0/s_A_ADDER[6] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[7]  ( .D(\DP/RegALU1/N10 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[7]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[7]  ( .D(\DP/RegALU2/N10 ), .CK(n2453), .Q(
        \DP/RegALU2_out[7] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[7]  ( .G(n2340), .D(\DP/B[7] ), .Q(
        \DP/ALU0/S_B_LHI[7] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[7]  ( .G(n2440), .D(n179), .Q(n29) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[7]  ( .D(\DP/B[7] ), .GN(n2447), .Q(
        \DP/ALU0/S_B_LOGIC[7] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[7]  ( .D(\DP/RegA1/N10 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[7] ) );
  DFF_X1 \PC/DOUT_reg[7]  ( .D(\PC/N10 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IROM_ADDR[7]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[7]  ( .D(\PC/N10 ), .CK(n2456), .Q(\DP/NPC1[7] )
         );
  DFF_X1 \DP/RegNPC1/DOUT_reg[7]  ( .D(\DP/RegNPC1/N10 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[7] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[7]  ( .G(n2440), .D(n178), .Q(n28) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[7]  ( .D(\DP/A[7] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[7] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[4]  ( .D(\DP/RegALU1/N7 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[4]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[4]  ( .D(\DP/RegALU2/N7 ), .CK(n2455), .Q(
        \DP/RegALU2_out[4] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[4]  ( .G(n2340), .D(\DP/B[4] ), .Q(
        \DP/ALU0/S_B_LHI[4] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[4]  ( .G(n2440), .D(\DP/B[4] ), .Q(
        \DP/ALU0/S_B_MULT[4] ) );
  DLL_X1 \DP/ALU0/S_B_SHIFT_reg[4]  ( .D(\DP/B[4] ), .GN(n2444), .Q(
        \DP/ALU0/S_B_SHIFT[4] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[4]  ( .D(\DP/B[4] ), .GN(n2446), .Q(
        \DP/ALU0/S_B_LOGIC[4] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[4]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N58 ), 
        .Q(\DP/ALU0/S_B_ADDER[4] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[4]  ( .D(\DP/RegA1/N7 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[4] ) );
  DFF_X1 \PC/DOUT_reg[4]  ( .D(\PC/N7 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IROM_ADDR[4]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[4]  ( .D(\PC/N7 ), .CK(\DP/RegNPC/net2366 ), .Q(
        \DP/NPC1[4] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[4]  ( .D(\DP/RegNPC1/N7 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[4] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[4]  ( .G(n2440), .D(\DP/A[4] ), .Q(
        \DP/ALU0/s_A_MULT[4] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[4]  ( .D(\DP/A[4] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[4] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[1]  ( .D(\DP/RegALU1/N4 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[1]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[1]  ( .D(\DP/RegALU2/N4 ), .CK(n2454), .Q(
        \DP/RegALU2_out[1] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[1]  ( .D(\DP/RegA1/N4 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[1] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[1]  ( .G(n2340), .D(\DP/B[1] ), .Q(
        \DP/ALU0/S_B_LHI[1] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[1]  ( .G(n2440), .D(\DP/B[1] ), .Q(
        \DP/ALU0/S_B_MULT[1] ) );
  DLL_X1 \DP/ALU0/S_B_SHIFT_reg[1]  ( .D(\DP/B[1] ), .GN(n2444), .Q(
        \DP/ALU0/S_B_SHIFT[1] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[1]  ( .D(\DP/B[1] ), .GN(n2447), .Q(
        \DP/ALU0/S_B_LOGIC[1] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[1]  ( .G(n2457), .D(\DP/ALU0/N55 ), .Q(
        \DP/ALU0/S_B_ADDER[1] ) );
  DFF_X1 \PC/DOUT_reg[1]  ( .D(\PC/N4 ), .CK(n2456), .Q(IROM_ADDR[1]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[1]  ( .D(\PC/N4 ), .CK(\DP/RegNPC/net2366 ), .Q(
        \DP/NPC1[1] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[1]  ( .D(\DP/RegNPC1/N4 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[1] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[1]  ( .G(n2440), .D(\DP/A[1] ), .Q(
        \DP/ALU0/s_A_MULT[1] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[1]  ( .D(\DP/A[1] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[1] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[1]  ( .D(\DP/A[1] ), .GN(n2447), .Q(
        \DP/ALU0/s_A_LOGIC[1] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[1]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N23 ), 
        .Q(\DP/ALU0/s_A_ADDER[1] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[2]  ( .D(\DP/RegALU1/N5 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[2]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[2]  ( .D(\DP/RegALU2/N5 ), .CK(n2452), .Q(
        \DP/RegALU2_out[2] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[2]  ( .D(\DP/RegA1/N5 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[2] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[2]  ( .G(n2340), .D(\DP/B[2] ), .Q(
        \DP/ALU0/S_B_LHI[2] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[2]  ( .G(n2440), .D(\DP/B[2] ), .Q(
        \DP/ALU0/S_B_MULT[2] ) );
  DLL_X1 \DP/ALU0/S_B_SHIFT_reg[2]  ( .D(\DP/B[2] ), .GN(n4740), .Q(
        \DP/ALU0/S_B_SHIFT[2] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[2]  ( .D(\DP/B[2] ), .GN(n2446), .Q(
        \DP/ALU0/S_B_LOGIC[2] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[2]  ( .G(n2457), .D(\DP/ALU0/N56 ), .Q(
        \DP/ALU0/S_B_ADDER[2] ) );
  DFF_X1 \PC/DOUT_reg[2]  ( .D(\PC/N5 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IROM_ADDR[2]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[2]  ( .D(\PC/N5 ), .CK(n2456), .Q(\DP/NPC1[2] )
         );
  DFF_X1 \DP/RegNPC1/DOUT_reg[2]  ( .D(\DP/RegNPC1/N5 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[2] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[2]  ( .G(n2440), .D(\DP/A[2] ), .Q(
        \DP/ALU0/s_A_MULT[2] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[2]  ( .D(\DP/A[2] ), .GN(n4740), .Q(
        \DP/ALU0/s_A_SHIFT[2] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[2]  ( .D(\DP/A[2] ), .GN(n2446), .Q(
        \DP/ALU0/s_A_LOGIC[2] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[2]  ( .G(\DP/ALU0/N21 ), .D(n196), .Q(
        \DP/ALU0/s_A_ADDER[2] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[3]  ( .D(\DP/RegALU1/N6 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[3]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[3]  ( .D(\DP/RegALU2/N6 ), .CK(n2455), .Q(
        \DP/RegALU2_out[3] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[3]  ( .D(\DP/RegA1/N6 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[3] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[3]  ( .G(n2340), .D(\DP/B[3] ), .Q(
        \DP/ALU0/S_B_LHI[3] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[3]  ( .G(n2440), .D(\DP/B[3] ), .Q(
        \DP/ALU0/S_B_MULT[3] ) );
  DLL_X1 \DP/ALU0/S_B_SHIFT_reg[3]  ( .D(\DP/B[3] ), .GN(n4740), .Q(
        \DP/ALU0/S_B_SHIFT[3] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[3]  ( .D(\DP/B[3] ), .GN(n2446), .Q(
        \DP/ALU0/S_B_LOGIC[3] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[3]  ( .G(n2457), .D(\DP/ALU0/N57 ), .Q(
        \DP/ALU0/S_B_ADDER[3] ) );
  DFF_X1 \PC/DOUT_reg[3]  ( .D(\PC/N6 ), .CK(\DP/RegNPC/net2366 ), .Q(
        IROM_ADDR[3]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[3]  ( .D(\PC/N6 ), .CK(n2456), .Q(\DP/NPC1[3] )
         );
  DFF_X1 \DP/RegNPC1/DOUT_reg[3]  ( .D(\DP/RegNPC1/N6 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[3] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[3]  ( .G(n2440), .D(\DP/A[3] ), .Q(
        \DP/ALU0/s_A_MULT[3] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[3]  ( .D(\DP/A[3] ), .GN(n4740), .Q(
        \DP/ALU0/s_A_SHIFT[3] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[24]  ( .D(\DP/RegALU2/N27 ), .CK(n2453), .Q(
        \DP/RegALU2_out[24] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[24]  ( .D(n128), .GN(n2446), .Q(n27) );
  DFF_X1 \DP/RegA1/DOUT_reg[24]  ( .D(\DP/RegA1/N27 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[24] ) );
  DFF_X1 \PC/DOUT_reg[24]  ( .D(\PC/N27 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[24]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[24]  ( .D(\PC/N27 ), .CK(\DP/RegNPC/net2366 ), 
        .Q(\DP/NPC1[24] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[24]  ( .D(\DP/RegNPC1/N27 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[24] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[24]  ( .D(\DP/A[24] ), .GN(n4740), .Q(
        \DP/ALU0/s_A_SHIFT[24] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[21]  ( .D(\DP/RegALU2/N24 ), .CK(n2455), .Q(
        \DP/RegALU2_out[21] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[21]  ( .D(n137), .GN(n2446), .Q(n26) );
  DFF_X1 \DP/RegA1/DOUT_reg[21]  ( .D(\DP/RegA1/N24 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[21] ) );
  DFF_X1 \PC/DOUT_reg[21]  ( .D(\PC/N24 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[21]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[21]  ( .D(\PC/N24 ), .CK(n2456), .Q(\DP/NPC1[21] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[21]  ( .D(\DP/RegNPC1/N24 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[21] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[21]  ( .D(n136), .GN(n4740), .Q(n25) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[21]  ( .D(n136), .GN(n2446), .Q(n24) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[21]  ( .G(n2457), .D(\DP/ALU0/N43 ), .Q(
        \DP/ALU0/s_A_ADDER[21] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[22]  ( .D(\DP/RegALU1/N25 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[22] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[22]  ( .D(\DP/RegALU2/N25 ), .CK(n2455), .Q(
        \DP/RegALU2_out[22] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[22]  ( .D(n134), .GN(n2446), .Q(n23) );
  DFF_X1 \DP/RegA1/DOUT_reg[22]  ( .D(\DP/RegA1/N25 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[22] ) );
  DFF_X1 \PC/DOUT_reg[22]  ( .D(\PC/N25 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[22]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[22]  ( .D(\PC/N25 ), .CK(n2456), .Q(\DP/NPC1[22] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[22]  ( .D(\DP/RegNPC1/N25 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[22] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[22]  ( .D(n133), .GN(n4740), .Q(n22) );
  DFF_X1 \DP/RegALU2/DOUT_reg[20]  ( .D(\DP/RegALU2/N23 ), .CK(n2454), .Q(
        \DP/RegALU2_out[20] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[20]  ( .D(n140), .GN(n2446), .Q(n21) );
  DFF_X1 \DP/RegA1/DOUT_reg[20]  ( .D(\DP/RegA1/N23 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[20] ) );
  DFF_X1 \PC/DOUT_reg[20]  ( .D(\PC/N23 ), .CK(n2456), .Q(w_PC_OUT[20]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[20]  ( .D(\PC/N23 ), .CK(\DP/RegNPC/net2366 ), 
        .Q(\DP/NPC1[20] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[20]  ( .D(\DP/RegNPC1/N23 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[20] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[20]  ( .D(n139), .GN(n2444), .Q(n20) );
  DFF_X1 \DP/RegALU1/DOUT_reg[17]  ( .D(\DP/RegALU1/N20 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[17] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[17]  ( .D(\DP/RegALU2/N20 ), .CK(n2452), .Q(
        \DP/RegALU2_out[17] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[17]  ( .D(n149), .GN(n2446), .Q(n19) );
  DFF_X1 \DP/RegA1/DOUT_reg[17]  ( .D(\DP/RegA1/N20 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[17] ) );
  DFF_X1 \PC/DOUT_reg[17]  ( .D(\PC/N20 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[17]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[17]  ( .D(\PC/N20 ), .CK(n2456), .Q(\DP/NPC1[17] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[17]  ( .D(\DP/RegNPC1/N20 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[17] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[17]  ( .D(n148), .GN(n2444), .Q(n18) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[17]  ( .D(n148), .GN(n2446), .Q(n17) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[17]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N39 ), 
        .Q(\DP/ALU0/s_A_ADDER[17] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[18]  ( .D(\DP/RegALU1/N21 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[18] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[18]  ( .D(\DP/RegALU2/N21 ), .CK(n2452), .Q(
        \DP/RegALU2_out[18] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[18]  ( .D(n146), .GN(n2446), .Q(n16) );
  DFF_X1 \PC/DOUT_reg[18]  ( .D(\PC/N21 ), .CK(n2456), .Q(w_PC_OUT[18]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[18]  ( .D(\PC/N21 ), .CK(n2456), .Q(\DP/NPC1[18] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[18]  ( .D(\DP/RegNPC1/N21 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[18] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[18]  ( .D(n145), .GN(n4740), .Q(n15) );
  DFF_X1 \DP/RegALU1/DOUT_reg[16]  ( .D(\DP/RegALU1/N19 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[16] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[16]  ( .D(\DP/RegALU2/N19 ), .CK(n2453), .Q(
        \DP/RegALU2_out[16] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[16]  ( .D(n152), .GN(n2446), .Q(n14) );
  DFF_X1 \DP/RegA1/DOUT_reg[16]  ( .D(\DP/RegA1/N19 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[16] ) );
  DFF_X1 \PC/DOUT_reg[16]  ( .D(\PC/N19 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[16]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[16]  ( .D(\PC/N19 ), .CK(\DP/RegNPC/net2366 ), 
        .Q(\DP/NPC1[16] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[16]  ( .D(\DP/RegNPC1/N19 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[16] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[16]  ( .D(n151), .GN(n4740), .Q(n13) );
  DFF_X1 \DP/RegALU1/DOUT_reg[13]  ( .D(\DP/RegALU1/N16 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[13] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[13]  ( .D(\DP/RegALU2/N16 ), .CK(n2453), .Q(
        \DP/RegALU2_out[13] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[13]  ( .G(n2340), .D(\DP/B[13] ), .Q(
        \DP/ALU0/S_B_LHI[13] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[13]  ( .G(n2440), .D(n161), .Q(n12) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[13]  ( .D(\DP/B[13] ), .GN(n2446), .Q(
        \DP/ALU0/S_B_LOGIC[13] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[13]  ( .D(\DP/RegA1/N16 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[13] ) );
  DFF_X1 \PC/DOUT_reg[13]  ( .D(\PC/N16 ), .CK(n2456), .Q(w_PC_OUT[13]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[13]  ( .D(\PC/N16 ), .CK(n2456), .Q(\DP/NPC1[13] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[13]  ( .D(\DP/RegNPC1/N16 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[13] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[13]  ( .G(n2440), .D(\DP/A[13] ), .Q(
        \DP/ALU0/s_A_MULT[13] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[13]  ( .D(\DP/A[13] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[13] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[10]  ( .D(\DP/RegALU1/N13 ), .CK(
        \DP/RegALU1/net2366 ), .Q(DRAM_ADDR[10]) );
  DFF_X1 \DP/RegALU2/DOUT_reg[10]  ( .D(\DP/RegALU2/N13 ), .CK(n2453), .Q(
        \DP/RegALU2_out[10] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[10]  ( .G(n2340), .D(\DP/B[10] ), .Q(
        \DP/ALU0/S_B_LHI[10] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[10]  ( .G(n2440), .D(n170), .Q(n11) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[10]  ( .D(\DP/B[10] ), .GN(n2446), .Q(
        \DP/ALU0/S_B_LOGIC[10] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[10]  ( .D(\DP/RegA1/N13 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[10] ) );
  DFF_X1 \PC/DOUT_reg[10]  ( .D(\PC/N13 ), .CK(n2456), .Q(IROM_ADDR[10]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[10]  ( .D(\PC/N13 ), .CK(\DP/RegNPC/net2366 ), 
        .Q(\DP/NPC1[10] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[10]  ( .D(\DP/RegNPC1/N13 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[10] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[10]  ( .G(n2440), .D(\DP/A[10] ), .Q(
        \DP/ALU0/s_A_MULT[10] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[12]  ( .G(n2457), .D(\DP/ALU0/N34 ), .Q(
        \DP/ALU0/s_A_ADDER[12] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[12]  ( .D(\DP/RegALU1/N15 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[12] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[12]  ( .D(\DP/RegALU2/N15 ), .CK(n2455), .Q(
        \DP/RegALU2_out[12] ) );
  DLH_X1 \DP/ALU0/S_B_LHI_reg[12]  ( .G(n2340), .D(\DP/B[12] ), .Q(
        \DP/ALU0/S_B_LHI[12] ) );
  DLH_X1 \DP/ALU0/S_B_MULT_reg[12]  ( .G(n2440), .D(n164), .Q(n10) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[12]  ( .D(\DP/B[12] ), .GN(n2446), .Q(
        \DP/ALU0/S_B_LOGIC[12] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[12]  ( .D(\DP/RegA1/N15 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[12] ) );
  DFF_X1 \PC/DOUT_reg[12]  ( .D(\PC/N15 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[12]) );
  DFF_X1 \DP/RegNPC/DOUT_reg[12]  ( .D(\PC/N15 ), .CK(\DP/RegNPC/net2366 ), 
        .Q(\DP/NPC1[12] ) );
  DFF_X1 \DP/RegNPC1/DOUT_reg[12]  ( .D(\DP/RegNPC1/N15 ), .CK(
        \DP/RegNPC1/net2366 ), .Q(\DP/NPC2[12] ) );
  DLH_X1 \DP/ALU0/s_A_MULT_reg[12]  ( .G(n2441), .D(\DP/A[12] ), .Q(
        \DP/ALU0/s_A_MULT[12] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[6]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N60 ), 
        .Q(\DP/ALU0/S_B_ADDER[6] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[7]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N61 ), 
        .Q(\DP/ALU0/S_B_ADDER[7] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[8]  ( .G(n2457), .D(\DP/ALU0/N62 ), .Q(
        \DP/ALU0/S_B_ADDER[8] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[9]  ( .G(n2457), .D(\DP/ALU0/N63 ), .Q(
        \DP/ALU0/S_B_ADDER[9] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[10]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N64 ), 
        .Q(\DP/ALU0/S_B_ADDER[10] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[11]  ( .G(n2457), .D(\DP/ALU0/N65 ), .Q(
        \DP/ALU0/S_B_ADDER[11] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[13]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N67 ), 
        .Q(\DP/ALU0/S_B_ADDER[13] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[12]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N66 ), 
        .Q(\DP/ALU0/S_B_ADDER[12] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[31]  ( .G(n2457), .D(\DP/ALU0/N53 ), .Q(
        \DP/ALU0/s_A_ADDER[31] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[30]  ( .G(n2457), .D(\DP/ALU0/N84 ), .Q(
        \DP/ALU0/S_B_ADDER[30] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[29]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N83 ), 
        .Q(\DP/ALU0/S_B_ADDER[29] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[28]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N82 ), 
        .Q(\DP/ALU0/S_B_ADDER[28] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[12]  ( .D(\DP/A[12] ), .GN(n4740), .Q(
        \DP/ALU0/s_A_SHIFT[12] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[12]  ( .D(\DP/A[12] ), .GN(n2446), .Q(
        \DP/ALU0/s_A_LOGIC[12] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[12]  ( .D(\DP/RegNPC2/N15 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[12] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[12]  ( .D(\DP/RegNPC3/N15 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[12] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[14]  ( .G(n2457), .D(\DP/ALU0/N68 ), .Q(
        \DP/ALU0/S_B_ADDER[14] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[15]  ( .G(n2457), .D(\DP/ALU0/N69 ), .Q(
        \DP/ALU0/S_B_ADDER[15] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[16]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N70 ), 
        .Q(\DP/ALU0/S_B_ADDER[16] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[17]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N71 ), 
        .Q(\DP/ALU0/S_B_ADDER[17] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[18]  ( .G(n2457), .D(\DP/ALU0/N72 ), .Q(
        \DP/ALU0/S_B_ADDER[18] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[19]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N73 ), 
        .Q(\DP/ALU0/S_B_ADDER[19] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[20]  ( .G(n2457), .D(\DP/ALU0/N74 ), .Q(
        \DP/ALU0/S_B_ADDER[20] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[21]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N75 ), 
        .Q(\DP/ALU0/S_B_ADDER[21] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[22]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N76 ), 
        .Q(\DP/ALU0/S_B_ADDER[22] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[23]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N77 ), 
        .Q(\DP/ALU0/S_B_ADDER[23] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[24]  ( .G(n2457), .D(\DP/ALU0/N78 ), .Q(
        \DP/ALU0/S_B_ADDER[24] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[25]  ( .G(n2457), .D(\DP/ALU0/N79 ), .Q(
        \DP/ALU0/S_B_ADDER[25] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[27]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N81 ), 
        .Q(\DP/ALU0/S_B_ADDER[27] ) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[26]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N80 ), 
        .Q(\DP/ALU0/S_B_ADDER[26] ) );
  DLL_X1 \DP/ALU0/s_A_SHIFT_reg[10]  ( .D(\DP/A[10] ), .GN(n2444), .Q(
        \DP/ALU0/s_A_SHIFT[10] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[10]  ( .D(\DP/A[10] ), .GN(n2446), .Q(
        \DP/ALU0/s_A_LOGIC[10] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[10]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N32 ), 
        .Q(\DP/ALU0/s_A_ADDER[10] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[10]  ( .D(\DP/RegNPC2/N13 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[10] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[10]  ( .D(\DP/RegNPC3/N13 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[10] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[13]  ( .D(\DP/A[13] ), .GN(n2447), .Q(
        \DP/ALU0/s_A_LOGIC[13] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[13]  ( .G(n2457), .D(\DP/ALU0/N35 ), .Q(
        \DP/ALU0/s_A_ADDER[13] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[13]  ( .D(\DP/RegNPC2/N16 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[13] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[13]  ( .D(\DP/RegNPC3/N16 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[13] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[16]  ( .D(n151), .GN(n2446), .Q(n9) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[16]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N38 ), 
        .Q(\DP/ALU0/s_A_ADDER[16] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[16]  ( .D(\DP/RegNPC2/N19 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[16] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[16]  ( .D(\DP/RegNPC3/N19 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[16] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[18]  ( .D(n145), .GN(n2447), .Q(n8) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[18]  ( .G(n2457), .D(\DP/ALU0/N40 ), .Q(
        \DP/ALU0/s_A_ADDER[18] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[18]  ( .D(\DP/RegNPC2/N21 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[18] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[18]  ( .D(\DP/RegNPC3/N21 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[18] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[17]  ( .D(\DP/RegNPC2/N20 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[17] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[17]  ( .D(\DP/RegNPC3/N20 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[17] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[20]  ( .D(n139), .GN(n2446), .Q(n7) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[20]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N42 ), 
        .Q(\DP/ALU0/s_A_ADDER[20] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[20]  ( .D(\DP/RegNPC2/N23 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[20] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[20]  ( .D(\DP/RegNPC3/N23 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[20] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[22]  ( .D(n133), .GN(n2447), .Q(n6) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[22]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N44 ), 
        .Q(\DP/ALU0/s_A_ADDER[22] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[22]  ( .D(\DP/RegNPC2/N25 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[22] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[22]  ( .D(\DP/RegNPC3/N25 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[22] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[21]  ( .D(\DP/RegNPC2/N24 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[21] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[21]  ( .D(\DP/RegNPC3/N24 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[21] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[24]  ( .D(n127), .GN(n2446), .Q(n5) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[24]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N46 ), 
        .Q(\DP/ALU0/s_A_ADDER[24] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[24]  ( .D(\DP/RegNPC2/N27 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[24] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[24]  ( .D(\DP/RegNPC3/N27 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[24] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[3]  ( .D(\DP/A[3] ), .GN(n2447), .Q(
        \DP/ALU0/s_A_LOGIC[3] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[3]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N25 ), 
        .Q(\DP/ALU0/s_A_ADDER[3] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[3]  ( .D(\DP/RegNPC2/N6 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[3] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[3]  ( .D(\DP/RegNPC3/N6 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[3] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[2]  ( .D(\DP/RegNPC2/N5 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[2] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[2]  ( .D(\DP/RegNPC3/N5 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[2] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[1]  ( .D(\DP/RegNPC2/N4 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[1] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[1]  ( .D(\DP/RegNPC3/N4 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[1] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[4]  ( .D(\DP/A[4] ), .GN(n2446), .Q(
        \DP/ALU0/s_A_LOGIC[4] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[4]  ( .G(\DP/ALU0/N21 ), .D(n189), .Q(
        \DP/ALU0/s_A_ADDER[4] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[4]  ( .D(\DP/RegNPC2/N7 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[4] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[4]  ( .D(\DP/RegNPC3/N7 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[4] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[7]  ( .D(\DP/A[7] ), .GN(n2447), .Q(
        \DP/ALU0/s_A_LOGIC[7] ) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[7]  ( .G(n2457), .D(\DP/ALU0/N29 ), .Q(
        \DP/ALU0/s_A_ADDER[7] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[7]  ( .D(\DP/RegNPC2/N10 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[7] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[7]  ( .D(\DP/RegNPC3/N10 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[7] ) );
  DFF_X1 \DP/RegA1/DOUT_reg[6]  ( .D(\DP/RegA1/N9 ), .CK(\DP/RegA1/net2366 ), 
        .Q(\DP/RegA1_out[6] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[25]  ( .D(n124), .GN(n2446), .Q(n4) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[25]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N47 ), 
        .Q(\DP/ALU0/s_A_ADDER[25] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[25]  ( .D(\DP/RegNPC2/N28 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[25] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[25]  ( .D(\DP/RegNPC3/N28 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[25] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[28]  ( .D(n115), .GN(n2447), .Q(n3) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[28]  ( .G(n2457), .D(\DP/ALU0/N50 ), .Q(
        \DP/ALU0/s_A_ADDER[28] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[28]  ( .D(\DP/RegNPC2/N31 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[28] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[28]  ( .D(\DP/RegNPC3/N31 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[28] ) );
  DLL_X1 \DP/ALU0/s_A_LOGIC_reg[30]  ( .D(n109), .GN(n2446), .Q(n2) );
  DLH_X1 \DP/ALU0/s_A_ADDER_reg[30]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N52 ), 
        .Q(\DP/ALU0/s_A_ADDER[30] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[30]  ( .D(\DP/RegNPC2/N33 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[30] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[30]  ( .D(\DP/RegNPC3/N33 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[30] ) );
  DFF_X1 \DP/RegALU1/DOUT_reg[31]  ( .D(\DP/RegALU1/N34 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[31] ) );
  DFF_X1 \DP/RegALU2/DOUT_reg[31]  ( .D(\DP/RegALU2/N34 ), .CK(n2454), .Q(
        \DP/RegALU2_out[31] ) );
  DLL_X1 \DP/ALU0/S_B_LOGIC_reg[31]  ( .D(n107), .GN(n2447), .Q(n1) );
  DLH_X1 \DP/ALU0/S_B_ADDER_reg[31]  ( .G(\DP/ALU0/N21 ), .D(\DP/ALU0/N85 ), 
        .Q(\DP/ALU0/S_B_ADDER[31] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[29]  ( .D(\DP/RegNPC2/N32 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[29] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[29]  ( .D(\DP/RegNPC3/N32 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[29] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[27]  ( .D(\DP/RegNPC2/N30 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[27] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[27]  ( .D(\DP/RegNPC3/N30 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[27] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[26]  ( .D(\DP/RegNPC2/N29 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[26] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[26]  ( .D(\DP/RegNPC3/N29 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[26] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[23]  ( .D(\DP/RegNPC2/N26 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[23] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[23]  ( .D(\DP/RegNPC3/N26 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[23] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[19]  ( .D(\DP/RegNPC2/N22 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[19] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[19]  ( .D(\DP/RegNPC3/N22 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[19] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[15]  ( .D(\DP/RegNPC2/N18 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[15] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[15]  ( .D(\DP/RegNPC3/N18 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[15] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[14]  ( .D(\DP/RegNPC2/N17 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[14] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[14]  ( .D(\DP/RegNPC3/N17 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[14] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[11]  ( .D(\DP/RegNPC2/N14 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[11] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[11]  ( .D(\DP/RegNPC3/N14 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[11] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[9]  ( .D(\DP/RegNPC2/N12 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[9] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[9]  ( .D(\DP/RegNPC3/N12 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[9] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[8]  ( .D(\DP/RegNPC2/N11 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[8] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[8]  ( .D(\DP/RegNPC3/N11 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[8] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[5]  ( .D(\DP/RegNPC2/N8 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[5] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[5]  ( .D(\DP/RegNPC3/N8 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[5] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[0]  ( .D(\DP/RegNPC2/N3 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[0] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[0]  ( .D(\DP/RegNPC3/N3 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[0] ) );
  DFF_X1 \DP/RegNPC2/DOUT_reg[31]  ( .D(\DP/RegNPC2/N34 ), .CK(
        \DP/RegNPC2/net2366 ), .Q(\DP/NPC3[31] ) );
  DFF_X1 \DP/RegNPC3/DOUT_reg[31]  ( .D(\DP/RegNPC3/N34 ), .CK(
        \DP/RegNPC3/net2366 ), .Q(\DP/NPC_out[31] ) );
  NOR2_X1 U3059 ( .A1(n3893), .A2(n3889), .ZN(n2343) );
  NOR2_X1 U3060 ( .A1(n3892), .A2(n2343), .ZN(n2344) );
  AOI21_X1 U3061 ( .B1(n3888), .B2(\DP/ALU0/s_A_ADDER[19] ), .A(n2344), .ZN(
        n3904) );
  NAND2_X1 U3062 ( .A1(n3904), .A2(n3954), .ZN(n2345) );
  XNOR2_X1 U3063 ( .A(n2345), .B(n3953), .ZN(n3997) );
  OAI22_X1 U3064 ( .A1(n4555), .A2(n4525), .B1(n2506), .B2(n2507), .ZN(n2346)
         );
  AOI211_X1 U3066 ( .C1(IR_OUT[1]), .C2(n2347), .A(n2512), .B(n2364), .ZN(
        n2348) );
  INV_X1 U3067 ( .A(IR_OUT[1]), .ZN(n2349) );
  AOI21_X1 U3069 ( .B1(n2543), .B2(n2560), .A(IR_OUT[0]), .ZN(n2351) );
  AOI211_X1 U3070 ( .C1(n2348), .C2(n2350), .A(n2555), .B(n2351), .ZN(n2352)
         );
  OAI211_X1 U3072 ( .C1(n2574), .C2(n2549), .A(n2511), .B(n2510), .ZN(n2354)
         );
  NOR2_X1 U3074 ( .A1(n2461), .A2(n2355), .ZN(\CU/N75 ) );
  OR3_X1 U3075 ( .A1(\DP/ALU0/S_B_MULT[1] ), .A2(\DP/ALU0/S_B_MULT[2] ), .A3(
        n2599), .ZN(n2356) );
  OR3_X1 U3076 ( .A1(n29), .A2(n2984), .A3(n3154), .ZN(n2357) );
  INV_X1 U3077 ( .A(n2357), .ZN(n2358) );
  INV_X1 U3078 ( .A(n2356), .ZN(n2359) );
  AOI21_X2 U3079 ( .B1(\DP/ALU0/s_A_MULT[3] ), .B2(n2606), .A(n2605), .ZN(
        n2912) );
  AOI21_X2 U3080 ( .B1(\DP/ALU0/s_A_MULT[4] ), .B2(n2615), .A(n2621), .ZN(
        n2955) );
  NOR2_X2 U3081 ( .A1(n2984), .A2(n3034), .ZN(n3078) );
  NOR2_X2 U3082 ( .A1(\DP/ALU0/S_B_MULT[5] ), .A2(n2622), .ZN(n3037) );
  NOR2_X2 U3083 ( .A1(n2810), .A2(n12), .ZN(n3304) );
  NOR2_X2 U3084 ( .A1(n3811), .A2(n3810), .ZN(n2340) );
  NOR3_X4 U3085 ( .A1(n31), .A2(n2652), .A3(n2650), .ZN(n3118) );
  NOR3_X4 U3086 ( .A1(n29), .A2(n54), .A3(n2691), .ZN(n3177) );
  AOI21_X2 U3087 ( .B1(n2637), .B2(n3032), .A(n2657), .ZN(n3029) );
  AOI21_X2 U3088 ( .B1(n2683), .B2(n3126), .A(n2705), .ZN(n3127) );
  NOR2_X2 U3089 ( .A1(\DP/ALU0/S_B_MULT[3] ), .A2(n2600), .ZN(n2962) );
  AOI21_X2 U3090 ( .B1(\DP/ALU0/s_A_MULT[10] ), .B2(n2735), .A(n2749), .ZN(
        n3222) );
  AOI21_X2 U3091 ( .B1(\DP/ALU0/s_A_MULT[12] ), .B2(n2777), .A(n2828), .ZN(
        n3276) );
  AOI21_X2 U3092 ( .B1(n2843), .B2(n3309), .A(n2922), .ZN(n3368) );
  NOR4_X4 U3094 ( .A1(w_LOAD_SIZE[1]), .A2(n202), .A3(w_LOAD_SIZE[2]), .A4(
        n2461), .ZN(n4306) );
  INV_X1 U3095 ( .A(n4623), .ZN(n2447) );
  INV_X1 U3096 ( .A(n2445), .ZN(n2444) );
  BUF_X1 U3097 ( .A(\DP/ALU0/N21 ), .Z(n2457) );
  AND2_X1 U3098 ( .A1(RST), .A2(\DP/RegALU1_out[25] ), .ZN(\DP/RegALU2/N28 )
         );
  AND2_X1 U3099 ( .A1(RST), .A2(\DP/RegALU1_out[17] ), .ZN(\DP/RegALU2/N20 )
         );
  AND2_X1 U3100 ( .A1(RST), .A2(\DP/RegALU1_out[12] ), .ZN(\DP/RegALU2/N15 )
         );
  AND2_X1 U3101 ( .A1(RST), .A2(DRAM_ADDR[10]), .ZN(\DP/RegALU2/N13 ) );
  AND2_X1 U3102 ( .A1(RST), .A2(\DP/RegALU1_out[13] ), .ZN(\DP/RegALU2/N16 )
         );
  AND2_X1 U3103 ( .A1(RST), .A2(DRAM_ADDR[7]), .ZN(\DP/RegALU2/N10 ) );
  AND2_X1 U3104 ( .A1(RST), .A2(DRAM_ADDR[4]), .ZN(\DP/RegALU2/N7 ) );
  AND2_X1 U3105 ( .A1(RST), .A2(DRAM_ADDR[1]), .ZN(\DP/RegALU2/N4 ) );
  AND2_X1 U3106 ( .A1(RST), .A2(DRAM_ADDR[2]), .ZN(\DP/RegALU2/N5 ) );
  AND2_X1 U3107 ( .A1(RST), .A2(DRAM_ADDR[3]), .ZN(\DP/RegALU2/N6 ) );
  AND2_X1 U3108 ( .A1(RST), .A2(\DP/RegALU1_out[21] ), .ZN(\DP/RegALU2/N24 )
         );
  AND2_X1 U3109 ( .A1(RST), .A2(\DP/RegALU1_out[22] ), .ZN(\DP/RegALU2/N25 )
         );
  AND2_X1 U3110 ( .A1(RST), .A2(\DP/RegALU1_out[20] ), .ZN(\DP/RegALU2/N23 )
         );
  AND2_X1 U3111 ( .A1(RST), .A2(\DP/RegALU1_out[16] ), .ZN(\DP/RegALU2/N19 )
         );
  AND2_X1 U3112 ( .A1(RST), .A2(IROM_DATA[31]), .ZN(\IR/N34 ) );
  AND2_X1 U3113 ( .A1(RST), .A2(IROM_DATA[30]), .ZN(\IR/N33 ) );
  AND2_X1 U3114 ( .A1(RST), .A2(IROM_DATA[29]), .ZN(\IR/N32 ) );
  AND2_X1 U3115 ( .A1(RST), .A2(IROM_DATA[28]), .ZN(\IR/N31 ) );
  AND2_X1 U3116 ( .A1(RST), .A2(IROM_DATA[27]), .ZN(\IR/N30 ) );
  AND2_X1 U3117 ( .A1(RST), .A2(IROM_DATA[26]), .ZN(\IR/N29 ) );
  AND2_X1 U3118 ( .A1(RST), .A2(IROM_DATA[25]), .ZN(\IR/N28 ) );
  AND2_X1 U3119 ( .A1(RST), .A2(IROM_DATA[24]), .ZN(\IR/N27 ) );
  AND2_X1 U3120 ( .A1(RST), .A2(IROM_DATA[23]), .ZN(\IR/N26 ) );
  AND2_X1 U3121 ( .A1(RST), .A2(IROM_DATA[22]), .ZN(\IR/N25 ) );
  AND2_X1 U3122 ( .A1(RST), .A2(IROM_DATA[21]), .ZN(\IR/N24 ) );
  AND2_X1 U3123 ( .A1(RST), .A2(IROM_DATA[20]), .ZN(\IR/N23 ) );
  AND2_X1 U3124 ( .A1(RST), .A2(IROM_DATA[19]), .ZN(\IR/N22 ) );
  AND2_X1 U3125 ( .A1(RST), .A2(IROM_DATA[18]), .ZN(\IR/N21 ) );
  AND2_X1 U3126 ( .A1(RST), .A2(IROM_DATA[17]), .ZN(\IR/N20 ) );
  AND2_X1 U3127 ( .A1(RST), .A2(IROM_DATA[16]), .ZN(\IR/N19 ) );
  AND2_X1 U3128 ( .A1(RST), .A2(IROM_DATA[15]), .ZN(\IR/N18 ) );
  AND2_X1 U3129 ( .A1(RST), .A2(IROM_DATA[14]), .ZN(\IR/N17 ) );
  AND2_X1 U3130 ( .A1(RST), .A2(IROM_DATA[13]), .ZN(\IR/N16 ) );
  AND2_X1 U3131 ( .A1(RST), .A2(IROM_DATA[12]), .ZN(\IR/N15 ) );
  AND2_X1 U3132 ( .A1(RST), .A2(IROM_DATA[11]), .ZN(\IR/N14 ) );
  AND2_X1 U3133 ( .A1(RST), .A2(IROM_DATA[10]), .ZN(\IR/N13 ) );
  AND2_X1 U3134 ( .A1(RST), .A2(IROM_DATA[9]), .ZN(\IR/N12 ) );
  AND2_X1 U3135 ( .A1(RST), .A2(IROM_DATA[8]), .ZN(\IR/N11 ) );
  AND2_X1 U3136 ( .A1(RST), .A2(IROM_DATA[7]), .ZN(\IR/N10 ) );
  AND2_X1 U3137 ( .A1(RST), .A2(IROM_DATA[6]), .ZN(\IR/N9 ) );
  AND2_X1 U3138 ( .A1(RST), .A2(IROM_DATA[5]), .ZN(\IR/N8 ) );
  AND2_X1 U3139 ( .A1(RST), .A2(IROM_DATA[4]), .ZN(\IR/N7 ) );
  AND2_X1 U3140 ( .A1(RST), .A2(IROM_DATA[3]), .ZN(\IR/N6 ) );
  AND2_X1 U3141 ( .A1(RST), .A2(IROM_DATA[2]), .ZN(\IR/N5 ) );
  AND2_X1 U3142 ( .A1(RST), .A2(IROM_DATA[1]), .ZN(\IR/N4 ) );
  AND2_X1 U3143 ( .A1(RST), .A2(IROM_DATA[0]), .ZN(\IR/N3 ) );
  NOR2_X1 U3144 ( .A1(n4306), .A2(n4287), .ZN(n4286) );
  NAND2_X1 U3145 ( .A1(n4289), .A2(n4288), .ZN(n4305) );
  NAND3_X1 U3146 ( .A1(n4277), .A2(\DP/LOAD8[7] ), .A3(w_SIGN_LD), .ZN(n4288)
         );
  INV_X1 U3147 ( .A(RST), .ZN(n2460) );
  AND2_X1 U3148 ( .A1(RST), .A2(\DP/RegALU1_out[18] ), .ZN(\DP/RegALU2/N21 )
         );
  AND2_X1 U3149 ( .A1(RST), .A2(DRAM_ADDR[6]), .ZN(\DP/RegALU2/N9 ) );
  AND2_X1 U3150 ( .A1(RST), .A2(\DP/RegALU1_out[14] ), .ZN(\DP/RegALU2/N17 )
         );
  AND2_X1 U3151 ( .A1(RST), .A2(\DP/RegALU1_out[15] ), .ZN(\DP/RegALU2/N18 )
         );
  AND2_X1 U3152 ( .A1(RST), .A2(\DP/RegALU1_out[19] ), .ZN(\DP/RegALU2/N22 )
         );
  BUF_X1 U3153 ( .A(n4515), .Z(n2442) );
  AND2_X1 U3155 ( .A1(RST), .A2(\DP/RegALU1_out[26] ), .ZN(\DP/RegALU2/N29 )
         );
  AND2_X1 U3156 ( .A1(RST), .A2(\DP/RegALU1_out[27] ), .ZN(\DP/RegALU2/N30 )
         );
  AND2_X1 U3157 ( .A1(n12), .A2(n2808), .ZN(n3310) );
  INV_X1 U3158 ( .A(n2760), .ZN(n3236) );
  AND2_X1 U3159 ( .A1(n2872), .A2(n3298), .ZN(n3270) );
  AND2_X1 U3160 ( .A1(RST), .A2(\DP/RegALU1_out[29] ), .ZN(\DP/RegALU2/N32 )
         );
  INV_X1 U3161 ( .A(n2441), .ZN(n2439) );
  INV_X1 U3162 ( .A(n3248), .ZN(n3364) );
  INV_X1 U3163 ( .A(n3345), .ZN(n3392) );
  AND2_X1 U3164 ( .A1(RST), .A2(\DP/RegALU1_out[30] ), .ZN(\DP/RegALU2/N33 )
         );
  AND2_X1 U3165 ( .A1(RST), .A2(n2340), .ZN(n4164) );
  BUF_X1 U3166 ( .A(n3690), .Z(n2420) );
  AND2_X1 U3167 ( .A1(\DP/RegALU1_out[31] ), .A2(RST), .ZN(\DP/RegALU2/N34 )
         );
  NAND3_X1 U3179 ( .A1(RST), .A2(n2508), .A3(n2502), .ZN(n4273) );
  AND2_X1 U3185 ( .A1(RST), .A2(DRAM_ADDR[0]), .ZN(\DP/RegALU2/N3 ) );
  INV_X1 U3186 ( .A(n2386), .ZN(n2408) );
  INV_X1 U3187 ( .A(n2383), .ZN(n2412) );
  INV_X1 U3188 ( .A(n4223), .ZN(n2427) );
  INV_X1 U3189 ( .A(n2389), .ZN(n2430) );
  AND2_X1 U3192 ( .A1(RST), .A2(DRAM_ADDR[5]), .ZN(\DP/RegALU2/N8 ) );
  BUF_X1 U3193 ( .A(n4515), .Z(n2443) );
  BUF_X1 U3195 ( .A(n3691), .Z(n2422) );
  INV_X1 U3196 ( .A(n2381), .ZN(n2438) );
  AND2_X1 U3197 ( .A1(RST), .A2(DRAM_ADDR[8]), .ZN(\DP/RegALU2/N11 ) );
  INV_X1 U3198 ( .A(n2361), .ZN(n2416) );
  INV_X1 U3199 ( .A(n2384), .ZN(n2417) );
  INV_X1 U3201 ( .A(n4267), .ZN(n100) );
  INV_X1 U3202 ( .A(n4270), .ZN(n103) );
  INV_X1 U3203 ( .A(n4272), .ZN(n104) );
  INV_X1 U3204 ( .A(n4269), .ZN(n102) );
  INV_X1 U3205 ( .A(n4268), .ZN(n101) );
  AND2_X1 U3206 ( .A1(RST), .A2(\DP/RegALU1_out[28] ), .ZN(\DP/RegALU2/N31 )
         );
  INV_X1 U3208 ( .A(n4498), .ZN(n2441) );
  INV_X1 U3209 ( .A(n2952), .ZN(n2876) );
  INV_X1 U3210 ( .A(n3076), .ZN(n2963) );
  INV_X1 U3211 ( .A(n2623), .ZN(n3033) );
  INV_X1 U3212 ( .A(n2604), .ZN(n2926) );
  AND3_X1 U3213 ( .A1(n2872), .A2(\DP/ALU0/S_B_MULT[1] ), .A3(
        \DP/ALU0/S_B_MULT[0] ), .ZN(n2886) );
  OR2_X1 U3214 ( .A1(\DP/ALU0/S_B_MULT[3] ), .A2(n2601), .ZN(n2960) );
  INV_X1 U3215 ( .A(n49), .ZN(n3309) );
  INV_X1 U3216 ( .A(n53), .ZN(n3126) );
  INV_X1 U3217 ( .A(n30), .ZN(n3032) );
  INV_X1 U3218 ( .A(\DP/ALU0/s_A_MULT[2] ), .ZN(n2951) );
  INV_X1 U3219 ( .A(\DP/ALU0/s_A_MULT[9] ), .ZN(n3220) );
  INV_X1 U3220 ( .A(\DP/ALU0/s_A_MULT[11] ), .ZN(n3274) );
  INV_X1 U3221 ( .A(\DP/ALU0/s_A_MULT[13] ), .ZN(n3350) );
  INV_X1 U3222 ( .A(n3420), .ZN(n4515) );
  OAI21_X1 U3223 ( .B1(n2586), .B2(w_ALU_OPCODE[3]), .A(n1272), .ZN(n3420) );
  NOR2_X1 U3224 ( .A1(n3695), .A2(\DP/ALU0/N91 ), .ZN(n1272) );
  AND2_X1 U3225 ( .A1(RST), .A2(DRAM_ADDR[11]), .ZN(\DP/RegALU2/N14 ) );
  INV_X1 U3227 ( .A(n4205), .ZN(n2425) );
  BUF_X1 U3228 ( .A(n4223), .Z(n2429) );
  BUF_X1 U3229 ( .A(n4413), .Z(n2435) );
  AND3_X1 U3230 ( .A1(RST), .A2(\DP/OUTCOME ), .A3(\DP/JREG ), .ZN(n4413) );
  BUF_X1 U3231 ( .A(n4414), .Z(n2436) );
  NOR2_X1 U3232 ( .A1(\DP/JREG ), .A2(n2405), .ZN(n4414) );
  INV_X1 U3233 ( .A(n2381), .ZN(n2437) );
  OR2_X1 U3234 ( .A1(n2460), .A2(\DP/OUTCOME ), .ZN(n2381) );
  BUF_X1 U3239 ( .A(n3386), .Z(n2410) );
  INV_X1 U3243 ( .A(n2426), .ZN(n2424) );
  INV_X1 U3244 ( .A(n4090), .ZN(n4083) );
  INV_X1 U3245 ( .A(n4171), .ZN(n4152) );
  BUF_X1 U3246 ( .A(n4205), .Z(n2426) );
  INV_X1 U3247 ( .A(n4223), .ZN(n2428) );
  XNOR2_X1 U3248 ( .A(n3819), .B(\DP/ALU0/S_B_SHIFT[1] ), .ZN(n4223) );
  INV_X1 U3249 ( .A(n2396), .ZN(n2432) );
  INV_X1 U3251 ( .A(n4096), .ZN(n4098) );
  NOR2_X1 U3252 ( .A1(\DP/ALU0/s_SHIFT[0] ), .A2(\DP/ALU0/s_SHIFT[1] ), .ZN(
        n3819) );
  INV_X1 U3254 ( .A(n4178), .ZN(n4231) );
  INV_X1 U3255 ( .A(n2389), .ZN(n2431) );
  OR2_X1 U3256 ( .A1(n4101), .A2(n2461), .ZN(n2389) );
  NOR3_X1 U3257 ( .A1(n3576), .A2(n2373), .A3(w_ALU_OPCODE[2]), .ZN(n3696) );
  BUF_X1 U3258 ( .A(n57), .Z(n2450) );
  BUF_X1 U3263 ( .A(n3387), .Z(n2411) );
  NOR2_X1 U3264 ( .A1(n2583), .A2(n2406), .ZN(n3387) );
  INV_X1 U3265 ( .A(n2386), .ZN(n2409) );
  NOR2_X1 U3266 ( .A1(w_MuxA_SEL), .A2(n2583), .ZN(n3386) );
  INV_X1 U3267 ( .A(n2383), .ZN(n2413) );
  AND3_X1 U3268 ( .A1(n407), .A2(n406), .A3(\DP/FwdC[1] ), .ZN(n2383) );
  BUF_X1 U3269 ( .A(n3569), .Z(n2419) );
  NOR2_X1 U3270 ( .A1(n3407), .A2(n2407), .ZN(n3569) );
  BUF_X1 U3271 ( .A(n3566), .Z(n2414) );
  NOR2_X1 U3272 ( .A1(w_MuxB_SEL), .A2(n3407), .ZN(n3566) );
  INV_X1 U3273 ( .A(n2361), .ZN(n2415) );
  OR3_X1 U3274 ( .A1(n405), .A2(\DP/FwdB[1] ), .A3(n2368), .ZN(n2361) );
  INV_X1 U3275 ( .A(n2384), .ZN(n2418) );
  AND3_X1 U3276 ( .A1(n405), .A2(n404), .A3(\DP/FwdB[1] ), .ZN(n2384) );
  INV_X1 U3277 ( .A(n4765), .ZN(n98) );
  OR2_X1 U3278 ( .A1(n2459), .A2(\DP/RD3[0] ), .ZN(\DP/RF_ADDR[0] ) );
  INV_X1 U3279 ( .A(n4421), .ZN(n94) );
  OR2_X1 U3280 ( .A1(n2459), .A2(\DP/RD3[2] ), .ZN(\DP/RF_ADDR[2] ) );
  OR2_X1 U3282 ( .A1(n2459), .A2(\DP/RD3[1] ), .ZN(\DP/RF_ADDR[1] ) );
  OR2_X1 U3284 ( .A1(n2459), .A2(\DP/RD3[3] ), .ZN(\DP/RF_ADDR[3] ) );
  INV_X1 U3285 ( .A(n4424), .ZN(n97) );
  OR2_X1 U3286 ( .A1(n2459), .A2(\DP/RD3[4] ), .ZN(\DP/RF_ADDR[4] ) );
  AND2_X1 U3288 ( .A1(RST), .A2(DRAM_ADDR[9]), .ZN(\DP/RegALU2/N12 ) );
  BUF_X1 U3289 ( .A(n3690), .Z(n2421) );
  AND2_X1 U3290 ( .A1(RST), .A2(n3655), .ZN(n3691) );
  BUF_X1 U3291 ( .A(n3693), .Z(n2423) );
  OR2_X1 U3292 ( .A1(n2461), .A2(n3654), .ZN(n3693) );
  INV_X1 U3293 ( .A(RST), .ZN(n2461) );
  BUF_X1 U3294 ( .A(\DP/RegLMD/net2366 ), .Z(n2455) );
  BUF_X1 U3295 ( .A(\DP/RegLMD/net2366 ), .Z(n2454) );
  BUF_X1 U3296 ( .A(\DP/RegLMD/net2366 ), .Z(n2453) );
  BUF_X1 U3297 ( .A(\DP/RegLMD/net2366 ), .Z(n2452) );
  BUF_X1 U3298 ( .A(\DP/RegNPC/net2366 ), .Z(n2456) );
  NAND2_X1 U3299 ( .A1(n204), .A2(DRAM_DATA_OUT[15]), .ZN(n4473) );
  AND2_X1 U3301 ( .A1(n205), .A2(n4482), .ZN(n4472) );
  NOR2_X1 U3302 ( .A1(\DP/FwdD ), .A2(n4489), .ZN(n4482) );
  INV_X1 U3303 ( .A(n4458), .ZN(n4475) );
  NOR2_X1 U3304 ( .A1(n2399), .A2(n4484), .ZN(n4458) );
  NAND2_X1 U3305 ( .A1(\DP/FwdD ), .A2(n4427), .ZN(n4484) );
  NOR2_X2 U3307 ( .A1(\DP/ALU0/S_B_MULT[1] ), .A2(n2591), .ZN(n2924) );
  INV_X1 U3308 ( .A(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .ZN(n2451) );
  OR3_X1 U3310 ( .A1(n407), .A2(\DP/FwdC[1] ), .A3(n2370), .ZN(n2386) );
  INV_X1 U3311 ( .A(n4498), .ZN(n2440) );
  NOR2_X1 U3317 ( .A1(n2467), .A2(IR_OUT[31]), .ZN(n2547) );
  NAND2_X1 U3320 ( .A1(n2527), .A2(n2528), .ZN(n2505) );
  INV_X1 U3322 ( .A(n2487), .ZN(n2488) );
  NOR2_X1 U3324 ( .A1(n2488), .A2(n4527), .ZN(n2497) );
  INV_X1 U3325 ( .A(n2497), .ZN(n2494) );
  NAND2_X1 U3326 ( .A1(n2505), .A2(n2494), .ZN(n2490) );
  NOR2_X1 U3327 ( .A1(IR_OUT[30]), .A2(n2479), .ZN(n2481) );
  NAND2_X1 U3328 ( .A1(n2481), .A2(n2547), .ZN(n2531) );
  INV_X1 U3329 ( .A(n2531), .ZN(n2464) );
  AOI211_X1 U3331 ( .C1(n2479), .C2(IR_OUT[27]), .A(n2371), .B(n2462), .ZN(
        n2463) );
  AOI211_X1 U3332 ( .C1(n224), .C2(n2464), .A(n2463), .B(n2516), .ZN(n2500) );
  NOR2_X1 U3333 ( .A1(n2397), .A2(n2467), .ZN(n2480) );
  INV_X1 U3334 ( .A(n2480), .ZN(n2466) );
  NAND2_X1 U3336 ( .A1(n2471), .A2(n4566), .ZN(n2569) );
  NAND2_X1 U3342 ( .A1(n2526), .A2(n2467), .ZN(n2469) );
  INV_X1 U3348 ( .A(n2469), .ZN(n2491) );
  INV_X1 U3350 ( .A(n2574), .ZN(n2483) );
  INV_X1 U3351 ( .A(n2528), .ZN(n2507) );
  AOI21_X1 U3352 ( .B1(n2506), .B2(n2483), .A(n2507), .ZN(n2470) );
  NAND2_X1 U3355 ( .A1(n2527), .A2(n2491), .ZN(n2566) );
  NOR2_X1 U3359 ( .A1(n2490), .A2(n2486), .ZN(n2476) );
  NOR4_X1 U3360 ( .A1(IR_OUT[8]), .A2(IR_OUT[7]), .A3(IR_OUT[6]), .A4(
        IR_OUT[10]), .ZN(n2473) );
  NAND2_X1 U3361 ( .A1(n2473), .A2(n2391), .ZN(n2513) );
  NOR2_X1 U3362 ( .A1(IR_OUT[1]), .A2(IR_OUT[0]), .ZN(n2535) );
  NOR2_X1 U3363 ( .A1(IR_OUT[4]), .A2(IR_OUT[3]), .ZN(n2520) );
  NAND4_X1 U3364 ( .A1(n2535), .A2(n2520), .A3(n2364), .A4(n2377), .ZN(n2475)
         );
  AOI21_X1 U3368 ( .B1(n2476), .B2(n2485), .A(n2460), .ZN(\CU/N40 ) );
  NAND2_X1 U3369 ( .A1(RST), .A2(n2525), .ZN(n2499) );
  NOR2_X1 U3370 ( .A1(n2478), .A2(n2499), .ZN(\CU/N43 ) );
  NOR3_X1 U3371 ( .A1(n2460), .A2(n2478), .A3(n4553), .ZN(\CU/N42 ) );
  NOR3_X1 U3372 ( .A1(n2460), .A2(n2478), .A3(n4527), .ZN(\CU/N41 ) );
  AND2_X1 U3373 ( .A1(n2516), .A2(RST), .ZN(\CU/N39 ) );
  NOR4_X1 U3374 ( .A1(n4559), .A2(n2460), .A3(n2479), .A4(n2478), .ZN(\CU/N44 ) );
  NAND2_X1 U3375 ( .A1(n2481), .A2(n2480), .ZN(n2484) );
  INV_X1 U3376 ( .A(n2484), .ZN(n2482) );
  NAND2_X1 U3377 ( .A1(n2482), .A2(n2506), .ZN(n2511) );
  NOR2_X1 U3378 ( .A1(n2461), .A2(n2511), .ZN(\CU/N48 ) );
  AND2_X1 U3379 ( .A1(n4559), .A2(\CU/N48 ), .ZN(\CU/N45 ) );
  NOR3_X1 U3380 ( .A1(n2460), .A2(n2484), .A3(n4553), .ZN(\CU/N46 ) );
  NOR2_X1 U3381 ( .A1(n2484), .A2(n2499), .ZN(\CU/N47 ) );
  NAND2_X1 U3384 ( .A1(n2487), .A2(n2509), .ZN(n2495) );
  INV_X1 U3386 ( .A(n2501), .ZN(n2489) );
  OAI21_X1 U3387 ( .B1(n2506), .B2(n2495), .A(n2489), .ZN(n2496) );
  NOR3_X1 U3388 ( .A1(n2491), .A2(n2496), .A3(n2490), .ZN(n2493) );
  NOR2_X1 U3389 ( .A1(n2372), .A2(n4273), .ZN(\CU/N53 ) );
  INV_X1 U3390 ( .A(\CU/N53 ), .ZN(n2492) );
  OAI221_X1 U3391 ( .B1(n2460), .B2(n4533), .C1(n2461), .C2(n2493), .A(n2492), 
        .ZN(\CU/N49 ) );
  NOR2_X1 U3392 ( .A1(n2460), .A2(n2494), .ZN(\CU/N50 ) );
  NOR3_X1 U3393 ( .A1(n2461), .A2(n4566), .A3(n2495), .ZN(\CU/N51 ) );
  NOR2_X1 U3397 ( .A1(n2515), .A2(n2499), .ZN(\CU/N52 ) );
  NAND3_X1 U3398 ( .A1(n2500), .A2(n2511), .A3(n2505), .ZN(n4266) );
  AOI211_X1 U3399 ( .C1(n2502), .C2(n4555), .A(n2501), .B(n4266), .ZN(n2503)
         );
  AOI21_X1 U3400 ( .B1(n2504), .B2(n2503), .A(n2461), .ZN(\CU/N54 ) );
  NOR2_X1 U3401 ( .A1(n2461), .A2(n4533), .ZN(\CU/N55 ) );
  NOR2_X1 U3403 ( .A1(n2460), .A2(n4524), .ZN(\CU/N56 ) );
  AND2_X1 U3404 ( .A1(RST), .A2(w_RF_WE_EX), .ZN(\CU/N57 ) );
  AND2_X1 U3405 ( .A1(RST), .A2(\CU/cw1[1] ), .ZN(\CU/N58 ) );
  AND2_X1 U3406 ( .A1(RST), .A2(\CU/cw1[2] ), .ZN(\CU/N59 ) );
  AND2_X1 U3407 ( .A1(RST), .A2(\CU/cw1[3] ), .ZN(\CU/N60 ) );
  AND2_X1 U3408 ( .A1(RST), .A2(\CU/cw1[4] ), .ZN(\CU/N61 ) );
  AND2_X1 U3409 ( .A1(RST), .A2(\CU/cw1[5] ), .ZN(\CU/N62 ) );
  AND2_X1 U3410 ( .A1(RST), .A2(\CU/cw1[6] ), .ZN(\CU/N63 ) );
  AND2_X1 U3411 ( .A1(RST), .A2(\CU/cw1[7] ), .ZN(\CU/N64 ) );
  AND2_X1 U3412 ( .A1(RST), .A2(\CU/cw1[8] ), .ZN(\CU/N65 ) );
  AND2_X1 U3413 ( .A1(RST), .A2(\CU/cw1[9] ), .ZN(\CU/N66 ) );
  AND2_X1 U3414 ( .A1(RST), .A2(\CU/cw1[10] ), .ZN(\CU/N67 ) );
  AND2_X1 U3415 ( .A1(RST), .A2(\CU/cw1[11] ), .ZN(\CU/N68 ) );
  NOR2_X1 U3416 ( .A1(n2460), .A2(n2395), .ZN(\CU/N69 ) );
  AND2_X1 U3417 ( .A1(RST), .A2(\CU/cw2[1] ), .ZN(\CU/N70 ) );
  AND2_X1 U3418 ( .A1(RST), .A2(\CU/cw2[2] ), .ZN(\CU/N71 ) );
  NOR2_X1 U3419 ( .A1(n2515), .A2(n2461), .ZN(\CU/N72 ) );
  AND2_X1 U3420 ( .A1(RST), .A2(n4535), .ZN(\CU/N73 ) );
  AND2_X1 U3421 ( .A1(n4532), .A2(RST), .ZN(\CU/N74 ) );
  NAND2_X1 U3422 ( .A1(n2547), .A2(n2509), .ZN(n2549) );
  INV_X1 U3425 ( .A(n2520), .ZN(n2523) );
  NOR2_X1 U3426 ( .A1(IR_OUT[1]), .A2(n2375), .ZN(n2568) );
  INV_X1 U3429 ( .A(n2512), .ZN(n2517) );
  NOR2_X1 U3431 ( .A1(n2568), .A2(n2571), .ZN(n2555) );
  NAND3_X1 U3432 ( .A1(n2520), .A2(IR_OUT[5]), .A3(n2512), .ZN(n2543) );
  NAND2_X1 U3433 ( .A1(n2512), .A2(n2364), .ZN(n2522) );
  OR3_X1 U3434 ( .A1(IR_OUT[4]), .A2(n2382), .A3(n2522), .ZN(n2560) );
  INV_X1 U3436 ( .A(n2576), .ZN(n2537) );
  AOI21_X1 U3437 ( .B1(IR_OUT[1]), .B2(n2375), .A(n2568), .ZN(n2544) );
  NOR2_X1 U3439 ( .A1(IR_OUT[1]), .A2(n2517), .ZN(n2557) );
  INV_X1 U3440 ( .A(n2539), .ZN(n2518) );
  OAI211_X1 U3441 ( .C1(n2519), .C2(n2557), .A(IR_OUT[4]), .B(n2518), .ZN(
        n2578) );
  AOI22_X1 U3442 ( .A1(n2520), .A2(n2519), .B1(n2535), .B2(n2556), .ZN(n2521)
         );
  OAI21_X1 U3443 ( .B1(n2544), .B2(n2578), .A(n2521), .ZN(n2524) );
  INV_X1 U3444 ( .A(n4275), .ZN(n4274) );
  NOR2_X1 U3445 ( .A1(n2364), .A2(n4274), .ZN(\DP/RegIMM/N8 ) );
  NOR2_X1 U3446 ( .A1(n2375), .A2(n4274), .ZN(\DP/RegIMM/N3 ) );
  NOR2_X1 U3448 ( .A1(n2377), .A2(n4274), .ZN(\DP/RegIMM/N5 ) );
  AOI222_X1 U3449 ( .A1(n2524), .A2(\DP/RegIMM/N8 ), .B1(\DP/RegIMM/N3 ), .B2(
        n2555), .C1(n2540), .C2(\DP/RegIMM/N5 ), .ZN(n2538) );
  NOR2_X1 U3450 ( .A1(n2537), .A2(n2543), .ZN(n2534) );
  INV_X1 U3451 ( .A(n2549), .ZN(n2575) );
  OAI21_X1 U3452 ( .B1(n2575), .B2(n2526), .A(n2525), .ZN(n2529) );
  OAI21_X1 U3453 ( .B1(n2575), .B2(n2528), .A(n2527), .ZN(n2562) );
  OAI211_X1 U3454 ( .C1(n4566), .C2(n4525), .A(n2529), .B(n2562), .ZN(n2532)
         );
  AOI211_X1 U3455 ( .C1(n2535), .C2(n2534), .A(n2533), .B(n2532), .ZN(n2536)
         );
  OAI22_X1 U3456 ( .A1(n2538), .A2(n2537), .B1(n2536), .B2(n2461), .ZN(
        \CU/N76 ) );
  NOR2_X1 U3457 ( .A1(IR_OUT[0]), .A2(n2539), .ZN(n2554) );
  OAI211_X1 U3458 ( .C1(n2556), .C2(n2554), .A(IR_OUT[5]), .B(n2557), .ZN(
        n2542) );
  OAI211_X1 U3460 ( .C1(n2544), .C2(n2543), .A(n2542), .B(n2541), .ZN(n2551)
         );
  NAND3_X1 U3462 ( .A1(n2547), .A2(n2546), .A3(n2388), .ZN(n2548) );
  OAI21_X1 U3463 ( .B1(n2372), .B2(n2549), .A(n2548), .ZN(n2564) );
  AOI211_X1 U3464 ( .C1(n2576), .C2(n2551), .A(n2550), .B(n2564), .ZN(n2552)
         );
  AOI21_X1 U3465 ( .B1(n2553), .B2(n2552), .A(n2461), .ZN(\CU/N77 ) );
  AOI21_X1 U3466 ( .B1(IR_OUT[0]), .B2(n2390), .A(n2554), .ZN(n2561) );
  INV_X1 U3467 ( .A(n2555), .ZN(n2559) );
  NAND3_X1 U3468 ( .A1(IR_OUT[5]), .A2(n2557), .A3(n2556), .ZN(n2558) );
  OAI211_X1 U3469 ( .C1(n2561), .C2(n2560), .A(n2559), .B(n2558), .ZN(n2565)
         );
  INV_X1 U3470 ( .A(n2562), .ZN(n2563) );
  AOI211_X1 U3471 ( .C1(n2576), .C2(n2565), .A(n2564), .B(n2563), .ZN(n2567)
         );
  AOI21_X1 U3472 ( .B1(n4529), .B2(n2567), .A(n2460), .ZN(\CU/N78 ) );
  NAND2_X1 U3473 ( .A1(n2568), .A2(n2576), .ZN(n2570) );
  OAI21_X1 U3474 ( .B1(n2571), .B2(n2570), .A(n2569), .ZN(n2572) );
  NAND2_X1 U3476 ( .A1(n2576), .A2(\DP/RegIMM/N8 ), .ZN(n2577) );
  OAI22_X1 U3477 ( .A1(n2579), .A2(n2461), .B1(n2578), .B2(n2577), .ZN(
        \CU/N79 ) );
  NAND2_X1 U3478 ( .A1(n2376), .A2(n2363), .ZN(n3576) );
  INV_X1 U3479 ( .A(n3576), .ZN(n2580) );
  NAND2_X1 U3480 ( .A1(w_ALU_OPCODE[3]), .A2(n2580), .ZN(n2581) );
  NOR3_X1 U3481 ( .A1(w_ALU_OPCODE[2]), .A2(n4744), .A3(n2581), .ZN(n4065) );
  NAND2_X1 U3482 ( .A1(w_ALU_OPCODE[2]), .A2(n4744), .ZN(n2582) );
  NAND3_X1 U3483 ( .A1(w_ALU_OPCODE[3]), .A2(n218), .A3(n2376), .ZN(n3810) );
  NOR2_X1 U3484 ( .A1(n2582), .A2(n3810), .ZN(n4068) );
  NOR3_X1 U3485 ( .A1(w_ALU_OPCODE[4]), .A2(n4744), .A3(n2362), .ZN(n4486) );
  NAND2_X1 U3486 ( .A1(w_ALU_OPCODE[3]), .A2(n4486), .ZN(n4059) );
  OAI22_X1 U3487 ( .A1(n2363), .A2(n4059), .B1(n2582), .B2(n2581), .ZN(n4104)
         );
  NOR3_X1 U3488 ( .A1(n4065), .A2(n4068), .A3(n4104), .ZN(n4522) );
  NAND4_X1 U3489 ( .A1(w_ALU_OPCODE[4]), .A2(n218), .A3(n4744), .A4(n2374), 
        .ZN(n4103) );
  NOR3_X1 U3490 ( .A1(n2376), .A2(w_ALU_OPCODE[3]), .A3(w_ALU_OPCODE[2]), .ZN(
        n4066) );
  INV_X1 U3491 ( .A(n4066), .ZN(n4067) );
  NAND4_X1 U3492 ( .A1(n4522), .A2(n4059), .A3(n4103), .A4(n4067), .ZN(
        \DP/ALU0/N91 ) );
  NAND2_X1 U3493 ( .A1(n2362), .A2(n2373), .ZN(n3811) );
  OR2_X1 U3494 ( .A1(n3811), .A2(w_ALU_OPCODE[3]), .ZN(n3575) );
  NOR3_X1 U3495 ( .A1(w_ALU_OPCODE[4]), .A2(n2363), .A3(n3575), .ZN(n3695) );
  NAND2_X1 U3496 ( .A1(w_ALU_OPCODE[3]), .A2(n3696), .ZN(n4498) );
  INV_X1 U3497 ( .A(n3696), .ZN(n2586) );
  NAND2_X1 U3498 ( .A1(n1272), .A2(n2586), .ZN(\DP/ALU0/N21 ) );
  AOI22_X1 U3499 ( .A1(n2449), .A2(\DP/RegALU2_out[0] ), .B1(
        \DP/RegLMD_out[0] ), .B2(n2360), .ZN(n4504) );
  NAND3_X1 U3500 ( .A1(n407), .A2(n2370), .A3(n2401), .ZN(n2583) );
  AOI22_X1 U3501 ( .A1(n3387), .A2(\DP/RegA_out[0] ), .B1(n2408), .B2(
        DRAM_ADDR[0]), .ZN(n2585) );
  NAND2_X1 U3502 ( .A1(n2410), .A2(\DP/NPC2[0] ), .ZN(n2584) );
  OAI211_X1 U3503 ( .C1(n4504), .C2(n2412), .A(n2585), .B(n2584), .ZN(
        \DP/A[0] ) );
  INV_X1 U3504 ( .A(\DP/A[0] ), .ZN(n2588) );
  INV_X1 U3505 ( .A(\DP/ALU0/S_B_MULT[0] ), .ZN(n2591) );
  NOR2_X1 U3506 ( .A1(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .A2(
        \DP/ALU0/s_A_MULT[1] ), .ZN(n2603) );
  NAND2_X1 U3507 ( .A1(n2603), .A2(n2951), .ZN(n2606) );
  NOR2_X1 U3508 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n2606), .ZN(n2605) );
  INV_X1 U3509 ( .A(n2605), .ZN(n2615) );
  NOR2_X1 U3510 ( .A1(n2615), .A2(\DP/ALU0/s_A_MULT[4] ), .ZN(n2621) );
  NAND2_X1 U3511 ( .A1(n2621), .A2(n55), .ZN(n2637) );
  NOR2_X1 U3512 ( .A1(n2637), .A2(n3032), .ZN(n2657) );
  NAND2_X1 U3513 ( .A1(n2657), .A2(n28), .ZN(n2683) );
  NOR2_X1 U3514 ( .A1(n2683), .A2(n3126), .ZN(n2705) );
  NAND2_X1 U3515 ( .A1(n3220), .A2(n2705), .ZN(n2735) );
  NOR2_X1 U3516 ( .A1(n2735), .A2(\DP/ALU0/s_A_MULT[10] ), .ZN(n2749) );
  NAND2_X1 U3517 ( .A1(n3274), .A2(n2749), .ZN(n2777) );
  NOR2_X1 U3518 ( .A1(n2777), .A2(\DP/ALU0/s_A_MULT[12] ), .ZN(n2828) );
  NAND2_X1 U3519 ( .A1(n3350), .A2(n2828), .ZN(n2843) );
  NOR2_X1 U3520 ( .A1(n2843), .A2(n3309), .ZN(n2922) );
  NAND2_X1 U3521 ( .A1(n2922), .A2(n47), .ZN(n2872) );
  NOR2_X1 U3522 ( .A1(n2924), .A2(n2886), .ZN(n2587) );
  NAND2_X1 U3523 ( .A1(n2441), .A2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .ZN(n2594)
         );
  OAI22_X1 U3524 ( .A1(n2443), .A2(n2588), .B1(n2587), .B2(n2594), .ZN(
        \DP/ALU0/N22 ) );
  AOI22_X1 U3525 ( .A1(n200), .A2(\DP/RegALU2_out[1] ), .B1(\DP/RegLMD_out[1] ), .B2(n2360), .ZN(n4502) );
  AOI22_X1 U3526 ( .A1(n2410), .A2(\DP/NPC2[1] ), .B1(n2409), .B2(DRAM_ADDR[1]), .ZN(n2590) );
  NAND2_X1 U3527 ( .A1(n2411), .A2(\DP/RegA_out[1] ), .ZN(n2589) );
  OAI211_X1 U3528 ( .C1(n4502), .C2(n2413), .A(n2590), .B(n2589), .ZN(
        \DP/A[1] ) );
  NAND3_X1 U3529 ( .A1(n2872), .A2(n2591), .A3(\DP/ALU0/S_B_MULT[1] ), .ZN(
        n2604) );
  INV_X1 U3530 ( .A(\DP/A[1] ), .ZN(n2593) );
  AOI21_X1 U3531 ( .B1(\DP/ALU0/s_A_MULT[1] ), .B2(
        \DP/ALU0/MULT/SHIFTERi_0/N19 ), .A(n2603), .ZN(n2874) );
  AOI22_X1 U3532 ( .A1(\DP/ALU0/s_A_MULT[1] ), .A2(n2924), .B1(n2874), .B2(
        n2886), .ZN(n2592) );
  OAI222_X1 U3533 ( .A1(n2594), .A2(n2604), .B1(n2443), .B2(n2593), .C1(n4498), 
        .C2(n2592), .ZN(\DP/ALU0/N23 ) );
  AOI22_X1 U3534 ( .A1(n2449), .A2(\DP/RegALU2_out[2] ), .B1(
        \DP/RegLMD_out[2] ), .B2(n2360), .ZN(n4494) );
  AOI22_X1 U3535 ( .A1(n3387), .A2(\DP/RegA_out[2] ), .B1(n2409), .B2(
        DRAM_ADDR[2]), .ZN(n2596) );
  NAND2_X1 U3536 ( .A1(n2410), .A2(\DP/NPC2[2] ), .ZN(n2595) );
  OAI211_X1 U3537 ( .C1(n4494), .C2(n2413), .A(n2596), .B(n2595), .ZN(
        \DP/A[2] ) );
  AOI22_X1 U3538 ( .A1(n200), .A2(\DP/RegALU2_out[3] ), .B1(\DP/RegLMD_out[3] ), .B2(n2360), .ZN(n4492) );
  AOI22_X1 U3539 ( .A1(n3387), .A2(\DP/RegA_out[3] ), .B1(n2409), .B2(
        DRAM_ADDR[3]), .ZN(n2598) );
  NAND2_X1 U3540 ( .A1(n2410), .A2(\DP/NPC2[3] ), .ZN(n2597) );
  OAI211_X1 U3541 ( .C1(n4492), .C2(n2413), .A(n2598), .B(n2597), .ZN(
        \DP/A[3] ) );
  INV_X1 U3542 ( .A(\DP/ALU0/S_B_MULT[3] ), .ZN(n2599) );
  NAND2_X1 U3543 ( .A1(\DP/ALU0/S_B_MULT[1] ), .A2(\DP/ALU0/S_B_MULT[2] ), 
        .ZN(n2600) );
  INV_X1 U3544 ( .A(\DP/ALU0/s_A_MULT[1] ), .ZN(n2908) );
  OAI21_X1 U3545 ( .B1(\DP/ALU0/S_B_MULT[1] ), .B2(\DP/ALU0/S_B_MULT[2] ), .A(
        n2600), .ZN(n2601) );
  INV_X1 U3546 ( .A(n2872), .ZN(n2984) );
  NOR2_X1 U3547 ( .A1(n2984), .A2(n2601), .ZN(n4496) );
  NAND2_X1 U3548 ( .A1(\DP/ALU0/S_B_MULT[3] ), .A2(n4496), .ZN(n2985) );
  INV_X1 U3549 ( .A(n2874), .ZN(n2909) );
  OAI22_X1 U3550 ( .A1(n2908), .A2(n2960), .B1(n2985), .B2(n2909), .ZN(n2602)
         );
  AOI221_X1 U3551 ( .B1(n2359), .B2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .C1(n2962), 
        .C2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .A(n2602), .ZN(n2631) );
  OAI21_X1 U3552 ( .B1(n2603), .B2(n2951), .A(n2606), .ZN(n2952) );
  AOI222_X1 U3553 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n2924), .B1(n2876), .B2(
        n2926), .C1(n2886), .C2(n2912), .ZN(n2630) );
  XNOR2_X1 U3554 ( .A(n2631), .B(n2630), .ZN(n2608) );
  AOI222_X1 U3555 ( .A1(n2926), .A2(n2874), .B1(n2924), .B2(
        \DP/ALU0/s_A_MULT[2] ), .C1(n2886), .C2(n2876), .ZN(n2607) );
  INV_X1 U3556 ( .A(n2607), .ZN(n4497) );
  NAND3_X1 U3557 ( .A1(n4496), .A2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .A3(n4497), 
        .ZN(n4495) );
  NOR2_X1 U3558 ( .A1(n2608), .A2(n4495), .ZN(n4507) );
  AOI211_X1 U3559 ( .C1(n2608), .C2(n4495), .A(n4507), .B(n4498), .ZN(n2609)
         );
  AOI21_X1 U3560 ( .B1(n3420), .B2(\DP/A[3] ), .A(n2609), .ZN(n2610) );
  INV_X1 U3561 ( .A(n2610), .ZN(\DP/ALU0/N25 ) );
  AOI22_X1 U3562 ( .A1(n2449), .A2(\DP/RegALU2_out[4] ), .B1(
        \DP/RegLMD_out[4] ), .B2(n2360), .ZN(n4506) );
  AOI22_X1 U3563 ( .A1(n2410), .A2(\DP/NPC2[4] ), .B1(n2409), .B2(DRAM_ADDR[4]), .ZN(n2612) );
  NAND2_X1 U3564 ( .A1(n2411), .A2(\DP/RegA_out[4] ), .ZN(n2611) );
  OAI211_X1 U3565 ( .C1(n4561), .C2(n2413), .A(n2612), .B(n2611), .ZN(
        \DP/A[4] ) );
  AOI22_X1 U3566 ( .A1(n200), .A2(\DP/RegALU2_out[5] ), .B1(\DP/RegLMD_out[5] ), .B2(n2360), .ZN(n4517) );
  AOI22_X1 U3567 ( .A1(n3386), .A2(\DP/NPC2[5] ), .B1(n2409), .B2(DRAM_ADDR[5]), .ZN(n2614) );
  NAND2_X1 U3568 ( .A1(n2411), .A2(\DP/RegA_out[5] ), .ZN(n2613) );
  OAI211_X1 U3569 ( .C1(n4517), .C2(n2413), .A(n2614), .B(n2613), .ZN(
        \DP/A[5] ) );
  INV_X1 U3570 ( .A(\DP/A[5] ), .ZN(n186) );
  AOI222_X1 U3571 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n2924), .B1(n2886), .B2(
        n2955), .C1(n2912), .C2(n2926), .ZN(n2627) );
  INV_X1 U3572 ( .A(\DP/ALU0/S_B_MULT[5] ), .ZN(n2650) );
  NAND2_X1 U3573 ( .A1(\DP/ALU0/S_B_MULT[3] ), .A2(\DP/ALU0/S_B_MULT[4] ), 
        .ZN(n2622) );
  OAI21_X1 U3574 ( .B1(\DP/ALU0/S_B_MULT[3] ), .B2(\DP/ALU0/S_B_MULT[4] ), .A(
        n2622), .ZN(n2616) );
  NOR2_X1 U3575 ( .A1(n2650), .A2(n2616), .ZN(n2988) );
  NAND2_X1 U3576 ( .A1(n2988), .A2(n2872), .ZN(n3076) );
  NOR2_X1 U3577 ( .A1(\DP/ALU0/S_B_MULT[5] ), .A2(n2616), .ZN(n2623) );
  OAI21_X1 U3578 ( .B1(n2963), .B2(n2623), .A(\DP/ALU0/MULT/SHIFTERi_0/N19 ), 
        .ZN(n2626) );
  INV_X1 U3579 ( .A(n2985), .ZN(n2958) );
  AOI22_X1 U3580 ( .A1(\DP/ALU0/s_A_MULT[1] ), .A2(n2962), .B1(n2958), .B2(
        n2876), .ZN(n2617) );
  OAI21_X1 U3581 ( .B1(n2951), .B2(n2960), .A(n2617), .ZN(n2618) );
  AOI21_X1 U3582 ( .B1(n2359), .B2(n2874), .A(n2618), .ZN(n2625) );
  INV_X1 U3583 ( .A(n4510), .ZN(n4508) );
  NAND2_X1 U3584 ( .A1(n4507), .A2(n4508), .ZN(n2632) );
  NAND2_X1 U3585 ( .A1(n2441), .A2(n2632), .ZN(n4512) );
  INV_X1 U3586 ( .A(\DP/ALU0/s_A_MULT[3] ), .ZN(n3002) );
  AOI22_X1 U3587 ( .A1(\DP/ALU0/s_A_MULT[2] ), .A2(n2962), .B1(n2958), .B2(
        n2912), .ZN(n2619) );
  OAI21_X1 U3588 ( .B1(n3002), .B2(n2960), .A(n2619), .ZN(n2620) );
  AOI21_X1 U3589 ( .B1(n2359), .B2(n2876), .A(n2620), .ZN(n2642) );
  INV_X1 U3590 ( .A(n55), .ZN(n3009) );
  OAI21_X1 U3591 ( .B1(n2621), .B2(n55), .A(n2637), .ZN(n3068) );
  INV_X1 U3592 ( .A(n3068), .ZN(n3006) );
  AOI222_X1 U3593 ( .A1(n3009), .A2(n2924), .B1(n2886), .B2(n3006), .C1(n2955), 
        .C2(n2926), .ZN(n2641) );
  NOR2_X1 U3594 ( .A1(\DP/ALU0/S_B_MULT[3] ), .A2(\DP/ALU0/S_B_MULT[4] ), .ZN(
        n3075) );
  NAND2_X1 U3595 ( .A1(\DP/ALU0/S_B_MULT[5] ), .A2(n3075), .ZN(n3034) );
  OAI22_X1 U3596 ( .A1(n2908), .A2(n3033), .B1(n3076), .B2(n2909), .ZN(n2624)
         );
  AOI221_X1 U3597 ( .B1(n3078), .B2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .C1(n3037), 
        .C2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .A(n2624), .ZN(n2640) );
  FA_X1 U3598 ( .A(n2627), .B(n2626), .CI(n2625), .CO(n2628), .S(n4510) );
  NOR2_X1 U3599 ( .A1(n2628), .A2(n2629), .ZN(n3435) );
  AOI21_X1 U3600 ( .B1(n2629), .B2(n2628), .A(n3435), .ZN(n3428) );
  NOR2_X1 U3601 ( .A1(n2631), .A2(n2630), .ZN(n4511) );
  INV_X1 U3602 ( .A(n4511), .ZN(n4509) );
  NOR2_X1 U3603 ( .A1(n4510), .A2(n4509), .ZN(n3427) );
  XNOR2_X1 U3604 ( .A(n3428), .B(n3427), .ZN(n3424) );
  OR2_X1 U3605 ( .A1(n4498), .A2(n2632), .ZN(n3423) );
  OAI222_X1 U3606 ( .A1(n4512), .A2(n3424), .B1(n2443), .B2(n186), .C1(n3423), 
        .C2(n3428), .ZN(\DP/ALU0/N27 ) );
  AOI22_X1 U3607 ( .A1(n200), .A2(\DP/RegALU2_out[6] ), .B1(\DP/RegLMD_out[6] ), .B2(n2360), .ZN(n4520) );
  AOI22_X1 U3608 ( .A1(n2410), .A2(\DP/NPC2[6] ), .B1(n2409), .B2(DRAM_ADDR[6]), .ZN(n2634) );
  NAND2_X1 U3609 ( .A1(n2411), .A2(\DP/RegA_out[6] ), .ZN(n2633) );
  OAI211_X1 U3610 ( .C1(n4520), .C2(n2413), .A(n2634), .B(n2633), .ZN(
        \DP/A[6] ) );
  INV_X1 U3611 ( .A(\DP/A[6] ), .ZN(n182) );
  INV_X1 U3612 ( .A(\DP/ALU0/s_A_MULT[4] ), .ZN(n3025) );
  AOI22_X1 U3613 ( .A1(n2958), .A2(n2955), .B1(n2359), .B2(n2912), .ZN(n2635)
         );
  OAI21_X1 U3614 ( .B1(n3025), .B2(n2960), .A(n2635), .ZN(n2636) );
  AOI21_X1 U3615 ( .B1(\DP/ALU0/s_A_MULT[3] ), .B2(n2962), .A(n2636), .ZN(
        n2662) );
  AOI222_X1 U3616 ( .A1(n3032), .A2(n2924), .B1(n2886), .B2(n3029), .C1(n3006), 
        .C2(n2926), .ZN(n2661) );
  AOI22_X1 U3617 ( .A1(\DP/ALU0/s_A_MULT[1] ), .A2(n3037), .B1(n2963), .B2(
        n2876), .ZN(n2638) );
  OAI21_X1 U3618 ( .B1(n2951), .B2(n3033), .A(n2638), .ZN(n2639) );
  AOI21_X1 U3619 ( .B1(n3078), .B2(n2874), .A(n2639), .ZN(n2660) );
  FA_X1 U3620 ( .A(n2642), .B(n2641), .CI(n2640), .CO(n2648), .S(n2629) );
  NAND2_X1 U3621 ( .A1(n31), .A2(n2650), .ZN(n3154) );
  OAI21_X1 U3622 ( .B1(n31), .B2(n2650), .A(n3154), .ZN(n2651) );
  NOR2_X1 U3623 ( .A1(n2984), .A2(n2651), .ZN(n2653) );
  NAND2_X1 U3624 ( .A1(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .A2(n2653), .ZN(n2647)
         );
  INV_X1 U3625 ( .A(n3430), .ZN(n3433) );
  AOI21_X1 U3626 ( .B1(n3428), .B2(n3427), .A(n3435), .ZN(n2643) );
  XOR2_X1 U3627 ( .A(n3433), .B(n2643), .Z(n2644) );
  OAI22_X1 U3628 ( .A1(n2442), .A2(n182), .B1(n2644), .B2(n4498), .ZN(
        \DP/ALU0/N28 ) );
  AOI22_X1 U3630 ( .A1(n2411), .A2(\DP/RegA_out[7] ), .B1(n2409), .B2(
        DRAM_ADDR[7]), .ZN(n2646) );
  NAND2_X1 U3631 ( .A1(n2410), .A2(\DP/NPC2[7] ), .ZN(n2645) );
  OAI211_X1 U3632 ( .C1(n3657), .C2(n2413), .A(n2646), .B(n2645), .ZN(
        \DP/A[7] ) );
  INV_X1 U3633 ( .A(\DP/A[7] ), .ZN(n178) );
  FA_X1 U3634 ( .A(n2649), .B(n2648), .CI(n2647), .CO(n2664), .S(n3430) );
  INV_X1 U3635 ( .A(n29), .ZN(n2652) );
  NOR2_X1 U3636 ( .A1(n2652), .A2(n2651), .ZN(n2693) );
  INV_X1 U3637 ( .A(n2693), .ZN(n3115) );
  NAND2_X1 U3638 ( .A1(n2653), .A2(n2652), .ZN(n3155) );
  OAI22_X1 U3639 ( .A1(n2908), .A2(n3115), .B1(n3155), .B2(n2909), .ZN(n2654)
         );
  AOI221_X1 U3640 ( .B1(n2358), .B2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .C1(n3118), 
        .C2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .A(n2654), .ZN(n2671) );
  AOI22_X1 U3641 ( .A1(n2958), .A2(n3006), .B1(n2359), .B2(n2955), .ZN(n2655)
         );
  OAI21_X1 U3642 ( .B1(n55), .B2(n2960), .A(n2655), .ZN(n2656) );
  AOI21_X1 U3643 ( .B1(\DP/ALU0/s_A_MULT[4] ), .B2(n2962), .A(n2656), .ZN(
        n2674) );
  INV_X1 U3644 ( .A(n28), .ZN(n3071) );
  OAI21_X1 U3645 ( .B1(n2657), .B2(n28), .A(n2683), .ZN(n3148) );
  INV_X1 U3646 ( .A(n3148), .ZN(n3072) );
  AOI222_X1 U3647 ( .A1(n3071), .A2(n2924), .B1(n2886), .B2(n3072), .C1(n3029), 
        .C2(n2926), .ZN(n2673) );
  AOI22_X1 U3648 ( .A1(n2963), .A2(n2912), .B1(n3078), .B2(n2876), .ZN(n2658)
         );
  OAI21_X1 U3649 ( .B1(n3002), .B2(n3033), .A(n2658), .ZN(n2659) );
  AOI21_X1 U3650 ( .B1(\DP/ALU0/s_A_MULT[2] ), .B2(n3037), .A(n2659), .ZN(
        n2672) );
  FA_X1 U3651 ( .A(n2662), .B(n2661), .CI(n2660), .CO(n2669), .S(n2649) );
  NOR2_X1 U3652 ( .A1(n2663), .A2(n2664), .ZN(n3439) );
  AOI21_X1 U3653 ( .B1(n2664), .B2(n2663), .A(n3439), .ZN(n3434) );
  NAND2_X1 U3654 ( .A1(n3435), .A2(n3433), .ZN(n2665) );
  XOR2_X1 U3655 ( .A(n3434), .B(n2665), .Z(n2666) );
  OAI22_X1 U3656 ( .A1(n2442), .A2(n178), .B1(n2666), .B2(n4498), .ZN(
        \DP/ALU0/N29 ) );
  AOI22_X1 U3657 ( .A1(n2449), .A2(\DP/RegALU2_out[8] ), .B1(
        \DP/RegLMD_out[8] ), .B2(n2448), .ZN(n4480) );
  AOI22_X1 U3658 ( .A1(n2411), .A2(\DP/RegA_out[8] ), .B1(n2409), .B2(
        DRAM_ADDR[8]), .ZN(n2668) );
  NAND2_X1 U3659 ( .A1(n2410), .A2(\DP/NPC2[8] ), .ZN(n2667) );
  OAI211_X1 U3660 ( .C1(n4548), .C2(n2413), .A(n2668), .B(n2667), .ZN(
        \DP/A[8] ) );
  INV_X1 U3661 ( .A(\DP/A[8] ), .ZN(n175) );
  FA_X1 U3662 ( .A(n2671), .B(n2670), .CI(n2669), .CO(n2689), .S(n2663) );
  FA_X1 U3663 ( .A(n2674), .B(n2673), .CI(n2672), .CO(n2708), .S(n2670) );
  AOI22_X1 U3664 ( .A1(\DP/ALU0/s_A_MULT[2] ), .A2(n2693), .B1(n2358), .B2(
        n2874), .ZN(n2676) );
  NAND2_X1 U3665 ( .A1(\DP/ALU0/s_A_MULT[1] ), .A2(n3118), .ZN(n2675) );
  OAI211_X1 U3666 ( .C1(n3155), .C2(n2952), .A(n2676), .B(n2675), .ZN(n2706)
         );
  NAND2_X1 U3667 ( .A1(n29), .A2(n54), .ZN(n3173) );
  OAI21_X1 U3668 ( .B1(n29), .B2(n54), .A(n3173), .ZN(n2690) );
  NOR2_X1 U3669 ( .A1(n2984), .A2(n2690), .ZN(n2707) );
  NAND2_X1 U3670 ( .A1(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .A2(n2707), .ZN(n2677)
         );
  XOR2_X1 U3671 ( .A(n2706), .B(n2677), .Z(n2678) );
  OR2_X1 U3672 ( .A1(n2708), .A2(n2678), .ZN(n2712) );
  NAND2_X1 U3673 ( .A1(n2708), .A2(n2678), .ZN(n2711) );
  NAND2_X1 U3674 ( .A1(n2712), .A2(n2711), .ZN(n2684) );
  AOI22_X1 U3675 ( .A1(n2958), .A2(n3029), .B1(n2359), .B2(n3006), .ZN(n2679)
         );
  OAI21_X1 U3676 ( .B1(n30), .B2(n2960), .A(n2679), .ZN(n2680) );
  AOI21_X1 U3677 ( .B1(n2962), .B2(n3009), .A(n2680), .ZN(n2700) );
  AOI22_X1 U3678 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n3037), .B1(n2963), .B2(
        n2955), .ZN(n2681) );
  OAI21_X1 U3679 ( .B1(n3025), .B2(n3033), .A(n2681), .ZN(n2682) );
  AOI21_X1 U3680 ( .B1(n3078), .B2(n2912), .A(n2682), .ZN(n2699) );
  AOI222_X1 U3681 ( .A1(n3126), .A2(n2924), .B1(n2886), .B2(n3127), .C1(n3072), 
        .C2(n2926), .ZN(n2698) );
  INV_X1 U3682 ( .A(n2709), .ZN(n2710) );
  XOR2_X1 U3683 ( .A(n2684), .B(n2710), .Z(n2688) );
  XOR2_X1 U3684 ( .A(n2689), .B(n2688), .Z(n3440) );
  XNOR2_X1 U3685 ( .A(n3440), .B(n3439), .ZN(n2685) );
  OAI22_X1 U3686 ( .A1(n4515), .A2(n175), .B1(n2685), .B2(n4498), .ZN(
        \DP/ALU0/N30 ) );
  AOI22_X1 U3687 ( .A1(n200), .A2(\DP/RegALU2_out[9] ), .B1(\DP/RegLMD_out[9] ), .B2(n2448), .ZN(n4485) );
  AOI22_X1 U3688 ( .A1(n3386), .A2(\DP/NPC2[9] ), .B1(n2409), .B2(DRAM_ADDR[9]), .ZN(n2687) );
  NAND2_X1 U3689 ( .A1(n2411), .A2(\DP/RegA_out[9] ), .ZN(n2686) );
  OAI211_X1 U3690 ( .C1(n4551), .C2(n2413), .A(n2687), .B(n2686), .ZN(
        \DP/A[9] ) );
  INV_X1 U3691 ( .A(\DP/A[9] ), .ZN(n2721) );
  NOR2_X1 U3692 ( .A1(n2689), .A2(n2688), .ZN(n3445) );
  INV_X1 U3693 ( .A(n52), .ZN(n2691) );
  NAND2_X1 U3694 ( .A1(n2707), .A2(n2691), .ZN(n3212) );
  NOR2_X1 U3695 ( .A1(n52), .A2(n3173), .ZN(n3240) );
  NAND2_X1 U3696 ( .A1(n2872), .A2(n3240), .ZN(n3214) );
  INV_X1 U3697 ( .A(n3214), .ZN(n3157) );
  NOR2_X1 U3698 ( .A1(n3157), .A2(n3177), .ZN(n2692) );
  OR2_X1 U3699 ( .A1(n2691), .A2(n2690), .ZN(n3159) );
  OAI222_X1 U3700 ( .A1(n2909), .A2(n3212), .B1(n2451), .B2(n2692), .C1(n2908), 
        .C2(n3159), .ZN(n2697) );
  INV_X1 U3701 ( .A(n3155), .ZN(n3086) );
  AOI22_X1 U3702 ( .A1(n3086), .A2(n2912), .B1(n2358), .B2(n2876), .ZN(n2695)
         );
  AOI22_X1 U3703 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n2693), .B1(
        \DP/ALU0/s_A_MULT[2] ), .B2(n3118), .ZN(n2694) );
  NAND2_X1 U3704 ( .A1(n2695), .A2(n2694), .ZN(n2696) );
  NAND2_X1 U3705 ( .A1(n2696), .A2(n2697), .ZN(n2770) );
  OAI21_X1 U3706 ( .B1(n2697), .B2(n2696), .A(n2770), .ZN(n2726) );
  FA_X1 U3707 ( .A(n2700), .B(n2699), .CI(n2698), .CO(n2725), .S(n2709) );
  AOI22_X1 U3708 ( .A1(n2958), .A2(n3072), .B1(n2359), .B2(n3029), .ZN(n2701)
         );
  OAI21_X1 U3709 ( .B1(n28), .B2(n2960), .A(n2701), .ZN(n2702) );
  AOI21_X1 U3710 ( .B1(n2962), .B2(n3032), .A(n2702), .ZN(n2740) );
  AOI22_X1 U3711 ( .A1(\DP/ALU0/s_A_MULT[4] ), .A2(n3037), .B1(n2963), .B2(
        n3006), .ZN(n2703) );
  OAI21_X1 U3712 ( .B1(n55), .B2(n3033), .A(n2703), .ZN(n2704) );
  AOI21_X1 U3713 ( .B1(n3078), .B2(n2955), .A(n2704), .ZN(n2739) );
  OAI21_X1 U3714 ( .B1(n3220), .B2(n2705), .A(n2735), .ZN(n3224) );
  INV_X1 U3715 ( .A(n3224), .ZN(n3151) );
  AOI222_X1 U3716 ( .A1(\DP/ALU0/s_A_MULT[9] ), .A2(n2924), .B1(n2886), .B2(
        n3151), .C1(n2926), .C2(n3127), .ZN(n2738) );
  NAND3_X1 U3717 ( .A1(n2707), .A2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .A3(n2706), 
        .ZN(n2714) );
  NOR3_X1 U3718 ( .A1(n2709), .A2(n2714), .A3(n2708), .ZN(n2716) );
  NAND2_X1 U3719 ( .A1(n2711), .A2(n2710), .ZN(n2713) );
  NAND3_X1 U3720 ( .A1(n2714), .A2(n2713), .A3(n2712), .ZN(n2742) );
  INV_X1 U3721 ( .A(n2742), .ZN(n2715) );
  NOR2_X1 U3722 ( .A1(n2716), .A2(n2715), .ZN(n2717) );
  NAND2_X1 U3723 ( .A1(n2718), .A2(n2717), .ZN(n2741) );
  OAI21_X1 U3724 ( .B1(n2718), .B2(n2717), .A(n2741), .ZN(n3444) );
  AOI21_X1 U3725 ( .B1(n3445), .B2(n3444), .A(n2439), .ZN(n2719) );
  OAI21_X1 U3726 ( .B1(n3445), .B2(n3444), .A(n2719), .ZN(n2720) );
  OAI21_X1 U3727 ( .B1(n2443), .B2(n2721), .A(n2720), .ZN(\DP/ALU0/N31 ) );
  AOI22_X1 U3728 ( .A1(n200), .A2(\DP/RegALU2_out[10] ), .B1(
        \DP/RegLMD_out[10] ), .B2(n2448), .ZN(n4430) );
  AOI22_X1 U3729 ( .A1(n2411), .A2(\DP/RegA_out[10] ), .B1(n2409), .B2(
        DRAM_ADDR[10]), .ZN(n2723) );
  NAND2_X1 U3730 ( .A1(n2410), .A2(\DP/NPC2[10] ), .ZN(n2722) );
  OAI211_X1 U3731 ( .C1(n4430), .C2(n2413), .A(n2723), .B(n2722), .ZN(
        \DP/A[10] ) );
  INV_X1 U3732 ( .A(\DP/A[10] ), .ZN(n2744) );
  FA_X1 U3733 ( .A(n2726), .B(n2725), .CI(n2724), .CO(n2769), .S(n2718) );
  NOR2_X1 U3734 ( .A1(n2951), .A2(n3159), .ZN(n2728) );
  OAI22_X1 U3735 ( .A1(n3212), .A2(n2952), .B1(n2909), .B2(n3214), .ZN(n2727)
         );
  AOI211_X1 U3736 ( .C1(n3177), .C2(\DP/ALU0/s_A_MULT[1] ), .A(n2728), .B(
        n2727), .ZN(n2767) );
  AOI22_X1 U3737 ( .A1(n3086), .A2(n2955), .B1(n2358), .B2(n2912), .ZN(n2729)
         );
  OAI21_X1 U3738 ( .B1(n3025), .B2(n3115), .A(n2729), .ZN(n2730) );
  AOI21_X1 U3739 ( .B1(\DP/ALU0/s_A_MULT[3] ), .B2(n3118), .A(n2730), .ZN(
        n2766) );
  NOR2_X1 U3740 ( .A1(n52), .A2(n11), .ZN(n2759) );
  AOI21_X1 U3741 ( .B1(n11), .B2(n52), .A(n2759), .ZN(n2731) );
  NAND2_X1 U3742 ( .A1(n51), .A2(n2731), .ZN(n3235) );
  INV_X1 U3743 ( .A(n3235), .ZN(n3207) );
  INV_X1 U3744 ( .A(n2731), .ZN(n2732) );
  NOR2_X1 U3745 ( .A1(n2732), .A2(n51), .ZN(n3206) );
  INV_X1 U3746 ( .A(n3206), .ZN(n3269) );
  NOR2_X1 U3747 ( .A1(n3269), .A2(n2984), .ZN(n2760) );
  OAI21_X1 U3748 ( .B1(n3207), .B2(n2760), .A(\DP/ALU0/MULT/SHIFTERi_0/N19 ), 
        .ZN(n2765) );
  AOI22_X1 U3749 ( .A1(n2958), .A2(n3127), .B1(n2359), .B2(n3072), .ZN(n2733)
         );
  OAI21_X1 U3750 ( .B1(n53), .B2(n2960), .A(n2733), .ZN(n2734) );
  AOI21_X1 U3751 ( .B1(n2962), .B2(n3071), .A(n2734), .ZN(n2754) );
  AOI222_X1 U3752 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n2924), .B1(n2886), .B2(
        n3222), .C1(n2926), .C2(n3151), .ZN(n2753) );
  AOI22_X1 U3753 ( .A1(n2963), .A2(n3029), .B1(n3078), .B2(n3006), .ZN(n2736)
         );
  OAI21_X1 U3754 ( .B1(n30), .B2(n3033), .A(n2736), .ZN(n2737) );
  AOI21_X1 U3755 ( .B1(n3037), .B2(n3009), .A(n2737), .ZN(n2752) );
  FA_X1 U3756 ( .A(n2740), .B(n2739), .CI(n2738), .CO(n2762), .S(n2724) );
  NAND2_X1 U3757 ( .A1(n2742), .A2(n2741), .ZN(n3449) );
  XNOR2_X1 U3758 ( .A(n3450), .B(n3449), .ZN(n2743) );
  OAI22_X1 U3759 ( .A1(n2442), .A2(n2744), .B1(n2743), .B2(n4498), .ZN(
        \DP/ALU0/N32 ) );
  AOI22_X1 U3760 ( .A1(n2449), .A2(\DP/RegALU2_out[11] ), .B1(
        \DP/RegLMD_out[11] ), .B2(n2448), .ZN(n4432) );
  AOI22_X1 U3761 ( .A1(n3386), .A2(\DP/NPC2[11] ), .B1(n2409), .B2(
        DRAM_ADDR[11]), .ZN(n2746) );
  NAND2_X1 U3762 ( .A1(n2411), .A2(\DP/RegA_out[11] ), .ZN(n2745) );
  OAI211_X1 U3763 ( .C1(n4565), .C2(n2413), .A(n2746), .B(n2745), .ZN(
        \DP/A[11] ) );
  INV_X1 U3764 ( .A(\DP/A[11] ), .ZN(n2772) );
  AOI22_X1 U3765 ( .A1(n2958), .A2(n3151), .B1(n2359), .B2(n3127), .ZN(n2747)
         );
  OAI21_X1 U3766 ( .B1(n3220), .B2(n2960), .A(n2747), .ZN(n2748) );
  AOI21_X1 U3767 ( .B1(n2962), .B2(n3126), .A(n2748), .ZN(n2782) );
  OAI21_X1 U3768 ( .B1(n3274), .B2(n2749), .A(n2777), .ZN(n3279) );
  INV_X1 U3769 ( .A(n3279), .ZN(n3215) );
  AOI222_X1 U3770 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n2924), .B1(n2886), .B2(
        n3215), .C1(n2926), .C2(n3222), .ZN(n2781) );
  AOI22_X1 U3771 ( .A1(n2963), .A2(n3072), .B1(n3078), .B2(n3029), .ZN(n2750)
         );
  OAI21_X1 U3772 ( .B1(n28), .B2(n3033), .A(n2750), .ZN(n2751) );
  AOI21_X1 U3773 ( .B1(n3037), .B2(n3032), .A(n2751), .ZN(n2780) );
  FA_X1 U3774 ( .A(n2754), .B(n2753), .CI(n2752), .CO(n2790), .S(n2763) );
  AOI22_X1 U3775 ( .A1(n3086), .A2(n3006), .B1(n2358), .B2(n2955), .ZN(n2755)
         );
  OAI21_X1 U3776 ( .B1(n55), .B2(n3115), .A(n2755), .ZN(n2756) );
  AOI21_X1 U3777 ( .B1(\DP/ALU0/s_A_MULT[4] ), .B2(n3118), .A(n2756), .ZN(
        n2794) );
  INV_X1 U3778 ( .A(n3212), .ZN(n3174) );
  AOI22_X1 U3779 ( .A1(n3174), .A2(n2912), .B1(n2876), .B2(n3157), .ZN(n2757)
         );
  OAI21_X1 U3780 ( .B1(n3002), .B2(n3159), .A(n2757), .ZN(n2758) );
  AOI21_X1 U3781 ( .B1(\DP/ALU0/s_A_MULT[2] ), .B2(n3177), .A(n2758), .ZN(
        n2793) );
  NAND2_X1 U3782 ( .A1(n51), .A2(n2759), .ZN(n3234) );
  INV_X1 U3783 ( .A(n3234), .ZN(n3208) );
  NAND2_X1 U3784 ( .A1(n52), .A2(n11), .ZN(n3267) );
  NOR2_X1 U3785 ( .A1(n51), .A2(n3267), .ZN(n3298) );
  OAI22_X1 U3786 ( .A1(n2908), .A2(n3235), .B1(n2909), .B2(n3236), .ZN(n2761)
         );
  AOI221_X1 U3787 ( .B1(n3208), .B2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .C1(n3270), 
        .C2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .A(n2761), .ZN(n2792) );
  FA_X1 U3788 ( .A(n2764), .B(n2763), .CI(n2762), .CO(n2799), .S(n2768) );
  FA_X1 U3789 ( .A(n2767), .B(n2766), .CI(n2765), .CO(n2798), .S(n2764) );
  FA_X1 U3790 ( .A(n2770), .B(n2769), .CI(n2768), .CO(n3454), .S(n3450) );
  XNOR2_X1 U3791 ( .A(n3455), .B(n3454), .ZN(n2771) );
  OAI22_X1 U3792 ( .A1(n2442), .A2(n2772), .B1(n2771), .B2(n4498), .ZN(
        \DP/ALU0/N33 ) );
  AOI22_X1 U3794 ( .A1(n3386), .A2(\DP/NPC2[12] ), .B1(n2409), .B2(
        \DP/RegALU1_out[12] ), .ZN(n2774) );
  NAND2_X1 U3795 ( .A1(n2411), .A2(\DP/RegA_out[12] ), .ZN(n2773) );
  INV_X1 U3797 ( .A(\DP/A[12] ), .ZN(n2802) );
  INV_X1 U3798 ( .A(\DP/ALU0/s_A_MULT[10] ), .ZN(n3246) );
  AOI22_X1 U3799 ( .A1(n2958), .A2(n3222), .B1(n2359), .B2(n3151), .ZN(n2775)
         );
  OAI21_X1 U3800 ( .B1(n3246), .B2(n2960), .A(n2775), .ZN(n2776) );
  AOI21_X1 U3801 ( .B1(\DP/ALU0/s_A_MULT[9] ), .B2(n2962), .A(n2776), .ZN(
        n2831) );
  AOI222_X1 U3802 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n2924), .B1(n2886), .B2(
        n3276), .C1(n2926), .C2(n3215), .ZN(n2830) );
  AOI22_X1 U3803 ( .A1(n3127), .A2(n2963), .B1(n3037), .B2(n3071), .ZN(n2778)
         );
  OAI21_X1 U3804 ( .B1(n53), .B2(n3033), .A(n2778), .ZN(n2779) );
  AOI21_X1 U3805 ( .B1(n3078), .B2(n3072), .A(n2779), .ZN(n2829) );
  FA_X1 U3806 ( .A(n2782), .B(n2781), .CI(n2780), .CO(n2816), .S(n2791) );
  AOI22_X1 U3807 ( .A1(n3174), .A2(n2955), .B1(n2912), .B2(n3157), .ZN(n2783)
         );
  OAI21_X1 U3808 ( .B1(n3025), .B2(n3159), .A(n2783), .ZN(n2784) );
  AOI21_X1 U3809 ( .B1(\DP/ALU0/s_A_MULT[3] ), .B2(n3177), .A(n2784), .ZN(
        n2814) );
  NOR2_X1 U3810 ( .A1(n2952), .A2(n3236), .ZN(n2786) );
  OAI22_X1 U3811 ( .A1(n2908), .A2(n3234), .B1(n2951), .B2(n3235), .ZN(n2785)
         );
  AOI211_X1 U3812 ( .C1(n3270), .C2(n2874), .A(n2786), .B(n2785), .ZN(n2813)
         );
  AOI22_X1 U3813 ( .A1(n3086), .A2(n3029), .B1(n2358), .B2(n3006), .ZN(n2787)
         );
  OAI21_X1 U3814 ( .B1(n30), .B2(n3115), .A(n2787), .ZN(n2788) );
  AOI21_X1 U3815 ( .B1(n3118), .B2(n3009), .A(n2788), .ZN(n2812) );
  FA_X1 U3816 ( .A(n2791), .B(n2790), .CI(n2789), .CO(n2806), .S(n2800) );
  NOR2_X1 U3817 ( .A1(n51), .A2(n10), .ZN(n2808) );
  AOI21_X1 U3818 ( .B1(n10), .B2(n51), .A(n2808), .ZN(n2809) );
  INV_X1 U3819 ( .A(n2809), .ZN(n2810) );
  NOR2_X1 U3820 ( .A1(n2451), .A2(n2810), .ZN(n2797) );
  FA_X1 U3821 ( .A(n2794), .B(n2793), .CI(n2792), .CO(n2795), .S(n2789) );
  INV_X1 U3822 ( .A(n2795), .ZN(n2796) );
  NAND3_X1 U3823 ( .A1(n2809), .A2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .A3(n2796), 
        .ZN(n3466) );
  OAI21_X1 U3824 ( .B1(n2797), .B2(n2796), .A(n3466), .ZN(n2805) );
  FA_X1 U3825 ( .A(n2800), .B(n2799), .CI(n2798), .CO(n3459), .S(n3455) );
  XNOR2_X1 U3826 ( .A(n3460), .B(n3459), .ZN(n2801) );
  OAI22_X1 U3827 ( .A1(n2442), .A2(n2802), .B1(n2801), .B2(n4498), .ZN(
        \DP/ALU0/N34 ) );
  AOI22_X1 U3828 ( .A1(n2449), .A2(\DP/RegALU2_out[13] ), .B1(
        \DP/RegLMD_out[13] ), .B2(n2448), .ZN(n4436) );
  AOI22_X1 U3829 ( .A1(n2411), .A2(\DP/RegA_out[13] ), .B1(n2409), .B2(
        \DP/RegALU1_out[13] ), .ZN(n2804) );
  NAND2_X1 U3830 ( .A1(n2410), .A2(\DP/NPC2[13] ), .ZN(n2803) );
  OAI211_X1 U3831 ( .C1(n4556), .C2(n2413), .A(n2804), .B(n2803), .ZN(
        \DP/A[13] ) );
  INV_X1 U3832 ( .A(\DP/A[13] ), .ZN(n2833) );
  FA_X1 U3833 ( .A(n2807), .B(n2806), .CI(n2805), .CO(n3465), .S(n3460) );
  NAND2_X1 U3834 ( .A1(n51), .A2(n10), .ZN(n3342) );
  NOR2_X1 U3835 ( .A1(n12), .A2(n3342), .ZN(n3362) );
  AND2_X1 U3836 ( .A1(n2872), .A2(n3362), .ZN(n3348) );
  NAND2_X1 U3837 ( .A1(n12), .A2(n2809), .ZN(n3307) );
  INV_X1 U3838 ( .A(n3304), .ZN(n3346) );
  OAI22_X1 U3839 ( .A1(n2908), .A2(n3307), .B1(n3346), .B2(n2909), .ZN(n2811)
         );
  AOI221_X1 U3840 ( .B1(n3348), .B2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .C1(n3310), 
        .C2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .A(n2811), .ZN(n2861) );
  FA_X1 U3841 ( .A(n2814), .B(n2813), .CI(n2812), .CO(n2860), .S(n2815) );
  XNOR2_X1 U3842 ( .A(n2861), .B(n2860), .ZN(n2864) );
  FA_X1 U3843 ( .A(n2817), .B(n2816), .CI(n2815), .CO(n2863), .S(n2807) );
  AOI22_X1 U3844 ( .A1(n3086), .A2(n3072), .B1(n2358), .B2(n3029), .ZN(n2818)
         );
  OAI21_X1 U3845 ( .B1(n28), .B2(n3115), .A(n2818), .ZN(n2819) );
  AOI21_X1 U3846 ( .B1(n3118), .B2(n3032), .A(n2819), .ZN(n2859) );
  AOI22_X1 U3847 ( .A1(n3174), .A2(n3006), .B1(n3157), .B2(n2955), .ZN(n2820)
         );
  OAI21_X1 U3848 ( .B1(n55), .B2(n3159), .A(n2820), .ZN(n2821) );
  AOI21_X1 U3849 ( .B1(\DP/ALU0/s_A_MULT[4] ), .B2(n3177), .A(n2821), .ZN(
        n2858) );
  INV_X1 U3850 ( .A(n2912), .ZN(n3003) );
  NOR2_X1 U3851 ( .A1(n3003), .A2(n3236), .ZN(n2823) );
  OAI22_X1 U3852 ( .A1(n3002), .A2(n3235), .B1(n2951), .B2(n3234), .ZN(n2822)
         );
  AOI211_X1 U3853 ( .C1(n3270), .C2(n2876), .A(n2823), .B(n2822), .ZN(n2857)
         );
  AOI22_X1 U3854 ( .A1(n2958), .A2(n3215), .B1(n2359), .B2(n3222), .ZN(n2824)
         );
  OAI21_X1 U3855 ( .B1(n3274), .B2(n2960), .A(n2824), .ZN(n2825) );
  AOI21_X1 U3856 ( .B1(\DP/ALU0/s_A_MULT[10] ), .B2(n2962), .A(n2825), .ZN(
        n2846) );
  AOI22_X1 U3857 ( .A1(n2963), .A2(n3151), .B1(n3078), .B2(n3127), .ZN(n2826)
         );
  OAI21_X1 U3858 ( .B1(n3220), .B2(n3033), .A(n2826), .ZN(n2827) );
  AOI21_X1 U3859 ( .B1(n3037), .B2(n3126), .A(n2827), .ZN(n2845) );
  OAI21_X1 U3860 ( .B1(n3350), .B2(n2828), .A(n2843), .ZN(n3349) );
  INV_X1 U3861 ( .A(n3349), .ZN(n3280) );
  AOI222_X1 U3862 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n2924), .B1(n2886), .B2(
        n3280), .C1(n2926), .C2(n3276), .ZN(n2844) );
  FA_X1 U3863 ( .A(n2831), .B(n2830), .CI(n2829), .CO(n2836), .S(n2817) );
  OAI22_X1 U3864 ( .A1(n2442), .A2(n2833), .B1(n2832), .B2(n4498), .ZN(
        \DP/ALU0/N35 ) );
  AOI22_X1 U3866 ( .A1(n3386), .A2(\DP/NPC2[14] ), .B1(n2408), .B2(
        \DP/RegALU1_out[14] ), .ZN(n2835) );
  NAND2_X1 U3867 ( .A1(n2411), .A2(\DP/RegA_out[14] ), .ZN(n2834) );
  OAI211_X1 U3868 ( .C1(n4542), .C2(n2412), .A(n2835), .B(n2834), .ZN(
        \DP/A[14] ) );
  INV_X1 U3869 ( .A(\DP/A[14] ), .ZN(n157) );
  FA_X1 U3870 ( .A(n2838), .B(n2837), .CI(n2836), .CO(n2901), .S(n2862) );
  INV_X1 U3871 ( .A(\DP/ALU0/s_A_MULT[12] ), .ZN(n3311) );
  AOI22_X1 U3872 ( .A1(n2958), .A2(n3276), .B1(n2359), .B2(n3215), .ZN(n2839)
         );
  OAI21_X1 U3873 ( .B1(n3311), .B2(n2960), .A(n2839), .ZN(n2840) );
  AOI21_X1 U3874 ( .B1(\DP/ALU0/s_A_MULT[11] ), .B2(n2962), .A(n2840), .ZN(
        n2889) );
  AOI22_X1 U3875 ( .A1(\DP/ALU0/s_A_MULT[9] ), .A2(n3037), .B1(n2963), .B2(
        n3222), .ZN(n2841) );
  OAI21_X1 U3876 ( .B1(n3246), .B2(n3033), .A(n2841), .ZN(n2842) );
  AOI21_X1 U3877 ( .B1(n3078), .B2(n3151), .A(n2842), .ZN(n2888) );
  AOI222_X1 U3878 ( .A1(n3309), .A2(n2924), .B1(n3368), .B2(n2886), .C1(n2926), 
        .C2(n3280), .ZN(n2887) );
  FA_X1 U3879 ( .A(n2846), .B(n2845), .CI(n2844), .CO(n2897), .S(n2837) );
  AOI22_X1 U3880 ( .A1(n3174), .A2(n3029), .B1(n3157), .B2(n3006), .ZN(n2847)
         );
  OAI21_X1 U3881 ( .B1(n30), .B2(n3159), .A(n2847), .ZN(n2848) );
  AOI21_X1 U3882 ( .B1(n3177), .B2(n3009), .A(n2848), .ZN(n2881) );
  INV_X1 U3883 ( .A(n2955), .ZN(n3026) );
  NOR2_X1 U3884 ( .A1(n3236), .A2(n3026), .ZN(n2850) );
  OAI22_X1 U3885 ( .A1(n3025), .A2(n3235), .B1(n3002), .B2(n3234), .ZN(n2849)
         );
  AOI211_X1 U3886 ( .C1(n3270), .C2(n2912), .A(n2850), .B(n2849), .ZN(n2880)
         );
  AOI22_X1 U3887 ( .A1(n3086), .A2(n3127), .B1(n2358), .B2(n3072), .ZN(n2851)
         );
  OAI21_X1 U3888 ( .B1(n53), .B2(n3115), .A(n2851), .ZN(n2852) );
  AOI21_X1 U3889 ( .B1(n3118), .B2(n3071), .A(n2852), .ZN(n2879) );
  AOI22_X1 U3890 ( .A1(n3304), .A2(n2876), .B1(n2874), .B2(n3348), .ZN(n2853)
         );
  OAI21_X1 U3891 ( .B1(n2951), .B2(n3307), .A(n2853), .ZN(n2854) );
  AOI21_X1 U3892 ( .B1(\DP/ALU0/s_A_MULT[1] ), .B2(n3310), .A(n2854), .ZN(
        n2870) );
  INV_X1 U3893 ( .A(n48), .ZN(n2855) );
  NAND2_X1 U3894 ( .A1(n12), .A2(n50), .ZN(n2871) );
  OAI21_X1 U3895 ( .B1(n12), .B2(n50), .A(n2871), .ZN(n2856) );
  NOR2_X1 U3896 ( .A1(n2855), .A2(n2856), .ZN(n3248) );
  NOR2_X1 U3897 ( .A1(n48), .A2(n2856), .ZN(n3376) );
  NAND2_X1 U3898 ( .A1(n3376), .A2(n2872), .ZN(n3365) );
  INV_X1 U3899 ( .A(n3365), .ZN(n3277) );
  OAI21_X1 U3900 ( .B1(n3248), .B2(n3277), .A(\DP/ALU0/MULT/SHIFTERi_0/N19 ), 
        .ZN(n2869) );
  FA_X1 U3901 ( .A(n2859), .B(n2858), .CI(n2857), .CO(n2868), .S(n2838) );
  OR2_X1 U3902 ( .A1(n2861), .A2(n2860), .ZN(n3471) );
  FA_X1 U3903 ( .A(n2864), .B(n2863), .CI(n2862), .CO(n3470), .S(n3464) );
  OAI22_X1 U3904 ( .A1(n2442), .A2(n157), .B1(n2865), .B2(n4498), .ZN(
        \DP/ALU0/N36 ) );
  AOI22_X1 U3905 ( .A1(n200), .A2(\DP/RegALU2_out[15] ), .B1(
        \DP/RegLMD_out[15] ), .B2(n2448), .ZN(n4440) );
  AOI22_X1 U3906 ( .A1(n2411), .A2(\DP/RegA_out[15] ), .B1(n2409), .B2(
        \DP/RegALU1_out[15] ), .ZN(n2867) );
  NAND2_X1 U3907 ( .A1(n2410), .A2(\DP/NPC2[15] ), .ZN(n2866) );
  OAI211_X1 U3908 ( .C1(n4440), .C2(n2412), .A(n2867), .B(n2866), .ZN(
        \DP/A[15] ) );
  INV_X1 U3909 ( .A(\DP/A[15] ), .ZN(n154) );
  FA_X1 U3910 ( .A(n2870), .B(n2869), .CI(n2868), .CO(n3478), .S(n2899) );
  NOR2_X1 U3911 ( .A1(n48), .A2(n2871), .ZN(n3393) );
  NAND2_X1 U3912 ( .A1(n3393), .A2(n2872), .ZN(n3377) );
  NOR2_X1 U3913 ( .A1(n12), .A2(n50), .ZN(n2873) );
  NAND2_X1 U3914 ( .A1(n48), .A2(n2873), .ZN(n3363) );
  NAND2_X1 U3915 ( .A1(n3377), .A2(n3363), .ZN(n2875) );
  AOI222_X1 U3916 ( .A1(n2875), .A2(\DP/ALU0/MULT/SHIFTERi_0/N19 ), .B1(n3277), 
        .B2(n2874), .C1(\DP/ALU0/s_A_MULT[1] ), .C2(n3248), .ZN(n2941) );
  AOI22_X1 U3917 ( .A1(n3304), .A2(n2912), .B1(n2876), .B2(n3348), .ZN(n2877)
         );
  OAI21_X1 U3918 ( .B1(n3002), .B2(n3307), .A(n2877), .ZN(n2878) );
  AOI21_X1 U3919 ( .B1(\DP/ALU0/s_A_MULT[2] ), .B2(n3310), .A(n2878), .ZN(
        n2940) );
  FA_X1 U3920 ( .A(n2881), .B(n2880), .CI(n2879), .CO(n2939), .S(n2896) );
  AOI22_X1 U3921 ( .A1(n2958), .A2(n3280), .B1(n2359), .B2(n3276), .ZN(n2882)
         );
  OAI21_X1 U3922 ( .B1(n3350), .B2(n2960), .A(n2882), .ZN(n2883) );
  AOI21_X1 U3923 ( .B1(\DP/ALU0/s_A_MULT[12] ), .B2(n2962), .A(n2883), .ZN(
        n2929) );
  AOI22_X1 U3924 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n3037), .B1(n2963), .B2(
        n3215), .ZN(n2884) );
  OAI21_X1 U3925 ( .B1(n3274), .B2(n3033), .A(n2884), .ZN(n2885) );
  AOI21_X1 U3926 ( .B1(n3078), .B2(n3222), .A(n2885), .ZN(n2928) );
  INV_X1 U3927 ( .A(n47), .ZN(n3343) );
  NOR2_X1 U3928 ( .A1(n2922), .A2(n47), .ZN(n3378) );
  INV_X1 U3929 ( .A(n3378), .ZN(n3347) );
  AOI222_X1 U3930 ( .A1(n3343), .A2(n2924), .B1(n2926), .B2(n3368), .C1(n3347), 
        .C2(n2886), .ZN(n2927) );
  FA_X1 U3931 ( .A(n2889), .B(n2888), .CI(n2887), .CO(n2937), .S(n2898) );
  AOI22_X1 U3932 ( .A1(n3174), .A2(n3072), .B1(n3157), .B2(n3029), .ZN(n2890)
         );
  OAI21_X1 U3933 ( .B1(n28), .B2(n3159), .A(n2890), .ZN(n2891) );
  AOI21_X1 U3934 ( .B1(n3177), .B2(n3032), .A(n2891), .ZN(n2917) );
  NOR2_X1 U3935 ( .A1(n3236), .A2(n3068), .ZN(n2893) );
  OAI22_X1 U3936 ( .A1(n55), .A2(n3235), .B1(n3025), .B2(n3234), .ZN(n2892) );
  AOI211_X1 U3937 ( .C1(n2955), .C2(n3270), .A(n2893), .B(n2892), .ZN(n2916)
         );
  AOI22_X1 U3938 ( .A1(n3086), .A2(n3151), .B1(n2358), .B2(n3127), .ZN(n2894)
         );
  OAI21_X1 U3939 ( .B1(n3220), .B2(n3115), .A(n2894), .ZN(n2895) );
  AOI21_X1 U3940 ( .B1(n3118), .B2(n3126), .A(n2895), .ZN(n2915) );
  FA_X1 U3941 ( .A(n2898), .B(n2897), .CI(n2896), .CO(n2905), .S(n2900) );
  FA_X1 U3942 ( .A(n2901), .B(n2900), .CI(n2899), .CO(n3476), .S(n3472) );
  OAI22_X1 U3943 ( .A1(n2442), .A2(n154), .B1(n2902), .B2(n2439), .ZN(
        \DP/ALU0/N37 ) );
  AOI22_X1 U3944 ( .A1(n2449), .A2(\DP/RegALU2_out[16] ), .B1(
        \DP/RegLMD_out[16] ), .B2(n2448), .ZN(n4442) );
  AOI22_X1 U3945 ( .A1(n3387), .A2(\DP/RegA_out[16] ), .B1(n2409), .B2(
        \DP/RegALU1_out[16] ), .ZN(n2903) );
  OAI21_X1 U3946 ( .B1(n4442), .B2(n2412), .A(n2903), .ZN(n2904) );
  AOI21_X1 U3947 ( .B1(n3386), .B2(\DP/NPC2[16] ), .A(n2904), .ZN(n151) );
  FA_X1 U3948 ( .A(n2907), .B(n2906), .CI(n2905), .CO(n3484), .S(n3477) );
  OAI22_X1 U3949 ( .A1(n2908), .A2(n3363), .B1(n2951), .B2(n3364), .ZN(n2911)
         );
  OAI22_X1 U3950 ( .A1(n3377), .A2(n2909), .B1(n3365), .B2(n2952), .ZN(n2910)
         );
  NOR2_X1 U3951 ( .A1(n2911), .A2(n2910), .ZN(n2980) );
  AOI22_X1 U3952 ( .A1(\DP/ALU0/s_A_MULT[3] ), .A2(n3310), .B1(n2912), .B2(
        n3348), .ZN(n2913) );
  OAI21_X1 U3953 ( .B1(n3025), .B2(n3307), .A(n2913), .ZN(n2914) );
  AOI21_X1 U3954 ( .B1(n3304), .B2(n2955), .A(n2914), .ZN(n2979) );
  FA_X1 U3955 ( .A(n2917), .B(n2916), .CI(n2915), .CO(n2978), .S(n2936) );
  AOI22_X1 U3956 ( .A1(n2958), .A2(n3368), .B1(n2359), .B2(n3280), .ZN(n2918)
         );
  OAI21_X1 U3957 ( .B1(n49), .B2(n2960), .A(n2918), .ZN(n2919) );
  AOI21_X1 U3958 ( .B1(\DP/ALU0/s_A_MULT[13] ), .B2(n2962), .A(n2919), .ZN(
        n2968) );
  AOI22_X1 U3959 ( .A1(n2963), .A2(n3276), .B1(n3078), .B2(n3215), .ZN(n2920)
         );
  OAI21_X1 U3960 ( .B1(n3311), .B2(n3033), .A(n2920), .ZN(n2921) );
  AOI21_X1 U3961 ( .B1(\DP/ALU0/s_A_MULT[11] ), .B2(n3037), .A(n2921), .ZN(
        n2967) );
  INV_X1 U3962 ( .A(n2922), .ZN(n2923) );
  NAND2_X1 U3963 ( .A1(n2923), .A2(n47), .ZN(n3345) );
  OAI22_X1 U3964 ( .A1(n3392), .A2(n2924), .B1(\DP/ALU0/S_B_MULT[1] ), .B2(
        n3343), .ZN(n3043) );
  INV_X1 U3965 ( .A(n3043), .ZN(n2925) );
  AOI21_X1 U3966 ( .B1(n2926), .B2(n3347), .A(n2925), .ZN(n2966) );
  FA_X1 U3967 ( .A(n2929), .B(n2928), .CI(n2927), .CO(n2976), .S(n2938) );
  AOI22_X1 U3968 ( .A1(n3174), .A2(n3127), .B1(n3157), .B2(n3072), .ZN(n2930)
         );
  OAI21_X1 U3969 ( .B1(n53), .B2(n3159), .A(n2930), .ZN(n2931) );
  AOI21_X1 U3970 ( .B1(n3177), .B2(n3071), .A(n2931), .ZN(n2950) );
  INV_X1 U3971 ( .A(n3029), .ZN(n3123) );
  NOR2_X1 U3972 ( .A1(n3236), .A2(n3123), .ZN(n2933) );
  OAI22_X1 U3973 ( .A1(n30), .A2(n3235), .B1(n55), .B2(n3234), .ZN(n2932) );
  AOI211_X1 U3974 ( .C1(n3006), .C2(n3270), .A(n2933), .B(n2932), .ZN(n2949)
         );
  AOI22_X1 U3975 ( .A1(n3086), .A2(n3222), .B1(n2358), .B2(n3151), .ZN(n2934)
         );
  OAI21_X1 U3976 ( .B1(n3246), .B2(n3115), .A(n2934), .ZN(n2935) );
  AOI21_X1 U3977 ( .B1(\DP/ALU0/s_A_MULT[9] ), .B2(n3118), .A(n2935), .ZN(
        n2948) );
  FA_X1 U3978 ( .A(n2938), .B(n2937), .CI(n2936), .CO(n2945), .S(n2906) );
  FA_X1 U3979 ( .A(n2941), .B(n2940), .CI(n2939), .CO(n3482), .S(n2907) );
  OAI22_X1 U3980 ( .A1(n2443), .A2(n151), .B1(n2942), .B2(n4498), .ZN(
        \DP/ALU0/N38 ) );
  AOI22_X1 U3981 ( .A1(n2449), .A2(\DP/RegALU2_out[17] ), .B1(
        \DP/RegLMD_out[17] ), .B2(n2448), .ZN(n4444) );
  AOI22_X1 U3982 ( .A1(n3387), .A2(\DP/RegA_out[17] ), .B1(n2408), .B2(
        \DP/RegALU1_out[17] ), .ZN(n2943) );
  OAI21_X1 U3983 ( .B1(n4444), .B2(n2412), .A(n2943), .ZN(n2944) );
  AOI21_X1 U3984 ( .B1(n2410), .B2(\DP/NPC2[17] ), .A(n2944), .ZN(n148) );
  FA_X1 U3985 ( .A(n2947), .B(n2946), .CI(n2945), .CO(n3490), .S(n3483) );
  FA_X1 U3986 ( .A(n2950), .B(n2949), .CI(n2948), .CO(n3018), .S(n2975) );
  OAI22_X1 U3987 ( .A1(n3002), .A2(n3364), .B1(n2951), .B2(n3363), .ZN(n2954)
         );
  OAI22_X1 U3988 ( .A1(n3377), .A2(n2952), .B1(n3365), .B2(n3003), .ZN(n2953)
         );
  NOR2_X1 U3989 ( .A1(n2954), .A2(n2953), .ZN(n3017) );
  AOI22_X1 U3990 ( .A1(n3304), .A2(n3006), .B1(n3348), .B2(n2955), .ZN(n2956)
         );
  OAI21_X1 U3991 ( .B1(n55), .B2(n3307), .A(n2956), .ZN(n2957) );
  AOI21_X1 U3992 ( .B1(\DP/ALU0/s_A_MULT[4] ), .B2(n3310), .A(n2957), .ZN(
        n3016) );
  AOI22_X1 U3993 ( .A1(n3368), .A2(n2359), .B1(n2958), .B2(n3347), .ZN(n2959)
         );
  OAI21_X1 U3994 ( .B1(n47), .B2(n2960), .A(n2959), .ZN(n2961) );
  AOI21_X1 U3995 ( .B1(n2962), .B2(n3309), .A(n2961), .ZN(n2992) );
  AOI22_X1 U3996 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n3037), .B1(n2963), .B2(
        n3280), .ZN(n2964) );
  OAI21_X1 U3997 ( .B1(n3350), .B2(n3033), .A(n2964), .ZN(n2965) );
  AOI21_X1 U3998 ( .B1(n3078), .B2(n3276), .A(n2965), .ZN(n2991) );
  FA_X1 U3999 ( .A(n2968), .B(n2967), .CI(n2966), .CO(n3011), .S(n2977) );
  AOI22_X1 U4000 ( .A1(n3174), .A2(n3151), .B1(n3157), .B2(n3127), .ZN(n2969)
         );
  OAI21_X1 U4001 ( .B1(n3220), .B2(n3159), .A(n2969), .ZN(n2970) );
  AOI21_X1 U4002 ( .B1(n3177), .B2(n3126), .A(n2970), .ZN(n3001) );
  NOR2_X1 U4003 ( .A1(n3236), .A2(n3148), .ZN(n2972) );
  OAI22_X1 U4004 ( .A1(n28), .A2(n3235), .B1(n30), .B2(n3234), .ZN(n2971) );
  AOI211_X1 U4005 ( .C1(n3029), .C2(n3270), .A(n2972), .B(n2971), .ZN(n3000)
         );
  AOI22_X1 U4006 ( .A1(n3086), .A2(n3215), .B1(n2358), .B2(n3222), .ZN(n2973)
         );
  OAI21_X1 U4007 ( .B1(n3274), .B2(n3115), .A(n2973), .ZN(n2974) );
  AOI21_X1 U4008 ( .B1(\DP/ALU0/s_A_MULT[10] ), .B2(n3118), .A(n2974), .ZN(
        n2999) );
  FA_X1 U4009 ( .A(n2977), .B(n2976), .CI(n2975), .CO(n3013), .S(n2946) );
  FA_X1 U4010 ( .A(n2980), .B(n2979), .CI(n2978), .CO(n3488), .S(n2947) );
  OAI22_X1 U4011 ( .A1(n4515), .A2(n148), .B1(n2981), .B2(n2439), .ZN(
        \DP/ALU0/N39 ) );
  AOI22_X1 U4013 ( .A1(n3386), .A2(\DP/NPC2[18] ), .B1(n2409), .B2(
        \DP/RegALU1_out[18] ), .ZN(n2982) );
  OAI21_X1 U4014 ( .B1(n4756), .B2(n2412), .A(n2982), .ZN(n2983) );
  AOI21_X1 U4015 ( .B1(n2411), .B2(\DP/RegA_out[18] ), .A(n2983), .ZN(n145) );
  NOR2_X1 U4016 ( .A1(n2984), .A2(n3378), .ZN(n3305) );
  NAND2_X1 U4017 ( .A1(\DP/ALU0/S_B_MULT[3] ), .A2(n3343), .ZN(n3039) );
  NOR2_X1 U4018 ( .A1(\DP/ALU0/S_B_MULT[1] ), .A2(\DP/ALU0/S_B_MULT[2] ), .ZN(
        n2986) );
  OAI21_X1 U4019 ( .B1(n47), .B2(n2986), .A(n2985), .ZN(n2987) );
  AOI22_X1 U4020 ( .A1(n3305), .A2(n2359), .B1(n3039), .B2(n2987), .ZN(n3042)
         );
  AOI22_X1 U4021 ( .A1(n2988), .A2(n3368), .B1(n3078), .B2(n3280), .ZN(n2989)
         );
  OAI21_X1 U4022 ( .B1(n49), .B2(n3033), .A(n2989), .ZN(n2990) );
  AOI21_X1 U4023 ( .B1(\DP/ALU0/s_A_MULT[13] ), .B2(n3037), .A(n2990), .ZN(
        n3041) );
  FA_X1 U4024 ( .A(n3043), .B(n2992), .CI(n2991), .CO(n3051), .S(n3012) );
  AOI22_X1 U4025 ( .A1(n3174), .A2(n3222), .B1(n3157), .B2(n3151), .ZN(n2993)
         );
  OAI21_X1 U4026 ( .B1(n3246), .B2(n3159), .A(n2993), .ZN(n2994) );
  AOI21_X1 U4027 ( .B1(\DP/ALU0/s_A_MULT[9] ), .B2(n3177), .A(n2994), .ZN(
        n3024) );
  INV_X1 U4028 ( .A(n3127), .ZN(n3185) );
  NOR2_X1 U4029 ( .A1(n3236), .A2(n3185), .ZN(n2996) );
  OAI22_X1 U4030 ( .A1(n53), .A2(n3235), .B1(n28), .B2(n3234), .ZN(n2995) );
  AOI211_X1 U4031 ( .C1(n3072), .C2(n3270), .A(n2996), .B(n2995), .ZN(n3023)
         );
  AOI22_X1 U4032 ( .A1(n3086), .A2(n3276), .B1(n2358), .B2(n3215), .ZN(n2997)
         );
  OAI21_X1 U4033 ( .B1(n3311), .B2(n3115), .A(n2997), .ZN(n2998) );
  AOI21_X1 U4034 ( .B1(\DP/ALU0/s_A_MULT[11] ), .B2(n3118), .A(n2998), .ZN(
        n3022) );
  FA_X1 U4035 ( .A(n3001), .B(n3000), .CI(n2999), .CO(n3058), .S(n3010) );
  OAI22_X1 U4036 ( .A1(n3025), .A2(n3364), .B1(n3002), .B2(n3363), .ZN(n3005)
         );
  OAI22_X1 U4037 ( .A1(n3377), .A2(n3003), .B1(n3365), .B2(n3026), .ZN(n3004)
         );
  NOR2_X1 U4038 ( .A1(n3005), .A2(n3004), .ZN(n3057) );
  AOI22_X1 U4039 ( .A1(n3304), .A2(n3029), .B1(n3348), .B2(n3006), .ZN(n3007)
         );
  OAI21_X1 U4040 ( .B1(n30), .B2(n3307), .A(n3007), .ZN(n3008) );
  AOI21_X1 U4041 ( .B1(n3310), .B2(n3009), .A(n3008), .ZN(n3056) );
  FA_X1 U4042 ( .A(n3012), .B(n3011), .CI(n3010), .CO(n3053), .S(n3014) );
  FA_X1 U4043 ( .A(n3015), .B(n3014), .CI(n3013), .CO(n3495), .S(n3489) );
  FA_X1 U4044 ( .A(n3018), .B(n3017), .CI(n3016), .CO(n3494), .S(n3015) );
  OAI22_X1 U4045 ( .A1(n2442), .A2(n145), .B1(n3019), .B2(n4498), .ZN(
        \DP/ALU0/N40 ) );
  AOI22_X1 U4046 ( .A1(n2449), .A2(\DP/RegALU2_out[19] ), .B1(
        \DP/RegLMD_out[19] ), .B2(n2360), .ZN(n4448) );
  AOI22_X1 U4047 ( .A1(n3387), .A2(\DP/RegA_out[19] ), .B1(n2408), .B2(
        \DP/RegALU1_out[19] ), .ZN(n3020) );
  OAI21_X1 U4048 ( .B1(n4448), .B2(n2412), .A(n3020), .ZN(n3021) );
  AOI21_X1 U4049 ( .B1(n3386), .B2(\DP/NPC2[19] ), .A(n3021), .ZN(n142) );
  FA_X1 U4050 ( .A(n3024), .B(n3023), .CI(n3022), .CO(n3096), .S(n3050) );
  OAI22_X1 U4051 ( .A1(n55), .A2(n3364), .B1(n3025), .B2(n3363), .ZN(n3028) );
  OAI22_X1 U4052 ( .A1(n3377), .A2(n3026), .B1(n3365), .B2(n3068), .ZN(n3027)
         );
  NOR2_X1 U4053 ( .A1(n3028), .A2(n3027), .ZN(n3095) );
  AOI22_X1 U4054 ( .A1(n3304), .A2(n3072), .B1(n3348), .B2(n3029), .ZN(n3030)
         );
  OAI21_X1 U4055 ( .B1(n28), .B2(n3307), .A(n3030), .ZN(n3031) );
  AOI21_X1 U4056 ( .B1(n3310), .B2(n3032), .A(n3031), .ZN(n3094) );
  NOR2_X1 U4057 ( .A1(n47), .A2(n3033), .ZN(n3036) );
  INV_X1 U4058 ( .A(n3368), .ZN(n3114) );
  OAI22_X1 U4059 ( .A1(n3378), .A2(n3076), .B1(n3114), .B2(n3034), .ZN(n3035)
         );
  AOI211_X1 U4060 ( .C1(n3037), .C2(n3309), .A(n3036), .B(n3035), .ZN(n3081)
         );
  INV_X1 U4061 ( .A(n3042), .ZN(n3038) );
  NAND2_X1 U4062 ( .A1(n3039), .A2(n3038), .ZN(n3040) );
  NAND2_X1 U4063 ( .A1(n3043), .A2(n3040), .ZN(n3104) );
  NOR2_X1 U4064 ( .A1(n3043), .A2(n3040), .ZN(n3105) );
  INV_X1 U4065 ( .A(n3105), .ZN(n3080) );
  NAND2_X1 U4066 ( .A1(n3104), .A2(n3080), .ZN(n3107) );
  XNOR2_X1 U4067 ( .A(n3081), .B(n3107), .ZN(n3093) );
  FA_X1 U4068 ( .A(n3043), .B(n3042), .CI(n3041), .CO(n3092), .S(n3052) );
  AOI22_X1 U4069 ( .A1(n3174), .A2(n3215), .B1(n3157), .B2(n3222), .ZN(n3044)
         );
  OAI21_X1 U4070 ( .B1(n3274), .B2(n3159), .A(n3044), .ZN(n3045) );
  AOI21_X1 U4071 ( .B1(\DP/ALU0/s_A_MULT[10] ), .B2(n3177), .A(n3045), .ZN(
        n3067) );
  NOR2_X1 U4072 ( .A1(n3236), .A2(n3224), .ZN(n3047) );
  OAI22_X1 U4073 ( .A1(n53), .A2(n3234), .B1(n3220), .B2(n3235), .ZN(n3046) );
  AOI211_X1 U4074 ( .C1(n3127), .C2(n3270), .A(n3047), .B(n3046), .ZN(n3066)
         );
  AOI22_X1 U4075 ( .A1(n3086), .A2(n3280), .B1(n2358), .B2(n3276), .ZN(n3048)
         );
  OAI21_X1 U4076 ( .B1(n3350), .B2(n3115), .A(n3048), .ZN(n3049) );
  AOI21_X1 U4077 ( .B1(\DP/ALU0/s_A_MULT[12] ), .B2(n3118), .A(n3049), .ZN(
        n3065) );
  FA_X1 U4078 ( .A(n3052), .B(n3051), .CI(n3050), .CO(n3062), .S(n3055) );
  FA_X1 U4079 ( .A(n3055), .B(n3054), .CI(n3053), .CO(n3501), .S(n3496) );
  FA_X1 U4080 ( .A(n3058), .B(n3057), .CI(n3056), .CO(n3500), .S(n3054) );
  OAI22_X1 U4081 ( .A1(n2442), .A2(n142), .B1(n3059), .B2(n2439), .ZN(
        \DP/ALU0/N41 ) );
  AOI22_X1 U4082 ( .A1(n200), .A2(\DP/RegALU2_out[20] ), .B1(
        \DP/RegLMD_out[20] ), .B2(n2360), .ZN(n4450) );
  AOI22_X1 U4083 ( .A1(n3387), .A2(\DP/RegA_out[20] ), .B1(n2408), .B2(
        \DP/RegALU1_out[20] ), .ZN(n3060) );
  OAI21_X1 U4084 ( .B1(n4450), .B2(n2412), .A(n3060), .ZN(n3061) );
  AOI21_X1 U4085 ( .B1(n2410), .B2(\DP/NPC2[20] ), .A(n3061), .ZN(n139) );
  FA_X1 U4086 ( .A(n3064), .B(n3063), .CI(n3062), .CO(n3508), .S(n3502) );
  FA_X1 U4087 ( .A(n3067), .B(n3066), .CI(n3065), .CO(n3137), .S(n3091) );
  OAI22_X1 U4088 ( .A1(n30), .A2(n3364), .B1(n55), .B2(n3363), .ZN(n3070) );
  OAI22_X1 U4089 ( .A1(n3377), .A2(n3068), .B1(n3365), .B2(n3123), .ZN(n3069)
         );
  NOR2_X1 U4090 ( .A1(n3070), .A2(n3069), .ZN(n3136) );
  AOI22_X1 U4091 ( .A1(n3072), .A2(n3348), .B1(n3310), .B2(n3071), .ZN(n3073)
         );
  OAI21_X1 U4092 ( .B1(n53), .B2(n3307), .A(n3073), .ZN(n3074) );
  AOI21_X1 U4093 ( .B1(n3304), .B2(n3127), .A(n3074), .ZN(n3135) );
  OAI21_X1 U4094 ( .B1(\DP/ALU0/S_B_MULT[5] ), .B2(n3075), .A(n3343), .ZN(
        n3108) );
  NAND2_X1 U4095 ( .A1(n47), .A2(n3076), .ZN(n3077) );
  AOI22_X1 U4096 ( .A1(n3078), .A2(n3347), .B1(n3108), .B2(n3077), .ZN(n3109)
         );
  XOR2_X1 U4097 ( .A(n3109), .B(n3107), .Z(n3133) );
  INV_X1 U4098 ( .A(n3104), .ZN(n3079) );
  AOI21_X1 U4099 ( .B1(n3081), .B2(n3080), .A(n3079), .ZN(n3132) );
  AOI22_X1 U4100 ( .A1(n3174), .A2(n3276), .B1(n3157), .B2(n3215), .ZN(n3082)
         );
  OAI21_X1 U4101 ( .B1(n3311), .B2(n3159), .A(n3082), .ZN(n3083) );
  AOI21_X1 U4102 ( .B1(\DP/ALU0/s_A_MULT[11] ), .B2(n3177), .A(n3083), .ZN(
        n3122) );
  INV_X1 U4103 ( .A(n3222), .ZN(n3245) );
  NOR2_X1 U4104 ( .A1(n3236), .A2(n3245), .ZN(n3085) );
  OAI22_X1 U4105 ( .A1(n3246), .A2(n3235), .B1(n3220), .B2(n3234), .ZN(n3084)
         );
  AOI211_X1 U4106 ( .C1(n3151), .C2(n3270), .A(n3085), .B(n3084), .ZN(n3121)
         );
  AOI22_X1 U4107 ( .A1(n3086), .A2(n3368), .B1(n2358), .B2(n3280), .ZN(n3087)
         );
  OAI21_X1 U4108 ( .B1(n49), .B2(n3115), .A(n3087), .ZN(n3088) );
  AOI21_X1 U4109 ( .B1(\DP/ALU0/s_A_MULT[13] ), .B2(n3118), .A(n3088), .ZN(
        n3120) );
  INV_X1 U4110 ( .A(n3089), .ZN(n3131) );
  INV_X1 U4111 ( .A(n3090), .ZN(n3101) );
  FA_X1 U4112 ( .A(n3093), .B(n3092), .CI(n3091), .CO(n3100), .S(n3063) );
  FA_X1 U4113 ( .A(n3096), .B(n3095), .CI(n3094), .CO(n3506), .S(n3064) );
  OAI22_X1 U4114 ( .A1(n2442), .A2(n139), .B1(n3097), .B2(n4498), .ZN(
        \DP/ALU0/N42 ) );
  AOI22_X1 U4115 ( .A1(n2449), .A2(\DP/RegALU2_out[21] ), .B1(
        \DP/RegLMD_out[21] ), .B2(n2360), .ZN(n4452) );
  AOI22_X1 U4116 ( .A1(n3387), .A2(\DP/RegA_out[21] ), .B1(n2408), .B2(
        \DP/RegALU1_out[21] ), .ZN(n3098) );
  OAI21_X1 U4117 ( .B1(n4554), .B2(n2412), .A(n3098), .ZN(n3099) );
  AOI21_X1 U4118 ( .B1(n2410), .B2(\DP/NPC2[21] ), .A(n3099), .ZN(n136) );
  FA_X1 U4119 ( .A(n3102), .B(n3101), .CI(n3100), .CO(n3514), .S(n3507) );
  INV_X1 U4120 ( .A(n3108), .ZN(n3103) );
  NOR2_X1 U4121 ( .A1(n3103), .A2(n3109), .ZN(n3106) );
  NOR2_X1 U4122 ( .A1(n3106), .A2(n3104), .ZN(n3302) );
  NAND2_X1 U4123 ( .A1(n3106), .A2(n3105), .ZN(n3337) );
  INV_X1 U4124 ( .A(n3337), .ZN(n3243) );
  NOR2_X1 U4125 ( .A1(n3302), .A2(n3243), .ZN(n3301) );
  INV_X1 U4126 ( .A(n3301), .ZN(n3300) );
  NOR3_X1 U4127 ( .A1(n3109), .A2(n3108), .A3(n3107), .ZN(n3165) );
  NOR2_X1 U4128 ( .A1(n3300), .A2(n3165), .ZN(n3119) );
  AOI22_X1 U4129 ( .A1(n3174), .A2(n3280), .B1(n3157), .B2(n3276), .ZN(n3110)
         );
  OAI21_X1 U4130 ( .B1(n3350), .B2(n3159), .A(n3110), .ZN(n3111) );
  AOI21_X1 U4131 ( .B1(\DP/ALU0/s_A_MULT[12] ), .B2(n3177), .A(n3111), .ZN(
        n3147) );
  NOR2_X1 U4132 ( .A1(n3236), .A2(n3279), .ZN(n3113) );
  OAI22_X1 U4133 ( .A1(n3274), .A2(n3235), .B1(n3246), .B2(n3234), .ZN(n3112)
         );
  AOI211_X1 U4134 ( .C1(n3222), .C2(n3270), .A(n3113), .B(n3112), .ZN(n3146)
         );
  NOR3_X1 U4135 ( .A1(n29), .A2(n3154), .A3(n3114), .ZN(n3117) );
  OAI22_X1 U4136 ( .A1(n47), .A2(n3115), .B1(n3378), .B2(n3155), .ZN(n3116) );
  AOI211_X1 U4137 ( .C1(n3118), .C2(n3309), .A(n3117), .B(n3116), .ZN(n3145)
         );
  XNOR2_X1 U4138 ( .A(n3119), .B(n3163), .ZN(n3143) );
  FA_X1 U4139 ( .A(n3122), .B(n3121), .CI(n3120), .CO(n3168), .S(n3089) );
  OAI22_X1 U4140 ( .A1(n28), .A2(n3364), .B1(n30), .B2(n3363), .ZN(n3125) );
  OAI22_X1 U4141 ( .A1(n3377), .A2(n3123), .B1(n3365), .B2(n3148), .ZN(n3124)
         );
  NOR2_X1 U4142 ( .A1(n3125), .A2(n3124), .ZN(n3167) );
  AOI22_X1 U4143 ( .A1(n3127), .A2(n3348), .B1(n3310), .B2(n3126), .ZN(n3128)
         );
  OAI21_X1 U4144 ( .B1(n3220), .B2(n3307), .A(n3128), .ZN(n3129) );
  AOI21_X1 U4145 ( .B1(n3304), .B2(n3151), .A(n3129), .ZN(n3166) );
  INV_X1 U4146 ( .A(n3130), .ZN(n3142) );
  FA_X1 U4147 ( .A(n3133), .B(n3132), .CI(n3131), .CO(n3141), .S(n3090) );
  INV_X1 U4148 ( .A(n3134), .ZN(n3513) );
  FA_X1 U4149 ( .A(n3137), .B(n3136), .CI(n3135), .CO(n3512), .S(n3102) );
  OAI22_X1 U4150 ( .A1(n2443), .A2(n136), .B1(n3138), .B2(n2439), .ZN(
        \DP/ALU0/N43 ) );
  AOI22_X1 U4151 ( .A1(n200), .A2(\DP/RegALU2_out[22] ), .B1(
        \DP/RegLMD_out[22] ), .B2(n2360), .ZN(n4454) );
  AOI22_X1 U4152 ( .A1(n3387), .A2(\DP/RegA_out[22] ), .B1(n2408), .B2(
        \DP/RegALU1_out[22] ), .ZN(n3139) );
  OAI21_X1 U4153 ( .B1(n4454), .B2(n2412), .A(n3139), .ZN(n3140) );
  AOI21_X1 U4154 ( .B1(n2410), .B2(\DP/NPC2[22] ), .A(n3140), .ZN(n133) );
  FA_X1 U4155 ( .A(n3143), .B(n3142), .CI(n3141), .CO(n3144), .S(n3134) );
  INV_X1 U4156 ( .A(n3144), .ZN(n3520) );
  FA_X1 U4157 ( .A(n3147), .B(n3146), .CI(n3145), .CO(n3198), .S(n3163) );
  OAI22_X1 U4158 ( .A1(n53), .A2(n3364), .B1(n28), .B2(n3363), .ZN(n3150) );
  OAI22_X1 U4159 ( .A1(n3377), .A2(n3148), .B1(n3365), .B2(n3185), .ZN(n3149)
         );
  NOR2_X1 U4160 ( .A1(n3150), .A2(n3149), .ZN(n3197) );
  AOI22_X1 U4161 ( .A1(n3304), .A2(n3222), .B1(n3348), .B2(n3151), .ZN(n3152)
         );
  OAI21_X1 U4162 ( .B1(n3246), .B2(n3307), .A(n3152), .ZN(n3153) );
  AOI21_X1 U4163 ( .B1(\DP/ALU0/s_A_MULT[9] ), .B2(n3310), .A(n3153), .ZN(
        n3196) );
  AOI21_X1 U4164 ( .B1(n29), .B2(n3154), .A(n47), .ZN(n3172) );
  AOI21_X1 U4165 ( .B1(n47), .B2(n3155), .A(n3172), .ZN(n3156) );
  AOI21_X1 U4166 ( .B1(n2358), .B2(n3347), .A(n3156), .ZN(n3190) );
  AOI22_X1 U4167 ( .A1(n3174), .A2(n3368), .B1(n3157), .B2(n3280), .ZN(n3158)
         );
  OAI21_X1 U4168 ( .B1(n49), .B2(n3159), .A(n3158), .ZN(n3160) );
  AOI21_X1 U4169 ( .B1(\DP/ALU0/s_A_MULT[13] ), .B2(n3177), .A(n3160), .ZN(
        n3189) );
  INV_X1 U4170 ( .A(n3276), .ZN(n3312) );
  NOR2_X1 U4171 ( .A1(n3236), .A2(n3312), .ZN(n3162) );
  OAI22_X1 U4172 ( .A1(n3311), .A2(n3235), .B1(n3274), .B2(n3234), .ZN(n3161)
         );
  AOI211_X1 U4173 ( .C1(n3215), .C2(n3270), .A(n3162), .B(n3161), .ZN(n3188)
         );
  XOR2_X1 U4174 ( .A(n3182), .B(n3301), .Z(n3194) );
  NAND2_X1 U4175 ( .A1(n3337), .A2(n3163), .ZN(n3164) );
  INV_X1 U4176 ( .A(n3302), .ZN(n3336) );
  OAI21_X1 U4177 ( .B1(n3165), .B2(n3164), .A(n3336), .ZN(n3193) );
  FA_X1 U4178 ( .A(n3168), .B(n3167), .CI(n3166), .CO(n3518), .S(n3130) );
  OAI22_X1 U4179 ( .A1(n2443), .A2(n133), .B1(n3169), .B2(n4498), .ZN(
        \DP/ALU0/N44 ) );
  MUX2_X1 U4180 ( .A(\DP/RegALU2_out[23] ), .B(\DP/RegLMD_out[23] ), .S(n2360), 
        .Z(n4455) );
  AOI22_X1 U4181 ( .A1(n2411), .A2(\DP/RegA_out[23] ), .B1(n2383), .B2(n4455), 
        .ZN(n3170) );
  OAI21_X1 U4182 ( .B1(n2386), .B2(n2366), .A(n3170), .ZN(n3171) );
  AOI21_X1 U4183 ( .B1(n2410), .B2(\DP/NPC2[23] ), .A(n3171), .ZN(n130) );
  NOR2_X1 U4184 ( .A1(n3172), .A2(n3190), .ZN(n3254) );
  NOR2_X1 U4185 ( .A1(n29), .A2(n54), .ZN(n3179) );
  NAND3_X1 U4186 ( .A1(n52), .A2(n3343), .A3(n3173), .ZN(n3211) );
  AOI22_X1 U4187 ( .A1(n3347), .A2(n3174), .B1(n3240), .B2(n3368), .ZN(n3175)
         );
  INV_X1 U4188 ( .A(n3175), .ZN(n3176) );
  AOI21_X1 U4189 ( .B1(n3177), .B2(n3309), .A(n3176), .ZN(n3178) );
  OAI21_X1 U4190 ( .B1(n3179), .B2(n3211), .A(n3178), .ZN(n3219) );
  OAI22_X1 U4191 ( .A1(n3350), .A2(n3235), .B1(n3311), .B2(n3234), .ZN(n3180)
         );
  AOI21_X1 U4192 ( .B1(n3270), .B2(n3276), .A(n3180), .ZN(n3181) );
  OAI21_X1 U4193 ( .B1(n3236), .B2(n3349), .A(n3181), .ZN(n3218) );
  XOR2_X1 U4194 ( .A(n3225), .B(n3301), .Z(n3204) );
  AOI21_X1 U4195 ( .B1(n3182), .B2(n3337), .A(n3302), .ZN(n3203) );
  AOI22_X1 U4196 ( .A1(\DP/ALU0/s_A_MULT[10] ), .A2(n3310), .B1(n3348), .B2(
        n3222), .ZN(n3183) );
  OAI21_X1 U4197 ( .B1(n3274), .B2(n3307), .A(n3183), .ZN(n3184) );
  AOI21_X1 U4198 ( .B1(n3304), .B2(n3215), .A(n3184), .ZN(n3230) );
  OAI22_X1 U4199 ( .A1(n53), .A2(n3363), .B1(n3220), .B2(n3364), .ZN(n3187) );
  OAI22_X1 U4200 ( .A1(n3377), .A2(n3185), .B1(n3365), .B2(n3224), .ZN(n3186)
         );
  NOR2_X1 U4201 ( .A1(n3187), .A2(n3186), .ZN(n3229) );
  FA_X1 U4202 ( .A(n3190), .B(n3189), .CI(n3188), .CO(n3228), .S(n3182) );
  INV_X1 U4203 ( .A(n3191), .ZN(n3202) );
  INV_X1 U4204 ( .A(n3192), .ZN(n3526) );
  FA_X1 U4205 ( .A(n3195), .B(n3194), .CI(n3193), .CO(n3525), .S(n3519) );
  FA_X1 U4206 ( .A(n3198), .B(n3197), .CI(n3196), .CO(n3524), .S(n3195) );
  OAI22_X1 U4207 ( .A1(n2443), .A2(n130), .B1(n3199), .B2(n2439), .ZN(
        \DP/ALU0/N45 ) );
  MUX2_X1 U4208 ( .A(\DP/RegALU2_out[24] ), .B(\DP/RegLMD_out[24] ), .S(n2360), 
        .Z(n4457) );
  AOI22_X1 U4209 ( .A1(n2408), .A2(\DP/RegALU1_out[24] ), .B1(n2383), .B2(
        n4457), .ZN(n3201) );
  AOI22_X1 U4210 ( .A1(n2411), .A2(\DP/RegA_out[24] ), .B1(n2410), .B2(
        \DP/NPC2[24] ), .ZN(n3200) );
  NAND2_X1 U4211 ( .A1(n3201), .A2(n3200), .ZN(\DP/A[24] ) );
  INV_X1 U4212 ( .A(\DP/A[24] ), .ZN(n127) );
  FA_X1 U4213 ( .A(n3204), .B(n3203), .CI(n3202), .CO(n3205), .S(n3192) );
  INV_X1 U4214 ( .A(n3205), .ZN(n3532) );
  AOI22_X1 U4215 ( .A1(n3206), .A2(n3368), .B1(n3270), .B2(n3280), .ZN(n3210)
         );
  AOI22_X1 U4216 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n3208), .B1(n3207), .B2(
        n3309), .ZN(n3209) );
  NAND2_X1 U4217 ( .A1(n3210), .A2(n3209), .ZN(n3253) );
  OAI21_X1 U4218 ( .B1(n3212), .B2(n3343), .A(n3211), .ZN(n3239) );
  INV_X1 U4219 ( .A(n3239), .ZN(n3213) );
  OAI21_X1 U4220 ( .B1(n3378), .B2(n3214), .A(n3213), .ZN(n3252) );
  XOR2_X1 U4221 ( .A(n3244), .B(n3301), .Z(n3259) );
  AOI22_X1 U4222 ( .A1(n3304), .A2(n3276), .B1(n3348), .B2(n3215), .ZN(n3217)
         );
  NAND2_X1 U4223 ( .A1(\DP/ALU0/s_A_MULT[11] ), .A2(n3310), .ZN(n3216) );
  OAI211_X1 U4224 ( .C1(n3307), .C2(n3311), .A(n3217), .B(n3216), .ZN(n3262)
         );
  FA_X1 U4225 ( .A(n3254), .B(n3219), .CI(n3218), .CO(n3261), .S(n3225) );
  OAI22_X1 U4226 ( .A1(n3246), .A2(n3364), .B1(n3220), .B2(n3363), .ZN(n3221)
         );
  AOI21_X1 U4227 ( .B1(n3277), .B2(n3222), .A(n3221), .ZN(n3223) );
  OAI21_X1 U4228 ( .B1(n3377), .B2(n3224), .A(n3223), .ZN(n3260) );
  NOR2_X1 U4229 ( .A1(n3225), .A2(n3300), .ZN(n3226) );
  NOR2_X1 U4230 ( .A1(n3302), .A2(n3226), .ZN(n3257) );
  INV_X1 U4231 ( .A(n3227), .ZN(n3531) );
  FA_X1 U4232 ( .A(n3230), .B(n3229), .CI(n3228), .CO(n3530), .S(n3191) );
  OAI22_X1 U4233 ( .A1(n4515), .A2(n127), .B1(n3231), .B2(n4498), .ZN(
        \DP/ALU0/N46 ) );
  AOI22_X1 U4234 ( .A1(n2449), .A2(\DP/RegALU2_out[25] ), .B1(
        \DP/RegLMD_out[25] ), .B2(n2448), .ZN(n4461) );
  AOI22_X1 U4235 ( .A1(n3386), .A2(\DP/NPC2[25] ), .B1(n2408), .B2(
        \DP/RegALU1_out[25] ), .ZN(n3233) );
  NAND2_X1 U4236 ( .A1(n2411), .A2(\DP/RegA_out[25] ), .ZN(n3232) );
  OAI211_X1 U4237 ( .C1(n4557), .C2(n2412), .A(n3233), .B(n3232), .ZN(
        \DP/A[25] ) );
  INV_X1 U4238 ( .A(\DP/A[25] ), .ZN(n124) );
  NOR2_X1 U4239 ( .A1(n49), .A2(n3234), .ZN(n3238) );
  OAI22_X1 U4240 ( .A1(n3378), .A2(n3236), .B1(n47), .B2(n3235), .ZN(n3237) );
  AOI211_X1 U4241 ( .C1(n3368), .C2(n3298), .A(n3238), .B(n3237), .ZN(n3273)
         );
  AOI21_X1 U4242 ( .B1(n3392), .B2(n3240), .A(n3239), .ZN(n3242) );
  INV_X1 U4243 ( .A(n3254), .ZN(n3241) );
  NOR2_X1 U4244 ( .A1(n3242), .A2(n3241), .ZN(n3341) );
  INV_X1 U4245 ( .A(n3341), .ZN(n3317) );
  NAND2_X1 U4246 ( .A1(n3242), .A2(n3241), .ZN(n3272) );
  NAND2_X1 U4247 ( .A1(n3317), .A2(n3272), .ZN(n3338) );
  XNOR2_X1 U4248 ( .A(n3273), .B(n3338), .ZN(n3271) );
  XOR2_X1 U4249 ( .A(n3271), .B(n3301), .Z(n3290) );
  AOI21_X1 U4250 ( .B1(n3244), .B2(n3336), .A(n3243), .ZN(n3289) );
  OAI22_X1 U4251 ( .A1(n3246), .A2(n3363), .B1(n3377), .B2(n3245), .ZN(n3247)
         );
  AOI21_X1 U4252 ( .B1(\DP/ALU0/s_A_MULT[11] ), .B2(n3248), .A(n3247), .ZN(
        n3249) );
  OAI21_X1 U4253 ( .B1(n3365), .B2(n3279), .A(n3249), .ZN(n3286) );
  AOI22_X1 U4254 ( .A1(\DP/ALU0/s_A_MULT[12] ), .A2(n3310), .B1(n3348), .B2(
        n3276), .ZN(n3251) );
  NAND2_X1 U4255 ( .A1(n3304), .A2(n3280), .ZN(n3250) );
  OAI211_X1 U4256 ( .C1(n3307), .C2(n3350), .A(n3251), .B(n3250), .ZN(n3285)
         );
  FA_X1 U4257 ( .A(n3254), .B(n3253), .CI(n3252), .CO(n3284), .S(n3244) );
  INV_X1 U4258 ( .A(n3255), .ZN(n3288) );
  INV_X1 U4259 ( .A(n3256), .ZN(n3538) );
  FA_X1 U4260 ( .A(n3259), .B(n3258), .CI(n3257), .CO(n3537), .S(n3227) );
  FA_X1 U4261 ( .A(n3262), .B(n3261), .CI(n3260), .CO(n3536), .S(n3258) );
  NAND2_X1 U4262 ( .A1(n3263), .A2(n2441), .ZN(n3264) );
  OAI21_X1 U4263 ( .B1(n2442), .B2(n124), .A(n3264), .ZN(\DP/ALU0/N47 ) );
  AOI22_X1 U4264 ( .A1(n200), .A2(\DP/RegALU2_out[26] ), .B1(
        \DP/RegLMD_out[26] ), .B2(n2360), .ZN(n4463) );
  AOI22_X1 U4265 ( .A1(n3387), .A2(\DP/RegA_out[26] ), .B1(n2408), .B2(
        \DP/RegALU1_out[26] ), .ZN(n3266) );
  NAND2_X1 U4266 ( .A1(n2410), .A2(\DP/NPC2[26] ), .ZN(n3265) );
  OAI211_X1 U4267 ( .C1(n4463), .C2(n2412), .A(n3266), .B(n3265), .ZN(
        \DP/A[26] ) );
  INV_X1 U4268 ( .A(\DP/A[26] ), .ZN(n121) );
  NAND3_X1 U4269 ( .A1(n51), .A2(n3343), .A3(n3267), .ZN(n3268) );
  OAI21_X1 U4270 ( .B1(n3269), .B2(n3345), .A(n3268), .ZN(n3297) );
  AOI21_X1 U4271 ( .B1(n3270), .B2(n3347), .A(n3297), .ZN(n3316) );
  XNOR2_X1 U4272 ( .A(n3316), .B(n3338), .ZN(n3303) );
  XOR2_X1 U4273 ( .A(n3300), .B(n3303), .Z(n3296) );
  AOI21_X1 U4274 ( .B1(n3271), .B2(n3337), .A(n3302), .ZN(n3295) );
  INV_X1 U4275 ( .A(n3272), .ZN(n3315) );
  AOI21_X1 U4276 ( .B1(n3273), .B2(n3317), .A(n3315), .ZN(n3322) );
  OAI22_X1 U4277 ( .A1(n3311), .A2(n3364), .B1(n3274), .B2(n3363), .ZN(n3275)
         );
  AOI21_X1 U4278 ( .B1(n3277), .B2(n3276), .A(n3275), .ZN(n3278) );
  OAI21_X1 U4279 ( .B1(n3377), .B2(n3279), .A(n3278), .ZN(n3321) );
  AOI22_X1 U4280 ( .A1(n3304), .A2(n3368), .B1(n3348), .B2(n3280), .ZN(n3282)
         );
  NAND2_X1 U4281 ( .A1(\DP/ALU0/s_A_MULT[13] ), .A2(n3310), .ZN(n3281) );
  OAI211_X1 U4282 ( .C1(n49), .C2(n3307), .A(n3282), .B(n3281), .ZN(n3320) );
  INV_X1 U4283 ( .A(n3283), .ZN(n3545) );
  FA_X1 U4284 ( .A(n3286), .B(n3285), .CI(n3284), .CO(n3287), .S(n3255) );
  INV_X1 U4285 ( .A(n3287), .ZN(n3544) );
  FA_X1 U4286 ( .A(n3290), .B(n3289), .CI(n3288), .CO(n3543), .S(n3256) );
  OAI22_X1 U4287 ( .A1(n4515), .A2(n121), .B1(n3291), .B2(n2439), .ZN(
        \DP/ALU0/N48 ) );
  AOI22_X1 U4288 ( .A1(n2449), .A2(\DP/RegALU2_out[27] ), .B1(
        \DP/RegLMD_out[27] ), .B2(n2448), .ZN(n4465) );
  AOI22_X1 U4289 ( .A1(n2411), .A2(\DP/RegA_out[27] ), .B1(n2408), .B2(
        \DP/RegALU1_out[27] ), .ZN(n3293) );
  NAND2_X1 U4290 ( .A1(n2410), .A2(\DP/NPC2[27] ), .ZN(n3292) );
  OAI211_X1 U4291 ( .C1(n4550), .C2(n2412), .A(n3293), .B(n3292), .ZN(
        \DP/A[27] ) );
  INV_X1 U4292 ( .A(\DP/A[27] ), .ZN(n118) );
  FA_X1 U4293 ( .A(n3296), .B(n3295), .CI(n3294), .CO(n3551), .S(n3283) );
  AOI21_X1 U4294 ( .B1(n3392), .B2(n3298), .A(n3297), .ZN(n3339) );
  XOR2_X1 U4295 ( .A(n3339), .B(n3338), .Z(n3335) );
  INV_X1 U4296 ( .A(n3335), .ZN(n3299) );
  AOI22_X1 U4297 ( .A1(n3335), .A2(n3301), .B1(n3300), .B2(n3299), .ZN(n3330)
         );
  AOI21_X1 U4298 ( .B1(n3303), .B2(n3337), .A(n3302), .ZN(n3329) );
  AOI22_X1 U4299 ( .A1(n3305), .A2(n3304), .B1(n3362), .B2(n3368), .ZN(n3306)
         );
  OAI21_X1 U4300 ( .B1(n47), .B2(n3307), .A(n3306), .ZN(n3308) );
  AOI21_X1 U4301 ( .B1(n3310), .B2(n3309), .A(n3308), .ZN(n3334) );
  OAI22_X1 U4302 ( .A1(n3350), .A2(n3364), .B1(n3311), .B2(n3363), .ZN(n3314)
         );
  OAI22_X1 U4303 ( .A1(n3377), .A2(n3312), .B1(n3365), .B2(n3349), .ZN(n3313)
         );
  NOR2_X1 U4304 ( .A1(n3314), .A2(n3313), .ZN(n3333) );
  AOI21_X1 U4305 ( .B1(n3317), .B2(n3316), .A(n3315), .ZN(n3318) );
  INV_X1 U4306 ( .A(n3318), .ZN(n3332) );
  INV_X1 U4307 ( .A(n3319), .ZN(n3328) );
  FA_X1 U4308 ( .A(n3322), .B(n3321), .CI(n3320), .CO(n3549), .S(n3294) );
  XOR2_X1 U4309 ( .A(n3550), .B(n3549), .Z(n3324) );
  NAND2_X1 U4310 ( .A1(n3551), .A2(n3324), .ZN(n3323) );
  OAI211_X1 U4311 ( .C1(n3551), .C2(n3324), .A(n2441), .B(n3323), .ZN(n3325)
         );
  OAI21_X1 U4312 ( .B1(n2443), .B2(n118), .A(n3325), .ZN(\DP/ALU0/N49 ) );
  AOI22_X1 U4314 ( .A1(n3386), .A2(\DP/NPC2[28] ), .B1(n2408), .B2(
        \DP/RegALU1_out[28] ), .ZN(n3327) );
  NAND2_X1 U4315 ( .A1(n2411), .A2(\DP/RegA_out[28] ), .ZN(n3326) );
  INV_X1 U4317 ( .A(\DP/A[28] ), .ZN(n115) );
  FA_X1 U4318 ( .A(n3330), .B(n3329), .CI(n3328), .CO(n3331), .S(n3550) );
  INV_X1 U4319 ( .A(n3331), .ZN(n3558) );
  FA_X1 U4320 ( .A(n3334), .B(n3333), .CI(n3332), .CO(n3557), .S(n3319) );
  NOR2_X1 U4321 ( .A1(n3336), .A2(n3335), .ZN(n3374) );
  INV_X1 U4322 ( .A(n3374), .ZN(n3400) );
  NOR2_X1 U4323 ( .A1(n3339), .A2(n3338), .ZN(n3340) );
  AOI211_X1 U4324 ( .C1(n3339), .C2(n3338), .A(n3340), .B(n3337), .ZN(n3360)
         );
  INV_X1 U4325 ( .A(n3360), .ZN(n3372) );
  NAND2_X1 U4326 ( .A1(n3400), .A2(n3372), .ZN(n3379) );
  NOR2_X1 U4327 ( .A1(n3341), .A2(n3340), .ZN(n3380) );
  NAND3_X1 U4328 ( .A1(n12), .A2(n3343), .A3(n3342), .ZN(n3344) );
  OAI21_X1 U4329 ( .B1(n3346), .B2(n3345), .A(n3344), .ZN(n3361) );
  AOI21_X1 U4330 ( .B1(n3348), .B2(n3347), .A(n3361), .ZN(n3357) );
  NOR2_X1 U4331 ( .A1(n49), .A2(n3364), .ZN(n3352) );
  OAI22_X1 U4332 ( .A1(n3350), .A2(n3363), .B1(n3377), .B2(n3349), .ZN(n3351)
         );
  AOI211_X1 U4333 ( .C1(n3368), .C2(n3376), .A(n3352), .B(n3351), .ZN(n3356)
         );
  XNOR2_X1 U4334 ( .A(n3379), .B(n3358), .ZN(n3556) );
  OAI22_X1 U4335 ( .A1(n2443), .A2(n115), .B1(n3353), .B2(n2439), .ZN(
        \DP/ALU0/N50 ) );
  AOI22_X1 U4336 ( .A1(n2449), .A2(\DP/RegALU2_out[29] ), .B1(
        \DP/RegLMD_out[29] ), .B2(n2448), .ZN(n4469) );
  AOI22_X1 U4337 ( .A1(n3387), .A2(\DP/RegA_out[29] ), .B1(n2408), .B2(
        \DP/RegALU1_out[29] ), .ZN(n3355) );
  NAND2_X1 U4338 ( .A1(n2410), .A2(\DP/NPC2[29] ), .ZN(n3354) );
  OAI211_X1 U4339 ( .C1(n4469), .C2(n2413), .A(n3355), .B(n3354), .ZN(
        \DP/A[29] ) );
  INV_X1 U4340 ( .A(\DP/A[29] ), .ZN(n112) );
  FA_X1 U4341 ( .A(n3380), .B(n3357), .CI(n3356), .CO(n3564), .S(n3358) );
  NOR2_X1 U4342 ( .A1(n3358), .A2(n3379), .ZN(n3359) );
  NOR2_X1 U4343 ( .A1(n3360), .A2(n3359), .ZN(n3563) );
  INV_X1 U4344 ( .A(n3379), .ZN(n3398) );
  AOI21_X1 U4345 ( .B1(n3392), .B2(n3362), .A(n3361), .ZN(n3381) );
  XOR2_X1 U4346 ( .A(n3381), .B(n3380), .Z(n3395) );
  NOR2_X1 U4347 ( .A1(n49), .A2(n3363), .ZN(n3367) );
  OAI22_X1 U4348 ( .A1(n3378), .A2(n3365), .B1(n47), .B2(n3364), .ZN(n3366) );
  AOI211_X1 U4349 ( .C1(n3393), .C2(n3368), .A(n3367), .B(n3366), .ZN(n3383)
         );
  XOR2_X1 U4350 ( .A(n3395), .B(n3383), .Z(n3373) );
  XOR2_X1 U4351 ( .A(n3398), .B(n3373), .Z(n3562) );
  OAI22_X1 U4352 ( .A1(n4515), .A2(n112), .B1(n3369), .B2(n2439), .ZN(
        \DP/ALU0/N51 ) );
  AOI22_X1 U4354 ( .A1(n2411), .A2(\DP/RegA_out[30] ), .B1(n2408), .B2(
        \DP/RegALU1_out[30] ), .ZN(n3371) );
  NAND2_X1 U4355 ( .A1(n2410), .A2(\DP/NPC2[30] ), .ZN(n3370) );
  INV_X1 U4357 ( .A(\DP/A[30] ), .ZN(n109) );
  OAI21_X1 U4358 ( .B1(n3374), .B2(n3373), .A(n3372), .ZN(n3572) );
  AOI21_X1 U4359 ( .B1(n12), .B2(n50), .A(n47), .ZN(n3375) );
  AOI22_X1 U4360 ( .A1(n3392), .A2(n3376), .B1(n48), .B2(n3375), .ZN(n3390) );
  OAI21_X1 U4361 ( .B1(n3378), .B2(n3377), .A(n3390), .ZN(n3394) );
  XOR2_X1 U4362 ( .A(n3395), .B(n3394), .Z(n3399) );
  XNOR2_X1 U4363 ( .A(n3399), .B(n3379), .ZN(n3571) );
  NAND2_X1 U4364 ( .A1(n3381), .A2(n3380), .ZN(n3397) );
  INV_X1 U4365 ( .A(n3397), .ZN(n3382) );
  AOI21_X1 U4366 ( .B1(n3395), .B2(n3383), .A(n3382), .ZN(n3570) );
  NAND2_X1 U4367 ( .A1(n3384), .A2(n2441), .ZN(n3385) );
  OAI21_X1 U4368 ( .B1(n2442), .B2(n109), .A(n3385), .ZN(\DP/ALU0/N52 ) );
  AOI22_X1 U4369 ( .A1(n2449), .A2(\DP/RegALU2_out[31] ), .B1(
        \DP/RegLMD_out[31] ), .B2(n2448), .ZN(n4476) );
  AOI22_X1 U4370 ( .A1(n3386), .A2(\DP/NPC2[31] ), .B1(n2408), .B2(
        \DP/RegALU1_out[31] ), .ZN(n3389) );
  NAND2_X1 U4371 ( .A1(n2411), .A2(\DP/RegA_out[31] ), .ZN(n3388) );
  OAI211_X1 U4372 ( .C1(n4549), .C2(n2413), .A(n3389), .B(n3388), .ZN(
        \DP/A[31] ) );
  INV_X1 U4373 ( .A(\DP/A[31] ), .ZN(n106) );
  INV_X1 U4374 ( .A(n3390), .ZN(n3391) );
  AOI21_X1 U4375 ( .B1(n3393), .B2(n3392), .A(n3391), .ZN(n3405) );
  NAND2_X1 U4376 ( .A1(n3395), .A2(n3394), .ZN(n3396) );
  NAND2_X1 U4377 ( .A1(n3397), .A2(n3396), .ZN(n3403) );
  NAND2_X1 U4378 ( .A1(n3399), .A2(n3398), .ZN(n3401) );
  NAND2_X1 U4379 ( .A1(n3401), .A2(n3400), .ZN(n3402) );
  XNOR2_X1 U4380 ( .A(n3403), .B(n3402), .ZN(n3404) );
  XNOR2_X1 U4381 ( .A(n3405), .B(n3404), .ZN(n3406) );
  OAI22_X1 U4382 ( .A1(n106), .A2(n2443), .B1(n3406), .B2(n2439), .ZN(
        \DP/ALU0/N53 ) );
  NAND3_X1 U4383 ( .A1(n2368), .A2(n2404), .A3(n405), .ZN(n3407) );
  AOI22_X1 U4384 ( .A1(n3569), .A2(\DP/RegIMM_out[0] ), .B1(n2416), .B2(
        DRAM_ADDR[0]), .ZN(n3409) );
  NAND2_X1 U4385 ( .A1(n2414), .A2(\DP/RegB_out[0] ), .ZN(n3408) );
  OAI211_X1 U4386 ( .C1(n4504), .C2(n2418), .A(n3409), .B(n3408), .ZN(
        \DP/B[0] ) );
  AND2_X1 U4387 ( .A1(n3420), .A2(\DP/B[0] ), .ZN(\DP/ALU0/N54 ) );
  AOI22_X1 U4388 ( .A1(n2419), .A2(\DP/RegIMM_out[1] ), .B1(n2415), .B2(
        DRAM_ADDR[1]), .ZN(n3411) );
  NAND2_X1 U4389 ( .A1(n2414), .A2(\DP/RegB_out[1] ), .ZN(n3410) );
  OAI211_X1 U4390 ( .C1(n4502), .C2(n2418), .A(n3411), .B(n3410), .ZN(
        \DP/B[1] ) );
  AND2_X1 U4391 ( .A1(n3420), .A2(\DP/B[1] ), .ZN(\DP/ALU0/N55 ) );
  AOI22_X1 U4392 ( .A1(n3566), .A2(\DP/RegB_out[2] ), .B1(n2416), .B2(
        DRAM_ADDR[2]), .ZN(n3413) );
  NAND2_X1 U4393 ( .A1(n2419), .A2(\DP/RegIMM_out[2] ), .ZN(n3412) );
  OAI211_X1 U4394 ( .C1(n4494), .C2(n2418), .A(n3413), .B(n3412), .ZN(
        \DP/B[2] ) );
  AND2_X1 U4395 ( .A1(n3420), .A2(\DP/B[2] ), .ZN(\DP/ALU0/N56 ) );
  AOI22_X1 U4396 ( .A1(n2419), .A2(\DP/RegIMM_out[3] ), .B1(n2416), .B2(
        DRAM_ADDR[3]), .ZN(n3415) );
  NAND2_X1 U4397 ( .A1(n2414), .A2(\DP/RegB_out[3] ), .ZN(n3414) );
  OAI211_X1 U4398 ( .C1(n4492), .C2(n2418), .A(n3415), .B(n3414), .ZN(
        \DP/B[3] ) );
  AND2_X1 U4399 ( .A1(n3420), .A2(\DP/B[3] ), .ZN(\DP/ALU0/N57 ) );
  AOI22_X1 U4400 ( .A1(n3566), .A2(\DP/RegB_out[4] ), .B1(n2416), .B2(
        DRAM_ADDR[4]), .ZN(n3417) );
  NAND2_X1 U4401 ( .A1(n2419), .A2(\DP/RegIMM_out[4] ), .ZN(n3416) );
  OAI211_X1 U4402 ( .C1(n4561), .C2(n2418), .A(n3417), .B(n3416), .ZN(
        \DP/B[4] ) );
  AND2_X1 U4403 ( .A1(n3420), .A2(\DP/B[4] ), .ZN(\DP/ALU0/N58 ) );
  AOI22_X1 U4404 ( .A1(n3569), .A2(\DP/RegIMM_out[5] ), .B1(n2416), .B2(
        DRAM_ADDR[5]), .ZN(n3419) );
  NAND2_X1 U4405 ( .A1(n2414), .A2(\DP/RegB_out[5] ), .ZN(n3418) );
  OAI211_X1 U4406 ( .C1(n4517), .C2(n2418), .A(n3419), .B(n3418), .ZN(
        \DP/B[5] ) );
  AND2_X1 U4407 ( .A1(n3420), .A2(\DP/B[5] ), .ZN(\DP/ALU0/N59 ) );
  AOI22_X1 U4408 ( .A1(n2419), .A2(\DP/RegIMM_out[6] ), .B1(n2416), .B2(
        DRAM_ADDR[6]), .ZN(n3422) );
  NAND2_X1 U4409 ( .A1(n2414), .A2(\DP/RegB_out[6] ), .ZN(n3421) );
  OAI211_X1 U4410 ( .C1(n4520), .C2(n2418), .A(n3422), .B(n3421), .ZN(
        \DP/B[6] ) );
  INV_X1 U4411 ( .A(\DP/B[6] ), .ZN(n183) );
  OAI22_X1 U4412 ( .A1(n2442), .A2(n183), .B1(n3424), .B2(n3423), .ZN(
        \DP/ALU0/N60 ) );
  AOI22_X1 U4413 ( .A1(n3569), .A2(\DP/RegIMM_out[7] ), .B1(n2416), .B2(
        DRAM_ADDR[7]), .ZN(n3426) );
  NAND2_X1 U4414 ( .A1(n2414), .A2(\DP/RegB_out[7] ), .ZN(n3425) );
  OAI211_X1 U4415 ( .C1(n3657), .C2(n2418), .A(n3426), .B(n3425), .ZN(
        \DP/B[7] ) );
  INV_X1 U4416 ( .A(\DP/B[7] ), .ZN(n179) );
  NAND3_X1 U4417 ( .A1(n2441), .A2(n3428), .A3(n3427), .ZN(n3429) );
  OAI22_X1 U4418 ( .A1(n3430), .A2(n3429), .B1(n2442), .B2(n179), .ZN(
        \DP/ALU0/N61 ) );
  AOI22_X1 U4419 ( .A1(DRAM_ADDR[8]), .A2(n2415), .B1(n2419), .B2(
        \DP/RegIMM_out[8] ), .ZN(n3432) );
  NAND2_X1 U4420 ( .A1(n2414), .A2(\DP/RegB_out[8] ), .ZN(n3431) );
  OAI211_X1 U4421 ( .C1(n4548), .C2(n2418), .A(n3432), .B(n3431), .ZN(
        \DP/B[8] ) );
  INV_X1 U4422 ( .A(\DP/B[8] ), .ZN(n176) );
  NAND3_X1 U4423 ( .A1(n3435), .A2(n3434), .A3(n3433), .ZN(n3436) );
  OAI22_X1 U4424 ( .A1(n4515), .A2(n176), .B1(n3436), .B2(n2439), .ZN(
        \DP/ALU0/N62 ) );
  AOI22_X1 U4425 ( .A1(DRAM_ADDR[9]), .A2(n2415), .B1(n2414), .B2(
        \DP/RegB_out[9] ), .ZN(n3438) );
  NAND2_X1 U4426 ( .A1(n2419), .A2(\DP/RegIMM_out[9] ), .ZN(n3437) );
  OAI211_X1 U4427 ( .C1(n4551), .C2(n2418), .A(n3438), .B(n3437), .ZN(
        \DP/B[9] ) );
  INV_X1 U4428 ( .A(\DP/B[9] ), .ZN(n173) );
  NAND3_X1 U4429 ( .A1(n2440), .A2(n3440), .A3(n3439), .ZN(n3441) );
  OAI21_X1 U4430 ( .B1(n2443), .B2(n173), .A(n3441), .ZN(\DP/ALU0/N63 ) );
  AOI22_X1 U4431 ( .A1(DRAM_ADDR[10]), .A2(n2415), .B1(n2419), .B2(
        \DP/RegIMM_out[10] ), .ZN(n3443) );
  NAND2_X1 U4432 ( .A1(n2414), .A2(\DP/RegB_out[10] ), .ZN(n3442) );
  OAI211_X1 U4433 ( .C1(n4430), .C2(n2418), .A(n3443), .B(n3442), .ZN(
        \DP/B[10] ) );
  INV_X1 U4434 ( .A(\DP/B[10] ), .ZN(n170) );
  NAND3_X1 U4435 ( .A1(n3445), .A2(n2441), .A3(n3444), .ZN(n3446) );
  OAI21_X1 U4436 ( .B1(n2442), .B2(n170), .A(n3446), .ZN(\DP/ALU0/N64 ) );
  AOI22_X1 U4437 ( .A1(n3569), .A2(\DP/RegIMM_out[11] ), .B1(n2416), .B2(
        DRAM_ADDR[11]), .ZN(n3448) );
  NAND2_X1 U4438 ( .A1(n2414), .A2(\DP/RegB_out[11] ), .ZN(n3447) );
  OAI211_X1 U4439 ( .C1(n4565), .C2(n2417), .A(n3448), .B(n3447), .ZN(
        \DP/B[11] ) );
  INV_X1 U4440 ( .A(\DP/B[11] ), .ZN(n167) );
  OR3_X1 U4441 ( .A1(n3450), .A2(n4498), .A3(n3449), .ZN(n3451) );
  OAI21_X1 U4442 ( .B1(n2443), .B2(n167), .A(n3451), .ZN(\DP/ALU0/N65 ) );
  AOI22_X1 U4443 ( .A1(n3566), .A2(\DP/RegB_out[12] ), .B1(n2416), .B2(
        \DP/RegALU1_out[12] ), .ZN(n3453) );
  NAND2_X1 U4444 ( .A1(n2419), .A2(\DP/RegIMM_out[12] ), .ZN(n3452) );
  INV_X1 U4446 ( .A(\DP/B[12] ), .ZN(n164) );
  OR2_X1 U4447 ( .A1(n3455), .A2(n3454), .ZN(n3456) );
  OAI22_X1 U4448 ( .A1(n2443), .A2(n164), .B1(n3456), .B2(n2439), .ZN(
        \DP/ALU0/N66 ) );
  AOI22_X1 U4449 ( .A1(n3569), .A2(\DP/RegIMM_out[13] ), .B1(n2416), .B2(
        \DP/RegALU1_out[13] ), .ZN(n3458) );
  NAND2_X1 U4450 ( .A1(n2414), .A2(\DP/RegB_out[13] ), .ZN(n3457) );
  OAI211_X1 U4451 ( .C1(n4556), .C2(n2417), .A(n3458), .B(n3457), .ZN(
        \DP/B[13] ) );
  INV_X1 U4452 ( .A(\DP/B[13] ), .ZN(n161) );
  OR2_X1 U4453 ( .A1(n3460), .A2(n3459), .ZN(n3461) );
  OAI22_X1 U4454 ( .A1(n4515), .A2(n161), .B1(n3461), .B2(n2439), .ZN(
        \DP/ALU0/N67 ) );
  AOI22_X1 U4455 ( .A1(n3566), .A2(\DP/RegB_out[14] ), .B1(n2416), .B2(
        \DP/RegALU1_out[14] ), .ZN(n3463) );
  NAND2_X1 U4456 ( .A1(n2419), .A2(\DP/RegIMM_out[14] ), .ZN(n3462) );
  OAI211_X1 U4457 ( .C1(n4542), .C2(n2418), .A(n3463), .B(n3462), .ZN(
        \DP/B[14] ) );
  INV_X1 U4458 ( .A(\DP/B[14] ), .ZN(n158) );
  FA_X1 U4459 ( .A(n3466), .B(n3465), .CI(n3464), .CO(n3467), .S(n2832) );
  OAI22_X1 U4460 ( .A1(n2442), .A2(n158), .B1(n3467), .B2(n2439), .ZN(
        \DP/ALU0/N68 ) );
  AOI22_X1 U4461 ( .A1(n3569), .A2(\DP/RegIMM_out[15] ), .B1(n2416), .B2(
        \DP/RegALU1_out[15] ), .ZN(n3469) );
  NAND2_X1 U4462 ( .A1(n2414), .A2(\DP/RegB_out[15] ), .ZN(n3468) );
  OAI211_X1 U4463 ( .C1(n4440), .C2(n2417), .A(n3469), .B(n3468), .ZN(
        \DP/B[15] ) );
  INV_X1 U4464 ( .A(\DP/B[15] ), .ZN(n155) );
  FA_X1 U4465 ( .A(n3472), .B(n3471), .CI(n3470), .CO(n3473), .S(n2865) );
  OAI22_X1 U4466 ( .A1(n2443), .A2(n155), .B1(n3473), .B2(n2439), .ZN(
        \DP/ALU0/N69 ) );
  AOI22_X1 U4467 ( .A1(n3566), .A2(\DP/RegB_out[16] ), .B1(n2416), .B2(
        \DP/RegALU1_out[16] ), .ZN(n3474) );
  OAI21_X1 U4468 ( .B1(n4442), .B2(n2418), .A(n3474), .ZN(n3475) );
  AOI21_X1 U4469 ( .B1(n3569), .B2(\DP/RegIMM_out[16] ), .A(n3475), .ZN(n152)
         );
  FA_X1 U4470 ( .A(n3478), .B(n3477), .CI(n3476), .CO(n3479), .S(n2902) );
  OAI22_X1 U4471 ( .A1(n2443), .A2(n152), .B1(n3479), .B2(n2439), .ZN(
        \DP/ALU0/N70 ) );
  AOI22_X1 U4472 ( .A1(n3569), .A2(\DP/RegIMM_out[17] ), .B1(n2415), .B2(
        \DP/RegALU1_out[17] ), .ZN(n3480) );
  OAI21_X1 U4473 ( .B1(n4444), .B2(n2418), .A(n3480), .ZN(n3481) );
  AOI21_X1 U4474 ( .B1(n3566), .B2(\DP/RegB_out[17] ), .A(n3481), .ZN(n149) );
  FA_X1 U4475 ( .A(n3484), .B(n3483), .CI(n3482), .CO(n3485), .S(n2942) );
  OAI22_X1 U4476 ( .A1(n4515), .A2(n149), .B1(n3485), .B2(n2439), .ZN(
        \DP/ALU0/N71 ) );
  AOI22_X1 U4477 ( .A1(n2419), .A2(\DP/RegIMM_out[18] ), .B1(n2416), .B2(
        \DP/RegALU1_out[18] ), .ZN(n3486) );
  OAI21_X1 U4478 ( .B1(n4756), .B2(n2417), .A(n3486), .ZN(n3487) );
  AOI21_X1 U4479 ( .B1(n2414), .B2(\DP/RegB_out[18] ), .A(n3487), .ZN(n146) );
  FA_X1 U4480 ( .A(n3490), .B(n3489), .CI(n3488), .CO(n3491), .S(n2981) );
  OAI22_X1 U4481 ( .A1(n2442), .A2(n146), .B1(n3491), .B2(n2439), .ZN(
        \DP/ALU0/N72 ) );
  AOI22_X1 U4482 ( .A1(n3566), .A2(\DP/RegB_out[19] ), .B1(n2415), .B2(
        \DP/RegALU1_out[19] ), .ZN(n3492) );
  OAI21_X1 U4483 ( .B1(n4448), .B2(n2417), .A(n3492), .ZN(n3493) );
  AOI21_X1 U4484 ( .B1(n2419), .B2(\DP/RegIMM_out[19] ), .A(n3493), .ZN(n143)
         );
  FA_X1 U4485 ( .A(n3496), .B(n3495), .CI(n3494), .CO(n3497), .S(n3019) );
  OAI22_X1 U4486 ( .A1(n4515), .A2(n143), .B1(n3497), .B2(n4498), .ZN(
        \DP/ALU0/N73 ) );
  AOI22_X1 U4487 ( .A1(n3569), .A2(\DP/RegIMM_out[20] ), .B1(n2416), .B2(
        \DP/RegALU1_out[20] ), .ZN(n3498) );
  OAI21_X1 U4488 ( .B1(n4450), .B2(n2417), .A(n3498), .ZN(n3499) );
  AOI21_X1 U4489 ( .B1(n2414), .B2(\DP/RegB_out[20] ), .A(n3499), .ZN(n140) );
  FA_X1 U4490 ( .A(n3502), .B(n3501), .CI(n3500), .CO(n3503), .S(n3059) );
  OAI22_X1 U4491 ( .A1(n4515), .A2(n140), .B1(n3503), .B2(n4498), .ZN(
        \DP/ALU0/N74 ) );
  AOI22_X1 U4492 ( .A1(n3569), .A2(\DP/RegIMM_out[21] ), .B1(n2415), .B2(
        \DP/RegALU1_out[21] ), .ZN(n3504) );
  OAI21_X1 U4493 ( .B1(n4554), .B2(n2417), .A(n3504), .ZN(n3505) );
  AOI21_X1 U4494 ( .B1(n3566), .B2(\DP/RegB_out[21] ), .A(n3505), .ZN(n137) );
  FA_X1 U4495 ( .A(n3508), .B(n3507), .CI(n3506), .CO(n3509), .S(n3097) );
  OAI22_X1 U4496 ( .A1(n4515), .A2(n137), .B1(n3509), .B2(n2439), .ZN(
        \DP/ALU0/N75 ) );
  AOI22_X1 U4497 ( .A1(n3566), .A2(\DP/RegB_out[22] ), .B1(n2415), .B2(
        \DP/RegALU1_out[22] ), .ZN(n3510) );
  OAI21_X1 U4498 ( .B1(n4454), .B2(n2417), .A(n3510), .ZN(n3511) );
  AOI21_X1 U4499 ( .B1(n2419), .B2(\DP/RegIMM_out[22] ), .A(n3511), .ZN(n134)
         );
  FA_X1 U4500 ( .A(n3514), .B(n3513), .CI(n3512), .CO(n3515), .S(n3138) );
  OAI22_X1 U4501 ( .A1(n4515), .A2(n134), .B1(n3515), .B2(n2439), .ZN(
        \DP/ALU0/N76 ) );
  AOI22_X1 U4502 ( .A1(n3566), .A2(\DP/RegB_out[23] ), .B1(n2384), .B2(n4455), 
        .ZN(n3516) );
  OAI21_X1 U4503 ( .B1(n2361), .B2(n2366), .A(n3516), .ZN(n3517) );
  AOI21_X1 U4504 ( .B1(n2419), .B2(\DP/RegIMM_out[23] ), .A(n3517), .ZN(n131)
         );
  FA_X1 U4505 ( .A(n3520), .B(n3519), .CI(n3518), .CO(n3521), .S(n3169) );
  OAI22_X1 U4506 ( .A1(n4515), .A2(n131), .B1(n3521), .B2(n4498), .ZN(
        \DP/ALU0/N77 ) );
  AOI22_X1 U4507 ( .A1(n2414), .A2(\DP/RegB_out[24] ), .B1(n2384), .B2(n4457), 
        .ZN(n3522) );
  OAI21_X1 U4508 ( .B1(n2361), .B2(n2393), .A(n3522), .ZN(n3523) );
  AOI21_X1 U4509 ( .B1(n2419), .B2(\DP/RegIMM_out[24] ), .A(n3523), .ZN(n128)
         );
  FA_X1 U4510 ( .A(n3526), .B(n3525), .CI(n3524), .CO(n3527), .S(n3199) );
  OAI22_X1 U4511 ( .A1(n4515), .A2(n128), .B1(n3527), .B2(n2439), .ZN(
        \DP/ALU0/N78 ) );
  AOI22_X1 U4512 ( .A1(n3569), .A2(\DP/RegIMM_out[25] ), .B1(n2415), .B2(
        \DP/RegALU1_out[25] ), .ZN(n3528) );
  OAI21_X1 U4513 ( .B1(n4557), .B2(n2417), .A(n3528), .ZN(n3529) );
  AOI21_X1 U4514 ( .B1(n2414), .B2(\DP/RegB_out[25] ), .A(n3529), .ZN(n125) );
  FA_X1 U4515 ( .A(n3532), .B(n3531), .CI(n3530), .CO(n3533), .S(n3231) );
  OAI22_X1 U4516 ( .A1(n4515), .A2(n125), .B1(n3533), .B2(n4498), .ZN(
        \DP/ALU0/N79 ) );
  AOI22_X1 U4517 ( .A1(n2414), .A2(\DP/RegB_out[26] ), .B1(n2415), .B2(
        \DP/RegALU1_out[26] ), .ZN(n3534) );
  OAI21_X1 U4518 ( .B1(n4463), .B2(n2417), .A(n3534), .ZN(n3535) );
  AOI21_X1 U4519 ( .B1(n2419), .B2(\DP/RegIMM_out[26] ), .A(n3535), .ZN(n122)
         );
  FA_X1 U4520 ( .A(n3538), .B(n3537), .CI(n3536), .CO(n3539), .S(n3263) );
  NAND2_X1 U4521 ( .A1(n3539), .A2(n2441), .ZN(n3540) );
  OAI21_X1 U4522 ( .B1(n2443), .B2(n122), .A(n3540), .ZN(\DP/ALU0/N80 ) );
  AOI22_X1 U4523 ( .A1(n2414), .A2(\DP/RegB_out[27] ), .B1(n2415), .B2(
        \DP/RegALU1_out[27] ), .ZN(n3541) );
  OAI21_X1 U4524 ( .B1(n4550), .B2(n2417), .A(n3541), .ZN(n3542) );
  AOI21_X1 U4525 ( .B1(n2419), .B2(\DP/RegIMM_out[27] ), .A(n3542), .ZN(n119)
         );
  FA_X1 U4526 ( .A(n3545), .B(n3544), .CI(n3543), .CO(n3546), .S(n3291) );
  OAI22_X1 U4527 ( .A1(n2443), .A2(n119), .B1(n3546), .B2(n2439), .ZN(
        \DP/ALU0/N81 ) );
  AOI22_X1 U4528 ( .A1(\DP/RegALU1_out[28] ), .A2(n2415), .B1(n2419), .B2(
        \DP/RegIMM_out[28] ), .ZN(n3547) );
  AOI21_X1 U4530 ( .B1(n3566), .B2(\DP/RegB_out[28] ), .A(n3548), .ZN(n116) );
  AOI21_X1 U4531 ( .B1(n3550), .B2(n3551), .A(n3549), .ZN(n3553) );
  OAI21_X1 U4532 ( .B1(n3551), .B2(n3550), .A(n2441), .ZN(n3552) );
  OAI22_X1 U4533 ( .A1(n3553), .A2(n3552), .B1(n2442), .B2(n116), .ZN(
        \DP/ALU0/N82 ) );
  AOI22_X1 U4534 ( .A1(\DP/RegALU1_out[29] ), .A2(n2415), .B1(n2414), .B2(
        \DP/RegB_out[29] ), .ZN(n3554) );
  OAI21_X1 U4535 ( .B1(n4469), .B2(n2417), .A(n3554), .ZN(n3555) );
  AOI21_X1 U4536 ( .B1(n2419), .B2(\DP/RegIMM_out[29] ), .A(n3555), .ZN(n113)
         );
  FA_X1 U4537 ( .A(n3558), .B(n3557), .CI(n3556), .CO(n3559), .S(n3353) );
  OAI22_X1 U4538 ( .A1(n4515), .A2(n113), .B1(n3559), .B2(n4498), .ZN(
        \DP/ALU0/N83 ) );
  AOI22_X1 U4539 ( .A1(\DP/RegALU1_out[30] ), .A2(n2415), .B1(n2414), .B2(
        \DP/RegB_out[30] ), .ZN(n3560) );
  AOI21_X1 U4541 ( .B1(n2419), .B2(\DP/RegIMM_out[30] ), .A(n3561), .ZN(n110)
         );
  FA_X1 U4542 ( .A(n3564), .B(n3563), .CI(n3562), .CO(n3565), .S(n3369) );
  OAI22_X1 U4543 ( .A1(n2443), .A2(n110), .B1(n3565), .B2(n2439), .ZN(
        \DP/ALU0/N84 ) );
  AOI22_X1 U4544 ( .A1(\DP/RegALU1_out[31] ), .A2(n2415), .B1(n2414), .B2(
        \DP/RegB_out[31] ), .ZN(n3567) );
  OAI21_X1 U4545 ( .B1(n4549), .B2(n2417), .A(n3567), .ZN(n3568) );
  AOI21_X1 U4546 ( .B1(n2419), .B2(\DP/RegIMM_out[31] ), .A(n3568), .ZN(n107)
         );
  FA_X1 U4547 ( .A(n3572), .B(n3571), .CI(n3570), .CO(n3573), .S(n3384) );
  NAND2_X1 U4548 ( .A1(n3573), .A2(n2441), .ZN(n3574) );
  OAI21_X1 U4549 ( .B1(n2443), .B2(n107), .A(n3574), .ZN(\DP/ALU0/N85 ) );
  NOR4_X1 U4551 ( .A1(w_ALU_OPCODE[3]), .A2(w_ALU_OPCODE[4]), .A3(n2362), .A4(
        n2373), .ZN(\DP/ALU0/N88 ) );
  OAI21_X1 U4552 ( .B1(n218), .B2(n3577), .A(n4623), .ZN(n3578) );
  INV_X1 U4553 ( .A(n3578), .ZN(\DP/ALU0/N89 ) );
  NAND2_X1 U4555 ( .A1(n4275), .A2(n208), .ZN(\DP/FFDBRANCH/N2 ) );
  NOR2_X1 U4556 ( .A1(n2460), .A2(n2392), .ZN(\DP/FFDJL1/N3 ) );
  NOR2_X1 U4557 ( .A1(n207), .A2(n2460), .ZN(\DP/FFDJREG/N3 ) );
  NAND4_X1 U4559 ( .A1(n4480), .A2(n4485), .A3(n3657), .A4(n4440), .ZN(n3587)
         );
  NAND4_X1 U4560 ( .A1(n4454), .A2(n4452), .A3(n4450), .A4(n4448), .ZN(n3579)
         );
  NAND4_X1 U4562 ( .A1(n4492), .A2(n4494), .A3(n4502), .A4(n4504), .ZN(n3583)
         );
  NAND4_X1 U4563 ( .A1(n4476), .A2(n4517), .A3(n4520), .A4(n4506), .ZN(n3582)
         );
  NAND3_X1 U4569 ( .A1(\DP/FwdC[1] ), .A2(n407), .A3(n406), .ZN(n3654) );
  NOR4_X1 U4570 ( .A1(\DP/RegALU1_out[18] ), .A2(\DP/RegALU1_out[17] ), .A3(
        \DP/RegALU1_out[16] ), .A4(\DP/RegALU1_out[15] ), .ZN(n3592) );
  NOR4_X1 U4571 ( .A1(\DP/RegALU1_out[22] ), .A2(\DP/RegALU1_out[21] ), .A3(
        \DP/RegALU1_out[20] ), .A4(\DP/RegALU1_out[19] ), .ZN(n3591) );
  NOR4_X1 U4572 ( .A1(DRAM_ADDR[10]), .A2(DRAM_ADDR[8]), .A3(DRAM_ADDR[9]), 
        .A4(DRAM_ADDR[7]), .ZN(n3590) );
  NOR4_X1 U4573 ( .A1(DRAM_ADDR[11]), .A2(\DP/RegALU1_out[14] ), .A3(
        \DP/RegALU1_out[13] ), .A4(\DP/RegALU1_out[12] ), .ZN(n3589) );
  NAND4_X1 U4574 ( .A1(n3592), .A2(n3591), .A3(n3590), .A4(n3589), .ZN(n3598)
         );
  NOR4_X1 U4575 ( .A1(\DP/RegALU1_out[30] ), .A2(DRAM_ADDR[5]), .A3(
        DRAM_ADDR[3]), .A4(DRAM_ADDR[1]), .ZN(n3596) );
  NOR4_X1 U4576 ( .A1(\DP/RegALU1_out[31] ), .A2(DRAM_ADDR[6]), .A3(
        DRAM_ADDR[4]), .A4(DRAM_ADDR[2]), .ZN(n3595) );
  NOR4_X1 U4577 ( .A1(\DP/RegALU1_out[26] ), .A2(\DP/RegALU1_out[25] ), .A3(
        \DP/RegALU1_out[24] ), .A4(\DP/RegALU1_out[23] ), .ZN(n3594) );
  NOR4_X1 U4578 ( .A1(\DP/RegALU1_out[29] ), .A2(\DP/RegALU1_out[28] ), .A3(
        \DP/RegALU1_out[27] ), .A4(DRAM_ADDR[0]), .ZN(n3593) );
  NAND4_X1 U4579 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(n3597)
         );
  NOR3_X1 U4580 ( .A1(\DP/FwdC[1] ), .A2(n407), .A3(n2370), .ZN(n3690) );
  OAI21_X1 U4581 ( .B1(n3598), .B2(n3597), .A(n2420), .ZN(n3610) );
  NOR4_X1 U4582 ( .A1(\DP/RegA_out[18] ), .A2(\DP/RegA_out[17] ), .A3(
        \DP/RegA_out[16] ), .A4(\DP/RegA_out[15] ), .ZN(n3602) );
  NOR4_X1 U4583 ( .A1(\DP/RegA_out[22] ), .A2(\DP/RegA_out[21] ), .A3(
        \DP/RegA_out[20] ), .A4(\DP/RegA_out[19] ), .ZN(n3601) );
  NOR4_X1 U4584 ( .A1(\DP/RegA_out[10] ), .A2(\DP/RegA_out[8] ), .A3(
        \DP/RegA_out[9] ), .A4(\DP/RegA_out[7] ), .ZN(n3600) );
  NOR4_X1 U4585 ( .A1(\DP/RegA_out[14] ), .A2(\DP/RegA_out[13] ), .A3(
        \DP/RegA_out[12] ), .A4(\DP/RegA_out[11] ), .ZN(n3599) );
  NAND4_X1 U4586 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3608)
         );
  NOR4_X1 U4587 ( .A1(\DP/RegA_out[5] ), .A2(\DP/RegA_out[3] ), .A3(
        \DP/RegA_out[1] ), .A4(\DP/RegA_out[30] ), .ZN(n3606) );
  NOR4_X1 U4588 ( .A1(\DP/RegA_out[31] ), .A2(\DP/RegA_out[6] ), .A3(
        \DP/RegA_out[4] ), .A4(\DP/RegA_out[2] ), .ZN(n3605) );
  NOR4_X1 U4589 ( .A1(\DP/RegA_out[26] ), .A2(\DP/RegA_out[25] ), .A3(
        \DP/RegA_out[24] ), .A4(\DP/RegA_out[23] ), .ZN(n3604) );
  NOR4_X1 U4590 ( .A1(\DP/RegA_out[0] ), .A2(\DP/RegA_out[29] ), .A3(
        \DP/RegA_out[28] ), .A4(\DP/RegA_out[27] ), .ZN(n3603) );
  NAND4_X1 U4591 ( .A1(n3606), .A2(n3605), .A3(n3604), .A4(n3603), .ZN(n3607)
         );
  NOR3_X1 U4592 ( .A1(\DP/FwdC[1] ), .A2(n406), .A3(n2398), .ZN(n3655) );
  OAI21_X1 U4593 ( .B1(n3608), .B2(n3607), .A(n3655), .ZN(n3609) );
  NAND2_X1 U4598 ( .A1(n3615), .A2(RST), .ZN(\DP/RegNPC1/N2 ) );
  NOR4_X1 U4607 ( .A1(\DP/RD2[1] ), .A2(\DP/RD2[0] ), .A3(n2365), .A4(n2385), 
        .ZN(n3618) );
  AOI21_X1 U4608 ( .B1(n3618), .B2(n2367), .A(n2395), .ZN(n4247) );
  AOI21_X1 U4610 ( .B1(n4421), .B2(\DP/RD2[2] ), .A(n3620), .ZN(n3621) );
  OAI221_X1 U4611 ( .B1(n97), .B2(n401), .C1(n4424), .C2(n2365), .A(n3621), 
        .ZN(n4262) );
  NOR2_X1 U4612 ( .A1(n2460), .A2(n4262), .ZN(\DP/FFDFD/N3 ) );
  NAND2_X1 U4613 ( .A1(RST), .A2(n2392), .ZN(\DP/RegNPC2/N2 ) );
  AND2_X1 U4615 ( .A1(RST), .A2(\DP/JL1 ), .ZN(\DP/FFDJL2/N3 ) );
  NAND2_X1 U4616 ( .A1(n4275), .A2(n207), .ZN(\DP/RegA1/N2 ) );
  NAND2_X1 U4617 ( .A1(n2459), .A2(\DP/NPC_out[0] ), .ZN(n3623) );
  NAND2_X1 U4618 ( .A1(n2459), .A2(\DP/NPC_out[10] ), .ZN(n3624) );
  NAND2_X1 U4619 ( .A1(n2458), .A2(\DP/NPC_out[11] ), .ZN(n3625) );
  NAND2_X1 U4620 ( .A1(n2458), .A2(\DP/NPC_out[12] ), .ZN(n3626) );
  NAND2_X1 U4622 ( .A1(n2458), .A2(\DP/NPC_out[13] ), .ZN(n3627) );
  NAND2_X1 U4624 ( .A1(n2459), .A2(\DP/NPC_out[14] ), .ZN(n3628) );
  NAND2_X1 U4626 ( .A1(n2458), .A2(\DP/NPC_out[15] ), .ZN(n3629) );
  NAND2_X1 U4628 ( .A1(n2458), .A2(\DP/NPC_out[16] ), .ZN(n3630) );
  NAND2_X1 U4630 ( .A1(n2458), .A2(\DP/NPC_out[17] ), .ZN(n3631) );
  NAND2_X1 U4632 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[18] ), .ZN(n3632) );
  NAND2_X1 U4635 ( .A1(n2458), .A2(\DP/NPC_out[1] ), .ZN(n3634) );
  NAND2_X1 U4637 ( .A1(n2458), .A2(\DP/NPC_out[20] ), .ZN(n3635) );
  NAND2_X1 U4638 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[21] ), .ZN(n3636) );
  NAND2_X1 U4640 ( .A1(n2459), .A2(\DP/NPC_out[22] ), .ZN(n3637) );
  MUX2_X1 U4642 ( .A(n4455), .B(\DP/NPC_out[23] ), .S(\DP/JL2 ), .Z(
        \DP/RF_DATA[23] ) );
  MUX2_X1 U4643 ( .A(n4457), .B(\DP/NPC_out[24] ), .S(\DP/JL2 ), .Z(
        \DP/RF_DATA[24] ) );
  NAND2_X1 U4644 ( .A1(n2458), .A2(\DP/NPC_out[25] ), .ZN(n3638) );
  NAND2_X1 U4645 ( .A1(n2458), .A2(\DP/NPC_out[26] ), .ZN(n3639) );
  NAND2_X1 U4646 ( .A1(n2458), .A2(\DP/NPC_out[27] ), .ZN(n3640) );
  NAND2_X1 U4647 ( .A1(n2458), .A2(\DP/NPC_out[28] ), .ZN(n3641) );
  NAND2_X1 U4649 ( .A1(n2458), .A2(\DP/NPC_out[29] ), .ZN(n3642) );
  NAND2_X1 U4651 ( .A1(n2458), .A2(\DP/NPC_out[2] ), .ZN(n3643) );
  NAND2_X1 U4653 ( .A1(n2458), .A2(\DP/NPC_out[30] ), .ZN(n3644) );
  NAND2_X1 U4655 ( .A1(n2459), .A2(\DP/NPC_out[31] ), .ZN(n3645) );
  NAND2_X1 U4657 ( .A1(n2459), .A2(\DP/NPC_out[3] ), .ZN(n3646) );
  NAND2_X1 U4659 ( .A1(n2459), .A2(\DP/NPC_out[4] ), .ZN(n3647) );
  NAND2_X1 U4661 ( .A1(n2459), .A2(\DP/NPC_out[5] ), .ZN(n3648) );
  NAND2_X1 U4663 ( .A1(n2459), .A2(\DP/NPC_out[6] ), .ZN(n3649) );
  NAND2_X1 U4667 ( .A1(n2459), .A2(\DP/NPC_out[8] ), .ZN(n3650) );
  NAND2_X1 U4669 ( .A1(n2459), .A2(\DP/NPC_out[9] ), .ZN(n3651) );
  AND2_X1 U4671 ( .A1(RST), .A2(\DP/RegA_in[7] ), .ZN(\DP/RegA/N10 ) );
  AND2_X1 U4672 ( .A1(RST), .A2(\DP/RegA_in[8] ), .ZN(\DP/RegA/N11 ) );
  AND2_X1 U4673 ( .A1(RST), .A2(\DP/RegA_in[9] ), .ZN(\DP/RegA/N12 ) );
  AND2_X1 U4674 ( .A1(RST), .A2(\DP/RegA_in[10] ), .ZN(\DP/RegA/N13 ) );
  AND2_X1 U4675 ( .A1(RST), .A2(\DP/RegA_in[11] ), .ZN(\DP/RegA/N14 ) );
  AND2_X1 U4676 ( .A1(RST), .A2(\DP/RegA_in[12] ), .ZN(\DP/RegA/N15 ) );
  AND2_X1 U4677 ( .A1(RST), .A2(\DP/RegA_in[13] ), .ZN(\DP/RegA/N16 ) );
  AND2_X1 U4678 ( .A1(RST), .A2(\DP/RegA_in[14] ), .ZN(\DP/RegA/N17 ) );
  AND2_X1 U4679 ( .A1(RST), .A2(\DP/RegA_in[15] ), .ZN(\DP/RegA/N18 ) );
  AND2_X1 U4680 ( .A1(RST), .A2(\DP/RegA_in[16] ), .ZN(\DP/RegA/N19 ) );
  NAND2_X1 U4681 ( .A1(n3653), .A2(n3652), .ZN(w_RF_RD1) );
  AND2_X1 U4683 ( .A1(RST), .A2(\DP/RegA_in[17] ), .ZN(\DP/RegA/N20 ) );
  AND2_X1 U4684 ( .A1(RST), .A2(\DP/RegA_in[18] ), .ZN(\DP/RegA/N21 ) );
  AND2_X1 U4685 ( .A1(RST), .A2(\DP/RegA_in[19] ), .ZN(\DP/RegA/N22 ) );
  AND2_X1 U4686 ( .A1(RST), .A2(\DP/RegA_in[20] ), .ZN(\DP/RegA/N23 ) );
  AND2_X1 U4687 ( .A1(RST), .A2(\DP/RegA_in[21] ), .ZN(\DP/RegA/N24 ) );
  AND2_X1 U4688 ( .A1(RST), .A2(\DP/RegA_in[22] ), .ZN(\DP/RegA/N25 ) );
  AND2_X1 U4689 ( .A1(RST), .A2(\DP/RegA_in[23] ), .ZN(\DP/RegA/N26 ) );
  AND2_X1 U4690 ( .A1(RST), .A2(\DP/RegA_in[24] ), .ZN(\DP/RegA/N27 ) );
  AND2_X1 U4691 ( .A1(RST), .A2(\DP/RegA_in[25] ), .ZN(\DP/RegA/N28 ) );
  AND2_X1 U4692 ( .A1(RST), .A2(\DP/RegA_in[26] ), .ZN(\DP/RegA/N29 ) );
  AND2_X1 U4693 ( .A1(RST), .A2(\DP/RegA_in[0] ), .ZN(\DP/RegA/N3 ) );
  AND2_X1 U4694 ( .A1(RST), .A2(\DP/RegA_in[27] ), .ZN(\DP/RegA/N30 ) );
  AND2_X1 U4695 ( .A1(RST), .A2(\DP/RegA_in[28] ), .ZN(\DP/RegA/N31 ) );
  AND2_X1 U4696 ( .A1(RST), .A2(\DP/RegA_in[29] ), .ZN(\DP/RegA/N32 ) );
  AND2_X1 U4697 ( .A1(RST), .A2(\DP/RegA_in[30] ), .ZN(\DP/RegA/N33 ) );
  AND2_X1 U4698 ( .A1(RST), .A2(\DP/RegA_in[31] ), .ZN(\DP/RegA/N34 ) );
  AND2_X1 U4699 ( .A1(RST), .A2(\DP/RegA_in[1] ), .ZN(\DP/RegA/N4 ) );
  AND2_X1 U4700 ( .A1(RST), .A2(\DP/RegA_in[2] ), .ZN(\DP/RegA/N5 ) );
  AND2_X1 U4701 ( .A1(RST), .A2(\DP/RegA_in[3] ), .ZN(\DP/RegA/N6 ) );
  AND2_X1 U4702 ( .A1(RST), .A2(\DP/RegA_in[4] ), .ZN(\DP/RegA/N7 ) );
  AND2_X1 U4703 ( .A1(RST), .A2(\DP/RegA_in[5] ), .ZN(\DP/RegA/N8 ) );
  AND2_X1 U4704 ( .A1(RST), .A2(\DP/RegA_in[6] ), .ZN(\DP/RegA/N9 ) );
  AOI22_X1 U4705 ( .A1(n2420), .A2(\DP/RegALU2/N10 ), .B1(\DP/RegA_out[7] ), 
        .B2(n3691), .ZN(n3656) );
  OAI21_X1 U4706 ( .B1(n3657), .B2(n2423), .A(n3656), .ZN(\DP/RegA1/N10 ) );
  AOI22_X1 U4707 ( .A1(\DP/RegA_out[8] ), .A2(n2422), .B1(n2421), .B2(
        \DP/RegALU2/N11 ), .ZN(n3658) );
  OAI21_X1 U4708 ( .B1(n4548), .B2(n3693), .A(n3658), .ZN(\DP/RegA1/N11 ) );
  AOI22_X1 U4709 ( .A1(\DP/RegA_out[9] ), .A2(n3691), .B1(n2421), .B2(
        \DP/RegALU2/N12 ), .ZN(n3659) );
  OAI21_X1 U4710 ( .B1(n4551), .B2(n2423), .A(n3659), .ZN(\DP/RegA1/N12 ) );
  AOI22_X1 U4711 ( .A1(\DP/RegA_out[10] ), .A2(n2422), .B1(\DP/RegALU2/N13 ), 
        .B2(n2420), .ZN(n3660) );
  OAI21_X1 U4712 ( .B1(n4430), .B2(n3693), .A(n3660), .ZN(\DP/RegA1/N13 ) );
  AOI22_X1 U4713 ( .A1(\DP/RegALU2/N14 ), .A2(n2421), .B1(\DP/RegA_out[11] ), 
        .B2(n2422), .ZN(n3661) );
  OAI21_X1 U4714 ( .B1(n4565), .B2(n2423), .A(n3661), .ZN(\DP/RegA1/N14 ) );
  AOI22_X1 U4715 ( .A1(\DP/RegALU2/N15 ), .A2(n2421), .B1(\DP/RegA_out[12] ), 
        .B2(n2422), .ZN(n3662) );
  AOI22_X1 U4717 ( .A1(\DP/RegALU2/N16 ), .A2(n2421), .B1(\DP/RegA_out[13] ), 
        .B2(n2422), .ZN(n3663) );
  OAI21_X1 U4718 ( .B1(n4556), .B2(n3693), .A(n3663), .ZN(\DP/RegA1/N16 ) );
  AOI22_X1 U4719 ( .A1(\DP/RegALU2/N17 ), .A2(n3690), .B1(\DP/RegA_out[14] ), 
        .B2(n2422), .ZN(n3664) );
  OAI21_X1 U4720 ( .B1(n4438), .B2(n3693), .A(n3664), .ZN(\DP/RegA1/N17 ) );
  AOI22_X1 U4721 ( .A1(\DP/RegALU2/N18 ), .A2(n3690), .B1(\DP/RegA_out[15] ), 
        .B2(n2422), .ZN(n3665) );
  OAI21_X1 U4722 ( .B1(n4440), .B2(n3693), .A(n3665), .ZN(\DP/RegA1/N18 ) );
  AOI22_X1 U4723 ( .A1(\DP/RegALU2/N19 ), .A2(n3690), .B1(\DP/RegA_out[16] ), 
        .B2(n2422), .ZN(n3666) );
  OAI21_X1 U4724 ( .B1(n4442), .B2(n3693), .A(n3666), .ZN(\DP/RegA1/N19 ) );
  AOI22_X1 U4725 ( .A1(\DP/RegALU2/N20 ), .A2(n3690), .B1(\DP/RegA_out[17] ), 
        .B2(n2422), .ZN(n3667) );
  OAI21_X1 U4726 ( .B1(n4444), .B2(n3693), .A(n3667), .ZN(\DP/RegA1/N20 ) );
  AOI22_X1 U4727 ( .A1(\DP/RegALU2/N21 ), .A2(n3690), .B1(\DP/RegA_out[18] ), 
        .B2(n2422), .ZN(n3668) );
  OAI21_X1 U4728 ( .B1(n4446), .B2(n3693), .A(n3668), .ZN(\DP/RegA1/N21 ) );
  AOI22_X1 U4729 ( .A1(\DP/RegALU2/N22 ), .A2(n2420), .B1(\DP/RegA_out[19] ), 
        .B2(n2422), .ZN(n3669) );
  OAI21_X1 U4730 ( .B1(n4448), .B2(n3693), .A(n3669), .ZN(\DP/RegA1/N22 ) );
  AOI22_X1 U4731 ( .A1(\DP/RegALU2/N23 ), .A2(n2420), .B1(\DP/RegA_out[20] ), 
        .B2(n3691), .ZN(n3670) );
  OAI21_X1 U4732 ( .B1(n4450), .B2(n2423), .A(n3670), .ZN(\DP/RegA1/N23 ) );
  AOI22_X1 U4733 ( .A1(\DP/RegALU2/N24 ), .A2(n2420), .B1(\DP/RegA_out[21] ), 
        .B2(n3691), .ZN(n3671) );
  OAI21_X1 U4734 ( .B1(n4554), .B2(n3693), .A(n3671), .ZN(\DP/RegA1/N24 ) );
  AOI22_X1 U4735 ( .A1(\DP/RegALU2/N25 ), .A2(n2420), .B1(\DP/RegA_out[22] ), 
        .B2(n2422), .ZN(n3672) );
  OAI21_X1 U4736 ( .B1(n4454), .B2(n2423), .A(n3672), .ZN(\DP/RegA1/N25 ) );
  INV_X1 U4737 ( .A(n4455), .ZN(n3674) );
  NOR2_X1 U4738 ( .A1(n2461), .A2(n2366), .ZN(\DP/RegALU2/N26 ) );
  AOI22_X1 U4739 ( .A1(\DP/RegALU2/N26 ), .A2(n2420), .B1(\DP/RegA_out[23] ), 
        .B2(n3691), .ZN(n3673) );
  OAI21_X1 U4740 ( .B1(n3674), .B2(n3693), .A(n3673), .ZN(\DP/RegA1/N26 ) );
  INV_X1 U4741 ( .A(n4457), .ZN(n3676) );
  NOR2_X1 U4742 ( .A1(n2460), .A2(n2393), .ZN(\DP/RegALU2/N27 ) );
  AOI22_X1 U4743 ( .A1(\DP/RegALU2/N27 ), .A2(n2420), .B1(\DP/RegA_out[24] ), 
        .B2(n2422), .ZN(n3675) );
  OAI21_X1 U4744 ( .B1(n3676), .B2(n2423), .A(n3675), .ZN(\DP/RegA1/N27 ) );
  AOI22_X1 U4745 ( .A1(\DP/RegALU2/N28 ), .A2(n2420), .B1(\DP/RegA_out[25] ), 
        .B2(n2422), .ZN(n3677) );
  OAI21_X1 U4746 ( .B1(n4557), .B2(n3693), .A(n3677), .ZN(\DP/RegA1/N28 ) );
  AOI22_X1 U4747 ( .A1(\DP/RegALU2/N29 ), .A2(n2420), .B1(\DP/RegA_out[26] ), 
        .B2(n3691), .ZN(n3678) );
  OAI21_X1 U4748 ( .B1(n4463), .B2(n2423), .A(n3678), .ZN(\DP/RegA1/N29 ) );
  AOI22_X1 U4749 ( .A1(\DP/RegA_out[0] ), .A2(n3691), .B1(n2421), .B2(
        \DP/RegALU2/N3 ), .ZN(n3679) );
  OAI21_X1 U4750 ( .B1(n4504), .B2(n3693), .A(n3679), .ZN(\DP/RegA1/N3 ) );
  AOI22_X1 U4751 ( .A1(\DP/RegALU2/N30 ), .A2(n2421), .B1(\DP/RegA_out[27] ), 
        .B2(n2422), .ZN(n3680) );
  OAI21_X1 U4752 ( .B1(n4550), .B2(n2423), .A(n3680), .ZN(\DP/RegA1/N30 ) );
  AOI22_X1 U4753 ( .A1(\DP/RegALU2/N31 ), .A2(n2420), .B1(\DP/RegA_out[28] ), 
        .B2(n3691), .ZN(n3681) );
  AOI22_X1 U4755 ( .A1(\DP/RegALU2/N32 ), .A2(n2421), .B1(\DP/RegA_out[29] ), 
        .B2(n2422), .ZN(n3682) );
  OAI21_X1 U4756 ( .B1(n4469), .B2(n3693), .A(n3682), .ZN(\DP/RegA1/N32 ) );
  AOI22_X1 U4757 ( .A1(\DP/RegALU2/N33 ), .A2(n2420), .B1(\DP/RegA_out[30] ), 
        .B2(n3691), .ZN(n3683) );
  AOI22_X1 U4759 ( .A1(\DP/RegA_out[31] ), .A2(n3691), .B1(\DP/RegALU2/N34 ), 
        .B2(n2420), .ZN(n3684) );
  OAI21_X1 U4760 ( .B1(n4549), .B2(n2423), .A(n3684), .ZN(\DP/RegA1/N34 ) );
  AOI22_X1 U4761 ( .A1(\DP/RegA_out[1] ), .A2(n3691), .B1(n2421), .B2(
        \DP/RegALU2/N4 ), .ZN(n3685) );
  OAI21_X1 U4762 ( .B1(n4502), .B2(n2423), .A(n3685), .ZN(\DP/RegA1/N4 ) );
  AOI22_X1 U4763 ( .A1(\DP/RegA_out[2] ), .A2(n3691), .B1(n2421), .B2(
        \DP/RegALU2/N5 ), .ZN(n3686) );
  OAI21_X1 U4764 ( .B1(n4494), .B2(n2423), .A(n3686), .ZN(\DP/RegA1/N5 ) );
  AOI22_X1 U4765 ( .A1(\DP/RegA_out[3] ), .A2(n3691), .B1(n2421), .B2(
        \DP/RegALU2/N6 ), .ZN(n3687) );
  OAI21_X1 U4766 ( .B1(n4492), .B2(n2423), .A(n3687), .ZN(\DP/RegA1/N6 ) );
  AOI22_X1 U4767 ( .A1(\DP/RegA_out[4] ), .A2(n3691), .B1(n2421), .B2(
        \DP/RegALU2/N7 ), .ZN(n3688) );
  OAI21_X1 U4768 ( .B1(n4561), .B2(n2423), .A(n3688), .ZN(\DP/RegA1/N7 ) );
  AOI22_X1 U4769 ( .A1(\DP/RegA_out[5] ), .A2(n3691), .B1(n2421), .B2(
        \DP/RegALU2/N8 ), .ZN(n3689) );
  OAI21_X1 U4770 ( .B1(n4517), .B2(n2423), .A(n3689), .ZN(\DP/RegA1/N8 ) );
  AOI22_X1 U4771 ( .A1(\DP/RegA_out[6] ), .A2(n3691), .B1(n2421), .B2(
        \DP/RegALU2/N9 ), .ZN(n3692) );
  OAI21_X1 U4772 ( .B1(n4520), .B2(n2423), .A(n3692), .ZN(\DP/RegA1/N9 ) );
  NAND2_X1 U4773 ( .A1(\DP/ALU0/s_A_LOGIC[7] ), .A2(\DP/ALU0/S_B_LOGIC[7] ), 
        .ZN(n3718) );
  XNOR2_X1 U4774 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[7] ), .ZN(n3720) );
  XNOR2_X1 U4775 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[5] ), .ZN(n4011) );
  XNOR2_X1 U4776 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[4] ), .ZN(n4031) );
  XNOR2_X1 U4777 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[3] ), .ZN(n4033) );
  XNOR2_X1 U4778 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[2] ), .ZN(n4035) );
  XNOR2_X1 U4779 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[1] ), .ZN(n4037) );
  INV_X1 U4780 ( .A(\DP/ALU0/S_B_ADDER[0] ), .ZN(n4014) );
  NOR2_X1 U4781 ( .A1(\DP/ALU0/s_A_ADDER[0] ), .A2(n4014), .ZN(n3694) );
  AOI21_X1 U4782 ( .B1(n2450), .B2(n4014), .A(n3694), .ZN(n4036) );
  XNOR2_X1 U4783 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[6] ), .ZN(n4012) );
  NOR2_X1 U4784 ( .A1(n3696), .A2(n3695), .ZN(n4101) );
  XOR2_X1 U4786 ( .A(\DP/ALU0/s_A_LOGIC[7] ), .B(\DP/ALU0/S_B_LOGIC[7] ), .Z(
        n3697) );
  AOI22_X1 U4787 ( .A1(n4009), .A2(n2430), .B1(n4231), .B2(n3697), .ZN(n3717)
         );
  XNOR2_X1 U4788 ( .A(n3819), .B(\DP/ALU0/S_B_SHIFT[0] ), .ZN(n4096) );
  XNOR2_X1 U4789 ( .A(n3819), .B(\DP/ALU0/S_B_SHIFT[2] ), .ZN(n4205) );
  INV_X1 U4790 ( .A(\DP/ALU0/s_A_SHIFT[6] ), .ZN(n4075) );
  INV_X1 U4791 ( .A(\DP/ALU0/S_B_SHIFT[3] ), .ZN(n3841) );
  INV_X1 U4792 ( .A(\DP/ALU0/S_B_SHIFT[4] ), .ZN(n3840) );
  NAND3_X1 U4793 ( .A1(n3841), .A2(n3840), .A3(n3819), .ZN(n4171) );
  AOI21_X1 U4794 ( .B1(\DP/ALU0/s_SHIFT[1] ), .B2(\DP/ALU0/s_SHIFT[0] ), .A(
        n3819), .ZN(n3698) );
  NOR2_X1 U4795 ( .A1(\DP/ALU0/S_B_SHIFT[3] ), .A2(n3840), .ZN(n3818) );
  NAND2_X1 U4796 ( .A1(n3698), .A2(n3818), .ZN(n4091) );
  INV_X1 U4797 ( .A(n4091), .ZN(n3713) );
  NAND3_X1 U4798 ( .A1(\DP/ALU0/S_B_SHIFT[3] ), .A2(n3698), .A3(n3840), .ZN(
        n4092) );
  NOR2_X1 U4799 ( .A1(\DP/ALU0/S_B_SHIFT[3] ), .A2(\DP/ALU0/S_B_SHIFT[4] ), 
        .ZN(n3842) );
  NAND2_X1 U4800 ( .A1(n3842), .A2(n3698), .ZN(n4090) );
  INV_X1 U4801 ( .A(\DP/ALU0/s_A_SHIFT[13] ), .ZN(n4088) );
  OAI22_X1 U4802 ( .A1(n25), .A2(n4092), .B1(n4090), .B2(n4088), .ZN(n3699) );
  AOI21_X1 U4803 ( .B1(n3713), .B2(\DP/ALU0/s_A_SHIFT[29] ), .A(n3699), .ZN(
        n3700) );
  OAI21_X1 U4804 ( .B1(n4075), .B2(n4171), .A(n3700), .ZN(n3747) );
  AOI22_X1 U4805 ( .A1(n4083), .A2(\DP/ALU0/s_A_SHIFT[9] ), .B1(n3713), .B2(
        \DP/ALU0/s_A_SHIFT[25] ), .ZN(n3702) );
  NAND2_X1 U4806 ( .A1(\DP/ALU0/s_A_SHIFT[2] ), .A2(n4152), .ZN(n3701) );
  OAI211_X1 U4807 ( .C1(n18), .C2(n4092), .A(n3702), .B(n3701), .ZN(n4197) );
  AOI22_X1 U4808 ( .A1(n2424), .A2(n3747), .B1(n4197), .B2(n4205), .ZN(n3725)
         );
  INV_X1 U4809 ( .A(n4092), .ZN(n4082) );
  INV_X1 U4810 ( .A(n45), .ZN(n3868) );
  AOI22_X1 U4811 ( .A1(n3713), .A2(\DP/ALU0/s_A_SHIFT[27] ), .B1(n4082), .B2(
        n3868), .ZN(n3704) );
  AOI22_X1 U4812 ( .A1(n4083), .A2(\DP/ALU0/s_A_SHIFT[11] ), .B1(
        \DP/ALU0/s_A_SHIFT[4] ), .B2(n4152), .ZN(n3703) );
  NAND2_X1 U4813 ( .A1(n3704), .A2(n3703), .ZN(n3724) );
  AOI22_X1 U4814 ( .A1(n4083), .A2(\DP/ALU0/s_A_SHIFT[7] ), .B1(n4082), .B2(
        \DP/ALU0/s_A_SHIFT[15] ), .ZN(n3706) );
  NAND2_X1 U4815 ( .A1(\DP/ALU0/s_A_SHIFT[0] ), .A2(n4152), .ZN(n3705) );
  OAI211_X1 U4816 ( .C1(n42), .C2(n4091), .A(n3706), .B(n3705), .ZN(n4086) );
  AOI22_X1 U4817 ( .A1(n2425), .A2(n3724), .B1(n4086), .B2(n2426), .ZN(n4216)
         );
  AOI22_X1 U4818 ( .A1(n2427), .A2(n3725), .B1(n4216), .B2(n2429), .ZN(n4233)
         );
  AOI22_X1 U4820 ( .A1(n4083), .A2(\DP/ALU0/s_A_SHIFT[14] ), .B1(n3713), .B2(
        \DP/ALU0/s_A_SHIFT[30] ), .ZN(n3708) );
  NAND2_X1 U4821 ( .A1(n4152), .A2(\DP/ALU0/s_A_SHIFT[7] ), .ZN(n3707) );
  OAI211_X1 U4822 ( .C1(n22), .C2(n4092), .A(n3708), .B(n3707), .ZN(n3758) );
  AOI22_X1 U4823 ( .A1(n4083), .A2(\DP/ALU0/s_A_SHIFT[10] ), .B1(
        \DP/ALU0/s_A_SHIFT[3] ), .B2(n4152), .ZN(n3710) );
  NAND2_X1 U4824 ( .A1(n3713), .A2(\DP/ALU0/s_A_SHIFT[26] ), .ZN(n3709) );
  OAI211_X1 U4825 ( .C1(n15), .C2(n4092), .A(n3710), .B(n3709), .ZN(n4207) );
  AOI22_X1 U4826 ( .A1(n2425), .A2(n3758), .B1(n4207), .B2(n2426), .ZN(n3737)
         );
  INV_X1 U4827 ( .A(\DP/ALU0/s_A_SHIFT[12] ), .ZN(n4125) );
  INV_X1 U4828 ( .A(\DP/ALU0/s_A_SHIFT[5] ), .ZN(n4087) );
  OAI22_X1 U4829 ( .A1(n4090), .A2(n4125), .B1(n4087), .B2(n4171), .ZN(n3711)
         );
  AOI21_X1 U4830 ( .B1(n3713), .B2(\DP/ALU0/s_A_SHIFT[28] ), .A(n3711), .ZN(
        n3712) );
  OAI21_X1 U4831 ( .B1(n20), .B2(n4092), .A(n3712), .ZN(n3736) );
  AOI22_X1 U4832 ( .A1(n4083), .A2(\DP/ALU0/s_A_SHIFT[8] ), .B1(n3713), .B2(
        \DP/ALU0/s_A_SHIFT[24] ), .ZN(n3715) );
  NAND2_X1 U4833 ( .A1(\DP/ALU0/s_A_SHIFT[1] ), .A2(n4152), .ZN(n3714) );
  OAI211_X1 U4834 ( .C1(n13), .C2(n4092), .A(n3715), .B(n3714), .ZN(n4188) );
  AOI22_X1 U4835 ( .A1(n2424), .A2(n3736), .B1(n4188), .B2(n2426), .ZN(n4225)
         );
  AOI22_X1 U4836 ( .A1(n2428), .A2(n3737), .B1(n4225), .B2(n4223), .ZN(n3726)
         );
  AOI22_X1 U4837 ( .A1(n2432), .A2(n4233), .B1(n4234), .B2(n3726), .ZN(n3716)
         );
  OAI211_X1 U4838 ( .C1(n4239), .C2(n3718), .A(n3717), .B(n3716), .ZN(
        \DP/RegALU1/N10 ) );
  NAND2_X1 U4839 ( .A1(\DP/ALU0/s_A_LOGIC[8] ), .A2(\DP/ALU0/S_B_LOGIC[8] ), 
        .ZN(n3729) );
  XNOR2_X1 U4840 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[8] ), .ZN(n3731) );
  FA_X1 U4841 ( .A(\DP/ALU0/s_A_ADDER[7] ), .B(n3720), .CI(n3719), .CO(n3730), 
        .S(n4009) );
  XOR2_X1 U4842 ( .A(\DP/ALU0/s_A_LOGIC[8] ), .B(\DP/ALU0/S_B_LOGIC[8] ), .Z(
        n3721) );
  AOI22_X1 U4843 ( .A1(n3998), .A2(n2431), .B1(n4231), .B2(n3721), .ZN(n3728)
         );
  INV_X1 U4844 ( .A(\DP/ALU0/s_A_SHIFT[31] ), .ZN(n4170) );
  NAND3_X1 U4845 ( .A1(n3840), .A2(\DP/ALU0/S_B_SHIFT[3] ), .A3(n3819), .ZN(
        n4150) );
  INV_X1 U4846 ( .A(n4150), .ZN(n4167) );
  AOI22_X1 U4847 ( .A1(\DP/ALU0/s_A_SHIFT[0] ), .A2(n4167), .B1(
        \DP/ALU0/s_A_SHIFT[8] ), .B2(n4152), .ZN(n3723) );
  INV_X1 U4848 ( .A(n42), .ZN(n4166) );
  AOI22_X1 U4849 ( .A1(n4083), .A2(\DP/ALU0/s_A_SHIFT[15] ), .B1(n4082), .B2(
        n4166), .ZN(n3722) );
  OAI211_X1 U4850 ( .C1(n4091), .C2(n4170), .A(n3723), .B(n3722), .ZN(n3769)
         );
  AOI22_X1 U4851 ( .A1(n2424), .A2(n3769), .B1(n3724), .B2(n2426), .ZN(n3748)
         );
  AOI22_X1 U4852 ( .A1(n2428), .A2(n3748), .B1(n3725), .B2(n4223), .ZN(n3738)
         );
  AOI22_X1 U4853 ( .A1(n2432), .A2(n3726), .B1(n4234), .B2(n3738), .ZN(n3727)
         );
  OAI211_X1 U4854 ( .C1(n2433), .C2(n3729), .A(n3728), .B(n3727), .ZN(
        \DP/RegALU1/N11 ) );
  NAND2_X1 U4855 ( .A1(\DP/ALU0/s_A_LOGIC[9] ), .A2(\DP/ALU0/S_B_LOGIC[9] ), 
        .ZN(n3741) );
  XNOR2_X1 U4856 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[9] ), .ZN(n3743) );
  FA_X1 U4857 ( .A(\DP/ALU0/s_A_ADDER[8] ), .B(n3731), .CI(n3730), .CO(n3742), 
        .S(n3998) );
  XOR2_X1 U4858 ( .A(\DP/ALU0/s_A_LOGIC[9] ), .B(\DP/ALU0/S_B_LOGIC[9] ), .Z(
        n3732) );
  AOI22_X1 U4859 ( .A1(n3999), .A2(n2431), .B1(n4231), .B2(n3732), .ZN(n3740)
         );
  INV_X1 U4860 ( .A(\DP/ALU0/s_SHIFT[1] ), .ZN(n3733) );
  NOR3_X1 U4861 ( .A1(\DP/ALU0/s_SHIFT[0] ), .A2(n3733), .A3(n4170), .ZN(n3839) );
  NAND2_X1 U4862 ( .A1(n3818), .A2(n3839), .ZN(n3820) );
  INV_X1 U4863 ( .A(n3820), .ZN(n3801) );
  AOI21_X1 U4864 ( .B1(n4152), .B2(\DP/ALU0/s_A_SHIFT[9] ), .A(n3801), .ZN(
        n3735) );
  AOI22_X1 U4865 ( .A1(n4082), .A2(\DP/ALU0/s_A_SHIFT[24] ), .B1(
        \DP/ALU0/s_A_SHIFT[1] ), .B2(n4167), .ZN(n3734) );
  OAI211_X1 U4866 ( .C1(n13), .C2(n4090), .A(n3735), .B(n3734), .ZN(n3780) );
  AOI22_X1 U4867 ( .A1(n2425), .A2(n3780), .B1(n3736), .B2(n2426), .ZN(n3759)
         );
  AOI22_X1 U4868 ( .A1(n2428), .A2(n3759), .B1(n3737), .B2(n4223), .ZN(n3749)
         );
  AOI22_X1 U4869 ( .A1(n2432), .A2(n3738), .B1(n4234), .B2(n3749), .ZN(n3739)
         );
  OAI211_X1 U4870 ( .C1(n2433), .C2(n3741), .A(n3740), .B(n3739), .ZN(
        \DP/RegALU1/N12 ) );
  NAND2_X1 U4871 ( .A1(\DP/ALU0/s_A_LOGIC[10] ), .A2(\DP/ALU0/S_B_LOGIC[10] ), 
        .ZN(n3752) );
  XNOR2_X1 U4872 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[10] ), .ZN(n3754) );
  FA_X1 U4873 ( .A(\DP/ALU0/s_A_ADDER[9] ), .B(n3743), .CI(n3742), .CO(n3753), 
        .S(n3999) );
  XOR2_X1 U4874 ( .A(\DP/ALU0/s_A_LOGIC[10] ), .B(\DP/ALU0/S_B_LOGIC[10] ), 
        .Z(n3744) );
  AOI22_X1 U4875 ( .A1(n4000), .A2(n2431), .B1(n4231), .B2(n3744), .ZN(n3751)
         );
  AOI21_X1 U4876 ( .B1(\DP/ALU0/s_A_SHIFT[2] ), .B2(n4167), .A(n3801), .ZN(
        n3746) );
  AOI22_X1 U4877 ( .A1(n4082), .A2(\DP/ALU0/s_A_SHIFT[25] ), .B1(
        \DP/ALU0/s_A_SHIFT[10] ), .B2(n4152), .ZN(n3745) );
  OAI211_X1 U4878 ( .C1(n18), .C2(n4090), .A(n3746), .B(n3745), .ZN(n3791) );
  AOI22_X1 U4879 ( .A1(n2424), .A2(n3791), .B1(n3747), .B2(n2426), .ZN(n3770)
         );
  AOI22_X1 U4880 ( .A1(n2428), .A2(n3770), .B1(n3748), .B2(n2429), .ZN(n3760)
         );
  AOI22_X1 U4881 ( .A1(n2432), .A2(n3749), .B1(n4234), .B2(n3760), .ZN(n3750)
         );
  OAI211_X1 U4882 ( .C1(n2433), .C2(n3752), .A(n3751), .B(n3750), .ZN(
        \DP/RegALU1/N13 ) );
  NAND2_X1 U4883 ( .A1(\DP/ALU0/s_A_LOGIC[11] ), .A2(\DP/ALU0/S_B_LOGIC[11] ), 
        .ZN(n3763) );
  XNOR2_X1 U4884 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[11] ), .ZN(n3765) );
  FA_X1 U4885 ( .A(\DP/ALU0/s_A_ADDER[10] ), .B(n3754), .CI(n3753), .CO(n3764), 
        .S(n4000) );
  XOR2_X1 U4886 ( .A(\DP/ALU0/s_A_LOGIC[11] ), .B(\DP/ALU0/S_B_LOGIC[11] ), 
        .Z(n3755) );
  AOI22_X1 U4887 ( .A1(n4001), .A2(n2431), .B1(n4231), .B2(n3755), .ZN(n3762)
         );
  AOI21_X1 U4888 ( .B1(n4152), .B2(\DP/ALU0/s_A_SHIFT[11] ), .A(n3801), .ZN(
        n3757) );
  AOI22_X1 U4889 ( .A1(n4082), .A2(\DP/ALU0/s_A_SHIFT[26] ), .B1(
        \DP/ALU0/s_A_SHIFT[3] ), .B2(n4167), .ZN(n3756) );
  OAI211_X1 U4890 ( .C1(n15), .C2(n4090), .A(n3757), .B(n3756), .ZN(n3804) );
  AOI22_X1 U4891 ( .A1(n2425), .A2(n3804), .B1(n3758), .B2(n2426), .ZN(n3781)
         );
  AOI22_X1 U4892 ( .A1(n2428), .A2(n3781), .B1(n3759), .B2(n2429), .ZN(n3771)
         );
  AOI22_X1 U4893 ( .A1(n2432), .A2(n3760), .B1(n4234), .B2(n3771), .ZN(n3761)
         );
  OAI211_X1 U4894 ( .C1(n2433), .C2(n3763), .A(n3762), .B(n3761), .ZN(
        \DP/RegALU1/N14 ) );
  NAND2_X1 U4895 ( .A1(\DP/ALU0/s_A_LOGIC[12] ), .A2(\DP/ALU0/S_B_LOGIC[12] ), 
        .ZN(n3774) );
  XNOR2_X1 U4896 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[12] ), .ZN(n3776) );
  FA_X1 U4897 ( .A(\DP/ALU0/s_A_ADDER[11] ), .B(n3765), .CI(n3764), .CO(n3775), 
        .S(n4001) );
  XOR2_X1 U4898 ( .A(\DP/ALU0/s_A_LOGIC[12] ), .B(\DP/ALU0/S_B_LOGIC[12] ), 
        .Z(n3766) );
  AOI22_X1 U4899 ( .A1(n4002), .A2(n2431), .B1(n4231), .B2(n3766), .ZN(n3773)
         );
  AOI21_X1 U4900 ( .B1(\DP/ALU0/s_A_SHIFT[4] ), .B2(n4167), .A(n3801), .ZN(
        n3768) );
  AOI22_X1 U4901 ( .A1(n4082), .A2(\DP/ALU0/s_A_SHIFT[27] ), .B1(
        \DP/ALU0/s_A_SHIFT[12] ), .B2(n4152), .ZN(n3767) );
  OAI211_X1 U4902 ( .C1(n45), .C2(n4090), .A(n3768), .B(n3767), .ZN(n3824) );
  AOI22_X1 U4903 ( .A1(n2425), .A2(n3824), .B1(n3769), .B2(n2426), .ZN(n3793)
         );
  AOI22_X1 U4904 ( .A1(n2428), .A2(n3793), .B1(n3770), .B2(n2429), .ZN(n3782)
         );
  AOI22_X1 U4905 ( .A1(n2432), .A2(n3771), .B1(n4234), .B2(n3782), .ZN(n3772)
         );
  OAI211_X1 U4906 ( .C1(n2433), .C2(n3774), .A(n3773), .B(n3772), .ZN(
        \DP/RegALU1/N15 ) );
  NAND2_X1 U4907 ( .A1(\DP/ALU0/s_A_LOGIC[13] ), .A2(\DP/ALU0/S_B_LOGIC[13] ), 
        .ZN(n3785) );
  XNOR2_X1 U4908 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[13] ), .ZN(n3787) );
  FA_X1 U4909 ( .A(\DP/ALU0/s_A_ADDER[12] ), .B(n3776), .CI(n3775), .CO(n3786), 
        .S(n4002) );
  XOR2_X1 U4910 ( .A(\DP/ALU0/s_A_LOGIC[13] ), .B(\DP/ALU0/S_B_LOGIC[13] ), 
        .Z(n3777) );
  AOI22_X1 U4911 ( .A1(n4003), .A2(n2431), .B1(n4231), .B2(n3777), .ZN(n3784)
         );
  AOI21_X1 U4912 ( .B1(n4152), .B2(\DP/ALU0/s_A_SHIFT[13] ), .A(n3801), .ZN(
        n3779) );
  AOI22_X1 U4913 ( .A1(n4082), .A2(\DP/ALU0/s_A_SHIFT[28] ), .B1(
        \DP/ALU0/s_A_SHIFT[5] ), .B2(n4167), .ZN(n3778) );
  OAI211_X1 U4914 ( .C1(n20), .C2(n4090), .A(n3779), .B(n3778), .ZN(n3845) );
  AOI22_X1 U4915 ( .A1(n2425), .A2(n3845), .B1(n3780), .B2(n4205), .ZN(n3805)
         );
  AOI22_X1 U4916 ( .A1(n2428), .A2(n3805), .B1(n3781), .B2(n2429), .ZN(n3794)
         );
  AOI22_X1 U4917 ( .A1(n2432), .A2(n3782), .B1(n4234), .B2(n3794), .ZN(n3783)
         );
  OAI211_X1 U4918 ( .C1(n2433), .C2(n3785), .A(n3784), .B(n3783), .ZN(
        \DP/RegALU1/N16 ) );
  NAND2_X1 U4919 ( .A1(\DP/ALU0/s_A_LOGIC[14] ), .A2(\DP/ALU0/S_B_LOGIC[14] ), 
        .ZN(n3797) );
  XNOR2_X1 U4920 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[14] ), .ZN(n3799) );
  FA_X1 U4921 ( .A(\DP/ALU0/s_A_ADDER[13] ), .B(n3787), .CI(n3786), .CO(n3798), 
        .S(n4003) );
  XOR2_X1 U4922 ( .A(\DP/ALU0/s_A_LOGIC[14] ), .B(\DP/ALU0/S_B_LOGIC[14] ), 
        .Z(n3788) );
  AOI22_X1 U4923 ( .A1(n4004), .A2(n2431), .B1(n4231), .B2(n3788), .ZN(n3796)
         );
  INV_X1 U4924 ( .A(\DP/ALU0/s_A_SHIFT[14] ), .ZN(n4149) );
  OAI21_X1 U4925 ( .B1(n4171), .B2(n4149), .A(n3820), .ZN(n3790) );
  OAI22_X1 U4926 ( .A1(n25), .A2(n4090), .B1(n4075), .B2(n4150), .ZN(n3789) );
  AOI211_X1 U4927 ( .C1(n4082), .C2(\DP/ALU0/s_A_SHIFT[29] ), .A(n3790), .B(
        n3789), .ZN(n3852) );
  INV_X1 U4928 ( .A(n3852), .ZN(n3792) );
  AOI22_X1 U4929 ( .A1(n2425), .A2(n3792), .B1(n3791), .B2(n2426), .ZN(n3826)
         );
  AOI22_X1 U4930 ( .A1(n2428), .A2(n3826), .B1(n3793), .B2(n2429), .ZN(n3806)
         );
  AOI22_X1 U4931 ( .A1(n2432), .A2(n3794), .B1(n4234), .B2(n3806), .ZN(n3795)
         );
  OAI211_X1 U4932 ( .C1(n4239), .C2(n3797), .A(n3796), .B(n3795), .ZN(
        \DP/RegALU1/N17 ) );
  NAND2_X1 U4933 ( .A1(\DP/ALU0/s_A_LOGIC[15] ), .A2(\DP/ALU0/S_B_LOGIC[15] ), 
        .ZN(n3809) );
  XNOR2_X1 U4934 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[15] ), .ZN(n3813) );
  FA_X1 U4935 ( .A(\DP/ALU0/s_A_ADDER[14] ), .B(n3799), .CI(n3798), .CO(n3812), 
        .S(n4004) );
  XOR2_X1 U4936 ( .A(\DP/ALU0/s_A_LOGIC[15] ), .B(\DP/ALU0/S_B_LOGIC[15] ), 
        .Z(n3800) );
  AOI22_X1 U4937 ( .A1(n4005), .A2(n2431), .B1(n4231), .B2(n3800), .ZN(n3808)
         );
  AOI21_X1 U4938 ( .B1(\DP/ALU0/s_A_SHIFT[15] ), .B2(n4152), .A(n3801), .ZN(
        n3803) );
  AOI22_X1 U4939 ( .A1(n4082), .A2(\DP/ALU0/s_A_SHIFT[30] ), .B1(
        \DP/ALU0/s_A_SHIFT[7] ), .B2(n4167), .ZN(n3802) );
  OAI211_X1 U4940 ( .C1(n22), .C2(n4090), .A(n3803), .B(n3802), .ZN(n3871) );
  AOI22_X1 U4941 ( .A1(n2425), .A2(n3871), .B1(n3804), .B2(n4205), .ZN(n3846)
         );
  AOI22_X1 U4942 ( .A1(n2428), .A2(n3846), .B1(n3805), .B2(n2429), .ZN(n3828)
         );
  AOI22_X1 U4943 ( .A1(n2432), .A2(n3806), .B1(n4234), .B2(n3828), .ZN(n3807)
         );
  OAI211_X1 U4944 ( .C1(n4239), .C2(n3809), .A(n3808), .B(n3807), .ZN(
        \DP/RegALU1/N18 ) );
  FA_X1 U4945 ( .A(\DP/ALU0/s_A_ADDER[15] ), .B(n3813), .CI(n3812), .CO(n3858), 
        .S(n4005) );
  XNOR2_X1 U4946 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[16] ), .ZN(n3814) );
  NAND2_X1 U4947 ( .A1(\DP/ALU0/s_A_ADDER[16] ), .A2(n3814), .ZN(n3854) );
  INV_X1 U4948 ( .A(n3854), .ZN(n3815) );
  NOR2_X1 U4949 ( .A1(\DP/ALU0/s_A_ADDER[16] ), .A2(n3814), .ZN(n3857) );
  NOR2_X1 U4950 ( .A1(n3815), .A2(n3857), .ZN(n3834) );
  XOR2_X1 U4951 ( .A(n3858), .B(n3834), .Z(n4049) );
  AOI22_X1 U4952 ( .A1(n4049), .A2(n2431), .B1(n4164), .B2(
        \DP/ALU0/S_B_LHI[0] ), .ZN(n3831) );
  NOR2_X1 U4953 ( .A1(n14), .A2(n9), .ZN(n3817) );
  AOI22_X1 U4954 ( .A1(n14), .A2(n9), .B1(n3817), .B2(n4239), .ZN(n3816) );
  OAI21_X1 U4955 ( .B1(n3817), .B2(n4231), .A(n3816), .ZN(n3830) );
  NOR2_X1 U4956 ( .A1(n42), .A2(n4090), .ZN(n3823) );
  NAND2_X1 U4957 ( .A1(n3819), .A2(n3818), .ZN(n4148) );
  INV_X1 U4958 ( .A(n4148), .ZN(n4168) );
  AOI22_X1 U4959 ( .A1(\DP/ALU0/s_A_SHIFT[0] ), .A2(n4168), .B1(
        \DP/ALU0/s_A_SHIFT[8] ), .B2(n4167), .ZN(n3821) );
  OAI211_X1 U4960 ( .C1(n13), .C2(n4171), .A(n3821), .B(n3820), .ZN(n3822) );
  AOI211_X1 U4961 ( .C1(\DP/ALU0/s_A_SHIFT[31] ), .C2(n4082), .A(n3823), .B(
        n3822), .ZN(n3881) );
  INV_X1 U4962 ( .A(n3824), .ZN(n3825) );
  OAI22_X1 U4963 ( .A1(n2426), .A2(n3881), .B1(n3825), .B2(n2425), .ZN(n3853)
         );
  INV_X1 U4964 ( .A(n3853), .ZN(n3827) );
  AOI22_X1 U4965 ( .A1(n2428), .A2(n3827), .B1(n3826), .B2(n2429), .ZN(n3847)
         );
  AOI22_X1 U4966 ( .A1(n2432), .A2(n3828), .B1(n4234), .B2(n3847), .ZN(n3829)
         );
  NAND3_X1 U4967 ( .A1(n3831), .A2(n3830), .A3(n3829), .ZN(\DP/RegALU1/N19 )
         );
  OR2_X1 U4968 ( .A1(w_EX_EN), .A2(n2461), .ZN(\DP/RegALU1/N2 ) );
  XNOR2_X1 U4969 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[17] ), .ZN(n3832) );
  NAND2_X1 U4970 ( .A1(\DP/ALU0/s_A_ADDER[17] ), .A2(n3832), .ZN(n3856) );
  NOR2_X1 U4971 ( .A1(\DP/ALU0/s_A_ADDER[17] ), .A2(n3832), .ZN(n3855) );
  INV_X1 U4972 ( .A(n3855), .ZN(n3833) );
  NAND2_X1 U4973 ( .A1(n3856), .A2(n3833), .ZN(n3890) );
  NAND2_X1 U4974 ( .A1(n3858), .A2(n3834), .ZN(n3891) );
  NAND2_X1 U4975 ( .A1(n3854), .A2(n3891), .ZN(n3835) );
  XOR2_X1 U4976 ( .A(n3890), .B(n3835), .Z(n4054) );
  NOR2_X1 U4977 ( .A1(n19), .A2(n17), .ZN(n3836) );
  AOI211_X1 U4978 ( .C1(n19), .C2(n17), .A(n3836), .B(n4178), .ZN(n3838) );
  NOR3_X1 U4979 ( .A1(n19), .A2(n17), .A3(n2433), .ZN(n3837) );
  AOI211_X1 U4980 ( .C1(\DP/ALU0/S_B_LHI[1] ), .C2(n4164), .A(n3838), .B(n3837), .ZN(n3849) );
  INV_X1 U4981 ( .A(\DP/ALU0/s_A_SHIFT[9] ), .ZN(n4093) );
  OAI21_X1 U4982 ( .B1(n3841), .B2(n3840), .A(n3839), .ZN(n4124) );
  NOR2_X1 U4983 ( .A1(n3842), .A2(n4124), .ZN(n3916) );
  INV_X1 U4984 ( .A(\DP/ALU0/s_A_SHIFT[1] ), .ZN(n4089) );
  OAI22_X1 U4985 ( .A1(n18), .A2(n4171), .B1(n4089), .B2(n4148), .ZN(n3843) );
  AOI211_X1 U4986 ( .C1(n4083), .C2(\DP/ALU0/s_A_SHIFT[24] ), .A(n3916), .B(
        n3843), .ZN(n3844) );
  OAI21_X1 U4987 ( .B1(n4093), .B2(n4150), .A(n3844), .ZN(n3909) );
  AOI22_X1 U4988 ( .A1(n2425), .A2(n3909), .B1(n3845), .B2(n4205), .ZN(n3872)
         );
  AOI22_X1 U4989 ( .A1(n2428), .A2(n3872), .B1(n3846), .B2(n2429), .ZN(n3863)
         );
  AOI22_X1 U4990 ( .A1(n2432), .A2(n3847), .B1(n4234), .B2(n3863), .ZN(n3848)
         );
  OAI211_X1 U4991 ( .C1(n4054), .C2(n2389), .A(n3849), .B(n3848), .ZN(
        \DP/RegALU1/N20 ) );
  AOI22_X1 U4992 ( .A1(\DP/ALU0/s_A_SHIFT[2] ), .A2(n4168), .B1(
        \DP/ALU0/s_A_SHIFT[10] ), .B2(n4167), .ZN(n3850) );
  OAI21_X1 U4993 ( .B1(n15), .B2(n4171), .A(n3850), .ZN(n3851) );
  AOI211_X1 U4994 ( .C1(n4083), .C2(\DP/ALU0/s_A_SHIFT[25] ), .A(n3916), .B(
        n3851), .ZN(n3917) );
  AOI22_X1 U4995 ( .A1(n2425), .A2(n3917), .B1(n3852), .B2(n2426), .ZN(n3882)
         );
  AOI22_X1 U4996 ( .A1(n2428), .A2(n3882), .B1(n3853), .B2(n2429), .ZN(n3878)
         );
  XNOR2_X1 U4997 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[18] ), .ZN(n3887) );
  OAI21_X1 U4998 ( .B1(n3855), .B2(n3854), .A(n3856), .ZN(n3889) );
  AOI21_X1 U4999 ( .B1(n3857), .B2(n3856), .A(n3855), .ZN(n3859) );
  MUX2_X1 U5000 ( .A(n3889), .B(n3859), .S(n3858), .Z(n3866) );
  AOI22_X1 U5001 ( .A1(n4008), .A2(n2431), .B1(n4164), .B2(
        \DP/ALU0/S_B_LHI[2] ), .ZN(n3865) );
  NOR2_X1 U5002 ( .A1(n16), .A2(n8), .ZN(n3860) );
  AOI211_X1 U5003 ( .C1(n16), .C2(n8), .A(n3860), .B(n4178), .ZN(n3862) );
  NOR3_X1 U5004 ( .A1(n16), .A2(n8), .A3(n4239), .ZN(n3861) );
  AOI211_X1 U5005 ( .C1(n3863), .C2(n2432), .A(n3862), .B(n3861), .ZN(n3864)
         );
  OAI211_X1 U5006 ( .C1(n4175), .C2(n3878), .A(n3865), .B(n3864), .ZN(
        \DP/RegALU1/N21 ) );
  FA_X1 U5007 ( .A(\DP/ALU0/s_A_ADDER[18] ), .B(n3887), .CI(n3866), .CO(n3867), 
        .S(n4008) );
  XNOR2_X1 U5008 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[19] ), .ZN(n3888) );
  XOR2_X1 U5009 ( .A(n3888), .B(\DP/ALU0/s_A_ADDER[19] ), .Z(n3886) );
  XOR2_X1 U5010 ( .A(n3867), .B(n3886), .Z(n4050) );
  AOI22_X1 U5011 ( .A1(n4050), .A2(n2431), .B1(n4164), .B2(
        \DP/ALU0/S_B_LHI[3] ), .ZN(n3877) );
  AOI22_X1 U5012 ( .A1(\DP/ALU0/s_A_SHIFT[11] ), .A2(n4167), .B1(n4152), .B2(
        n3868), .ZN(n3870) );
  AOI22_X1 U5013 ( .A1(n4083), .A2(\DP/ALU0/s_A_SHIFT[26] ), .B1(
        \DP/ALU0/s_A_SHIFT[3] ), .B2(n4168), .ZN(n3869) );
  INV_X1 U5014 ( .A(n3916), .ZN(n3948) );
  NAND3_X1 U5015 ( .A1(n3870), .A2(n3869), .A3(n3948), .ZN(n3936) );
  AOI22_X1 U5016 ( .A1(n2425), .A2(n3936), .B1(n3871), .B2(n4205), .ZN(n3910)
         );
  AOI22_X1 U5017 ( .A1(n2427), .A2(n3910), .B1(n3872), .B2(n2429), .ZN(n3896)
         );
  NOR2_X1 U5018 ( .A1(n46), .A2(n44), .ZN(n3873) );
  AOI211_X1 U5019 ( .C1(n46), .C2(n44), .A(n3873), .B(n4178), .ZN(n3875) );
  NOR3_X1 U5020 ( .A1(n46), .A2(n44), .A3(n2433), .ZN(n3874) );
  AOI211_X1 U5021 ( .C1(n3896), .C2(n4234), .A(n3875), .B(n3874), .ZN(n3876)
         );
  OAI211_X1 U5022 ( .C1(n2396), .C2(n3878), .A(n3877), .B(n3876), .ZN(
        \DP/RegALU1/N22 ) );
  INV_X1 U5023 ( .A(\DP/ALU0/s_A_SHIFT[4] ), .ZN(n4078) );
  OAI22_X1 U5024 ( .A1(n20), .A2(n4171), .B1(n4078), .B2(n4148), .ZN(n3880) );
  OAI21_X1 U5025 ( .B1(n4150), .B2(n4125), .A(n3948), .ZN(n3879) );
  AOI211_X1 U5026 ( .C1(n4083), .C2(\DP/ALU0/s_A_SHIFT[27] ), .A(n3880), .B(
        n3879), .ZN(n3951) );
  AOI22_X1 U5027 ( .A1(n2425), .A2(n3951), .B1(n3881), .B2(n2426), .ZN(n3918)
         );
  AOI22_X1 U5028 ( .A1(n2428), .A2(n3918), .B1(n3882), .B2(n2429), .ZN(n3913)
         );
  NOR2_X1 U5029 ( .A1(n21), .A2(n7), .ZN(n3883) );
  AOI211_X1 U5030 ( .C1(n21), .C2(n7), .A(n3883), .B(n4178), .ZN(n3885) );
  NOR3_X1 U5031 ( .A1(n21), .A2(n7), .A3(n2433), .ZN(n3884) );
  AOI211_X1 U5032 ( .C1(\DP/ALU0/S_B_LHI[4] ), .C2(n4164), .A(n3885), .B(n3884), .ZN(n3898) );
  AND2_X1 U5033 ( .A1(\DP/ALU0/s_A_ADDER[18] ), .A2(n3887), .ZN(n3893) );
  OAI21_X1 U5034 ( .B1(\DP/ALU0/s_A_ADDER[18] ), .B2(n3887), .A(n3886), .ZN(
        n3892) );
  NOR4_X1 U5035 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3905)
         );
  INV_X1 U5036 ( .A(n3905), .ZN(n3954) );
  XNOR2_X1 U5037 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[20] ), .ZN(n3894) );
  NAND2_X1 U5038 ( .A1(\DP/ALU0/s_A_ADDER[20] ), .A2(n3894), .ZN(n3903) );
  NOR2_X1 U5039 ( .A1(\DP/ALU0/s_A_ADDER[20] ), .A2(n3894), .ZN(n3922) );
  INV_X1 U5040 ( .A(n3922), .ZN(n3895) );
  NAND2_X1 U5041 ( .A1(n3903), .A2(n3895), .ZN(n3953) );
  AOI22_X1 U5042 ( .A1(n3896), .A2(n2432), .B1(n2431), .B2(n3997), .ZN(n3897)
         );
  OAI211_X1 U5043 ( .C1(n4175), .C2(n3913), .A(n3898), .B(n3897), .ZN(
        \DP/RegALU1/N23 ) );
  NOR2_X1 U5044 ( .A1(n26), .A2(n24), .ZN(n3899) );
  AOI211_X1 U5045 ( .C1(n26), .C2(n24), .A(n3899), .B(n4178), .ZN(n3901) );
  NOR3_X1 U5046 ( .A1(n26), .A2(n24), .A3(n4239), .ZN(n3900) );
  AOI211_X1 U5047 ( .C1(\DP/ALU0/S_B_LHI[5] ), .C2(n4164), .A(n3901), .B(n3900), .ZN(n3912) );
  XNOR2_X1 U5048 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[21] ), .ZN(n3902) );
  NAND2_X1 U5049 ( .A1(\DP/ALU0/s_A_ADDER[21] ), .A2(n3902), .ZN(n3924) );
  INV_X1 U5050 ( .A(n3924), .ZN(n3962) );
  NOR2_X1 U5051 ( .A1(\DP/ALU0/s_A_ADDER[21] ), .A2(n3902), .ZN(n3923) );
  NOR2_X1 U5052 ( .A1(n3962), .A2(n3923), .ZN(n3958) );
  NAND2_X1 U5053 ( .A1(n3904), .A2(n3903), .ZN(n3960) );
  NOR2_X1 U5054 ( .A1(n3905), .A2(n3960), .ZN(n3926) );
  NOR2_X1 U5055 ( .A1(n3926), .A2(n3922), .ZN(n3906) );
  XOR2_X1 U5056 ( .A(n3958), .B(n3906), .Z(n4058) );
  OAI22_X1 U5057 ( .A1(n25), .A2(n4171), .B1(n4087), .B2(n4148), .ZN(n3907) );
  AOI211_X1 U5058 ( .C1(n4083), .C2(\DP/ALU0/s_A_SHIFT[28] ), .A(n3916), .B(
        n3907), .ZN(n3908) );
  OAI21_X1 U5059 ( .B1(n4088), .B2(n4150), .A(n3908), .ZN(n3976) );
  AOI22_X1 U5060 ( .A1(n2425), .A2(n3976), .B1(n3909), .B2(n2426), .ZN(n3937)
         );
  AOI22_X1 U5061 ( .A1(n2427), .A2(n3937), .B1(n3910), .B2(n2429), .ZN(n3928)
         );
  AOI22_X1 U5062 ( .A1(n4058), .A2(n2431), .B1(n4234), .B2(n3928), .ZN(n3911)
         );
  OAI211_X1 U5063 ( .C1(n2396), .C2(n3913), .A(n3912), .B(n3911), .ZN(
        \DP/RegALU1/N24 ) );
  AOI22_X1 U5064 ( .A1(\DP/ALU0/s_A_SHIFT[6] ), .A2(n4168), .B1(
        \DP/ALU0/s_A_SHIFT[14] ), .B2(n4167), .ZN(n3914) );
  OAI21_X1 U5065 ( .B1(n22), .B2(n4171), .A(n3914), .ZN(n3915) );
  AOI211_X1 U5066 ( .C1(n4083), .C2(\DP/ALU0/s_A_SHIFT[29] ), .A(n3916), .B(
        n3915), .ZN(n3987) );
  AOI22_X1 U5067 ( .A1(n2425), .A2(n3987), .B1(n3917), .B2(n2426), .ZN(n3952)
         );
  AOI22_X1 U5068 ( .A1(n2427), .A2(n3952), .B1(n3918), .B2(n2429), .ZN(n3947)
         );
  NOR2_X1 U5069 ( .A1(n23), .A2(n6), .ZN(n3919) );
  AOI211_X1 U5070 ( .C1(n23), .C2(n6), .A(n3919), .B(n4178), .ZN(n3921) );
  NOR3_X1 U5071 ( .A1(n23), .A2(n6), .A3(n2433), .ZN(n3920) );
  AOI211_X1 U5072 ( .C1(\DP/ALU0/S_B_LHI[6] ), .C2(n4164), .A(n3921), .B(n3920), .ZN(n3930) );
  NOR2_X1 U5073 ( .A1(n3923), .A2(n3922), .ZN(n3961) );
  INV_X1 U5074 ( .A(n3961), .ZN(n3925) );
  OAI21_X1 U5075 ( .B1(n3926), .B2(n3925), .A(n3924), .ZN(n3938) );
  XNOR2_X1 U5076 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[22] ), .ZN(n3927) );
  NAND2_X1 U5077 ( .A1(\DP/ALU0/s_A_ADDER[22] ), .A2(n3927), .ZN(n3940) );
  INV_X1 U5078 ( .A(n3940), .ZN(n3956) );
  NOR2_X1 U5079 ( .A1(\DP/ALU0/s_A_ADDER[22] ), .A2(n3927), .ZN(n3955) );
  NOR2_X1 U5080 ( .A1(n3956), .A2(n3955), .ZN(n3959) );
  XOR2_X1 U5081 ( .A(n3938), .B(n3959), .Z(n4051) );
  AOI22_X1 U5082 ( .A1(n4051), .A2(n2430), .B1(n2432), .B2(n3928), .ZN(n3929)
         );
  OAI211_X1 U5083 ( .C1(n3947), .C2(n4175), .A(n3930), .B(n3929), .ZN(
        \DP/RegALU1/N25 ) );
  NOR2_X1 U5084 ( .A1(n43), .A2(n41), .ZN(n3931) );
  AOI211_X1 U5085 ( .C1(n43), .C2(n41), .A(n3931), .B(n4178), .ZN(n3933) );
  NOR3_X1 U5086 ( .A1(n43), .A2(n41), .A3(n4239), .ZN(n3932) );
  AOI211_X1 U5087 ( .C1(\DP/ALU0/S_B_LHI[7] ), .C2(n4164), .A(n3933), .B(n3932), .ZN(n3946) );
  AOI22_X1 U5088 ( .A1(n4152), .A2(n4166), .B1(\DP/ALU0/s_A_SHIFT[7] ), .B2(
        n4168), .ZN(n3935) );
  AOI22_X1 U5089 ( .A1(n4083), .A2(\DP/ALU0/s_A_SHIFT[30] ), .B1(
        \DP/ALU0/s_A_SHIFT[15] ), .B2(n4167), .ZN(n3934) );
  NAND3_X1 U5090 ( .A1(n3935), .A2(n3934), .A3(n3948), .ZN(n4116) );
  AOI22_X1 U5091 ( .A1(n2424), .A2(n4116), .B1(n3936), .B2(n2426), .ZN(n3977)
         );
  AOI22_X1 U5092 ( .A1(n2428), .A2(n3977), .B1(n3937), .B2(n2429), .ZN(n3970)
         );
  NAND2_X1 U5093 ( .A1(n3959), .A2(n3938), .ZN(n3939) );
  NAND2_X1 U5094 ( .A1(n3940), .A2(n3939), .ZN(n3944) );
  XNOR2_X1 U5095 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[23] ), .ZN(n3941) );
  NAND2_X1 U5096 ( .A1(\DP/ALU0/s_A_ADDER[23] ), .A2(n3941), .ZN(n3963) );
  NOR2_X1 U5097 ( .A1(\DP/ALU0/s_A_ADDER[23] ), .A2(n3941), .ZN(n3966) );
  INV_X1 U5098 ( .A(n3966), .ZN(n3942) );
  NAND2_X1 U5099 ( .A1(n3963), .A2(n3942), .ZN(n3943) );
  XNOR2_X1 U5100 ( .A(n3944), .B(n3943), .ZN(n4057) );
  AOI22_X1 U5101 ( .A1(n3970), .A2(n4234), .B1(n2431), .B2(n4057), .ZN(n3945)
         );
  OAI211_X1 U5102 ( .C1(n2396), .C2(n3947), .A(n3946), .B(n3945), .ZN(
        \DP/RegALU1/N26 ) );
  AOI22_X1 U5103 ( .A1(\DP/ALU0/s_A_SHIFT[8] ), .A2(n4168), .B1(n4152), .B2(
        \DP/ALU0/s_A_SHIFT[24] ), .ZN(n3949) );
  OAI211_X1 U5104 ( .C1(n13), .C2(n4150), .A(n3949), .B(n3948), .ZN(n3950) );
  AOI21_X1 U5105 ( .B1(n4083), .B2(\DP/ALU0/s_A_SHIFT[31] ), .A(n3950), .ZN(
        n4128) );
  AOI22_X1 U5106 ( .A1(n2424), .A2(n4128), .B1(n3951), .B2(n2426), .ZN(n3988)
         );
  AOI22_X1 U5107 ( .A1(n2427), .A2(n3988), .B1(n3952), .B2(n2429), .ZN(n3983)
         );
  XNOR2_X1 U5108 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[24] ), .ZN(n3974) );
  NOR3_X1 U5109 ( .A1(n3955), .A2(n3954), .A3(n3953), .ZN(n3957) );
  AOI21_X1 U5110 ( .B1(n3958), .B2(n3957), .A(n3956), .ZN(n3965) );
  OAI221_X1 U5111 ( .B1(n3962), .B2(n3961), .C1(n3962), .C2(n3960), .A(n3959), 
        .ZN(n3964) );
  OAI221_X1 U5112 ( .B1(n3966), .B2(n3965), .C1(n3966), .C2(n3964), .A(n3963), 
        .ZN(n3973) );
  AOI22_X1 U5113 ( .A1(n4016), .A2(n2431), .B1(n4164), .B2(
        \DP/ALU0/S_B_LHI[8] ), .ZN(n3972) );
  NOR2_X1 U5114 ( .A1(n27), .A2(n5), .ZN(n3967) );
  AOI211_X1 U5115 ( .C1(n27), .C2(n5), .A(n3967), .B(n4178), .ZN(n3969) );
  NOR3_X1 U5116 ( .A1(n27), .A2(n5), .A3(n4239), .ZN(n3968) );
  AOI211_X1 U5117 ( .C1(n3970), .C2(n2432), .A(n3969), .B(n3968), .ZN(n3971)
         );
  OAI211_X1 U5118 ( .C1(n4175), .C2(n3983), .A(n3972), .B(n3971), .ZN(
        \DP/RegALU1/N27 ) );
  XNOR2_X1 U5119 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[25] ), .ZN(n3990) );
  FA_X1 U5120 ( .A(\DP/ALU0/s_A_ADDER[24] ), .B(n3974), .CI(n3973), .CO(n3989), 
        .S(n4016) );
  AOI22_X1 U5121 ( .A1(n4006), .A2(n2430), .B1(n4164), .B2(
        \DP/ALU0/S_B_LHI[9] ), .ZN(n3982) );
  AOI22_X1 U5122 ( .A1(\DP/ALU0/s_A_SHIFT[9] ), .A2(n4168), .B1(n4152), .B2(
        \DP/ALU0/s_A_SHIFT[25] ), .ZN(n3975) );
  OAI211_X1 U5123 ( .C1(n18), .C2(n4150), .A(n3975), .B(n4124), .ZN(n4140) );
  AOI22_X1 U5124 ( .A1(n2424), .A2(n4140), .B1(n3976), .B2(n4205), .ZN(n4117)
         );
  AOI22_X1 U5125 ( .A1(n2428), .A2(n4117), .B1(n3977), .B2(n2429), .ZN(n3994)
         );
  NOR2_X1 U5126 ( .A1(n32), .A2(n4), .ZN(n3978) );
  AOI211_X1 U5127 ( .C1(n32), .C2(n4), .A(n3978), .B(n4178), .ZN(n3980) );
  NOR3_X1 U5128 ( .A1(n32), .A2(n4), .A3(n4239), .ZN(n3979) );
  AOI211_X1 U5129 ( .C1(n3994), .C2(n4234), .A(n3980), .B(n3979), .ZN(n3981)
         );
  OAI211_X1 U5130 ( .C1(n2396), .C2(n3983), .A(n3982), .B(n3981), .ZN(
        \DP/RegALU1/N28 ) );
  INV_X1 U5131 ( .A(n4124), .ZN(n3986) );
  INV_X1 U5132 ( .A(\DP/ALU0/s_A_SHIFT[10] ), .ZN(n3984) );
  OAI22_X1 U5133 ( .A1(n15), .A2(n4150), .B1(n3984), .B2(n4148), .ZN(n3985) );
  AOI211_X1 U5134 ( .C1(n4152), .C2(\DP/ALU0/s_A_SHIFT[26] ), .A(n3986), .B(
        n3985), .ZN(n4154) );
  AOI22_X1 U5135 ( .A1(n2424), .A2(n4154), .B1(n3987), .B2(n4205), .ZN(n4129)
         );
  AOI22_X1 U5136 ( .A1(n2427), .A2(n4129), .B1(n3988), .B2(n2429), .ZN(n4123)
         );
  XNOR2_X1 U5137 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[26] ), .ZN(n4022) );
  FA_X1 U5138 ( .A(\DP/ALU0/s_A_ADDER[25] ), .B(n3990), .CI(n3989), .CO(n4021), 
        .S(n4006) );
  AOI22_X1 U5139 ( .A1(n4007), .A2(n2430), .B1(n4164), .B2(
        \DP/ALU0/S_B_LHI[10] ), .ZN(n3996) );
  NOR2_X1 U5140 ( .A1(n40), .A2(n39), .ZN(n3991) );
  AOI211_X1 U5141 ( .C1(n40), .C2(n39), .A(n3991), .B(n4178), .ZN(n3993) );
  NOR3_X1 U5142 ( .A1(n40), .A2(n39), .A3(n4239), .ZN(n3992) );
  AOI211_X1 U5143 ( .C1(n3994), .C2(n2432), .A(n3993), .B(n3992), .ZN(n3995)
         );
  OAI211_X1 U5144 ( .C1(n4175), .C2(n4123), .A(n3996), .B(n3995), .ZN(
        \DP/RegALU1/N29 ) );
  INV_X1 U5145 ( .A(n3997), .ZN(n4055) );
  NOR4_X1 U5146 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(n4020)
         );
  NOR4_X1 U5147 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4019)
         );
  NOR4_X1 U5148 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4018)
         );
  FA_X1 U5149 ( .A(\DP/ALU0/s_A_ADDER[5] ), .B(n4011), .CI(n4010), .CO(n4013), 
        .S(n4222) );
  FA_X1 U5150 ( .A(\DP/ALU0/s_A_ADDER[6] ), .B(n4013), .CI(n4012), .CO(n3719), 
        .S(n4232) );
  XOR2_X1 U5151 ( .A(n4014), .B(\DP/ALU0/s_A_ADDER[0] ), .Z(n4102) );
  INV_X1 U5152 ( .A(n4102), .ZN(n4015) );
  NOR4_X1 U5153 ( .A1(n4222), .A2(n4232), .A3(n4016), .A4(n4015), .ZN(n4017)
         );
  NAND4_X1 U5154 ( .A1(n4020), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(n4048)
         );
  XNOR2_X1 U5155 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[30] ), .ZN(n4027) );
  XNOR2_X1 U5156 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[29] ), .ZN(n4023) );
  XNOR2_X1 U5157 ( .A(n2450), .B(\DP/ALU0/S_B_ADDER[28] ), .ZN(n4041) );
  AOI22_X1 U5158 ( .A1(\DP/ALU0/s_A_ADDER[29] ), .A2(n4023), .B1(
        \DP/ALU0/s_A_ADDER[28] ), .B2(n4041), .ZN(n4025) );
  XNOR2_X1 U5159 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[27] ), .ZN(n4029) );
  FA_X1 U5160 ( .A(\DP/ALU0/s_A_ADDER[26] ), .B(n4022), .CI(n4021), .CO(n4028), 
        .S(n4007) );
  OAI21_X1 U5161 ( .B1(\DP/ALU0/s_A_ADDER[28] ), .B2(n4041), .A(n4040), .ZN(
        n4024) );
  INV_X1 U5162 ( .A(n4023), .ZN(n4038) );
  INV_X1 U5163 ( .A(\DP/ALU0/s_A_ADDER[29] ), .ZN(n4039) );
  AOI22_X1 U5164 ( .A1(n4025), .A2(n4024), .B1(n4038), .B2(n4039), .ZN(n4026)
         );
  XNOR2_X1 U5165 ( .A(n57), .B(\DP/ALU0/S_B_ADDER[31] ), .ZN(n4062) );
  FA_X1 U5166 ( .A(\DP/ALU0/s_A_ADDER[30] ), .B(n4027), .CI(n4026), .CO(n4063), 
        .S(n4157) );
  FA_X1 U5167 ( .A(\DP/ALU0/s_A_ADDER[27] ), .B(n4029), .CI(n4028), .CO(n4040), 
        .S(n4114) );
  NOR4_X1 U5168 ( .A1(n4165), .A2(n4157), .A3(n4130), .A4(n4114), .ZN(n4046)
         );
  FA_X1 U5169 ( .A(\DP/ALU0/s_A_ADDER[4] ), .B(n4031), .CI(n4030), .CO(n4010), 
        .S(n4214) );
  FA_X1 U5170 ( .A(\DP/ALU0/s_A_ADDER[3] ), .B(n4033), .CI(n4032), .CO(n4030), 
        .S(n4204) );
  FA_X1 U5171 ( .A(\DP/ALU0/s_A_ADDER[2] ), .B(n4035), .CI(n4034), .CO(n4032), 
        .S(n4195) );
  FA_X1 U5172 ( .A(\DP/ALU0/s_A_ADDER[1] ), .B(n4037), .CI(n4036), .CO(n4034), 
        .S(n4186) );
  NOR4_X1 U5173 ( .A1(n4214), .A2(n4204), .A3(n4195), .A4(n4186), .ZN(n4045)
         );
  XOR2_X1 U5174 ( .A(n4039), .B(n4038), .Z(n4043) );
  FA_X1 U5175 ( .A(\DP/ALU0/s_A_ADDER[28] ), .B(n4041), .CI(n4040), .CO(n4042), 
        .S(n4130) );
  XOR2_X1 U5176 ( .A(n4043), .B(n4042), .Z(n4137) );
  INV_X1 U5177 ( .A(n4137), .ZN(n4044) );
  NAND3_X1 U5178 ( .A1(n4046), .A2(n4045), .A3(n4044), .ZN(n4047) );
  NOR4_X1 U5179 ( .A1(n4050), .A2(n4049), .A3(n4048), .A4(n4047), .ZN(n4053)
         );
  INV_X1 U5180 ( .A(n4051), .ZN(n4052) );
  NAND4_X1 U5181 ( .A1(n4055), .A2(n4054), .A3(n4053), .A4(n4052), .ZN(n4056)
         );
  NOR3_X1 U5182 ( .A1(n4058), .A2(n4057), .A3(n4056), .ZN(n4071) );
  NOR2_X1 U5183 ( .A1(w_ALU_OPCODE[2]), .A2(n4103), .ZN(n4061) );
  OAI211_X1 U5184 ( .C1(n4103), .C2(n2362), .A(n4059), .B(n4071), .ZN(n4060)
         );
  OAI21_X1 U5185 ( .B1(n4071), .B2(n4061), .A(n4060), .ZN(n4113) );
  FA_X1 U5186 ( .A(\DP/ALU0/s_A_ADDER[31] ), .B(n4063), .CI(n4062), .CO(n4064), 
        .S(n4165) );
  XOR2_X1 U5187 ( .A(\DP/ALU0/s_SIGN ), .B(n4064), .Z(n4111) );
  AOI21_X1 U5188 ( .B1(n4744), .B2(n4066), .A(n4065), .ZN(n4070) );
  NOR2_X1 U5189 ( .A1(n4744), .A2(n4067), .ZN(n4106) );
  AOI21_X1 U5190 ( .B1(n218), .B2(n4106), .A(n4068), .ZN(n4069) );
  OAI21_X1 U5191 ( .B1(n4071), .B2(n4070), .A(n4069), .ZN(n4110) );
  NAND2_X1 U5192 ( .A1(\DP/ALU0/S_B_LOGIC[0] ), .A2(\DP/ALU0/s_A_LOGIC[0] ), 
        .ZN(n4074) );
  OAI21_X1 U5193 ( .B1(\DP/ALU0/S_B_LOGIC[0] ), .B2(\DP/ALU0/s_A_LOGIC[0] ), 
        .A(\DP/ALU0/s_LOGIC[2] ), .ZN(n4072) );
  OAI21_X1 U5195 ( .B1(\DP/ALU0/s_LOGIC[3] ), .B2(n4074), .A(n4073), .ZN(n4100) );
  OAI222_X1 U5196 ( .A1(n4149), .A2(n4092), .B1(n4091), .B2(n22), .C1(n4090), 
        .C2(n4075), .ZN(n4206) );
  AOI22_X1 U5197 ( .A1(n4083), .A2(\DP/ALU0/s_A_SHIFT[2] ), .B1(n4082), .B2(
        \DP/ALU0/s_A_SHIFT[10] ), .ZN(n4076) );
  OAI21_X1 U5198 ( .B1(n15), .B2(n4091), .A(n4076), .ZN(n4077) );
  AOI22_X1 U5199 ( .A1(n2424), .A2(n4206), .B1(n4077), .B2(n2426), .ZN(n4189)
         );
  OAI222_X1 U5200 ( .A1(n4125), .A2(n4092), .B1(n4091), .B2(n20), .C1(n4090), 
        .C2(n4078), .ZN(n4187) );
  AOI22_X1 U5201 ( .A1(\DP/ALU0/s_A_SHIFT[0] ), .A2(n4083), .B1(n4082), .B2(
        \DP/ALU0/s_A_SHIFT[8] ), .ZN(n4079) );
  OAI21_X1 U5202 ( .B1(n13), .B2(n4091), .A(n4079), .ZN(n4080) );
  AOI22_X1 U5203 ( .A1(n2424), .A2(n4187), .B1(n4080), .B2(n2426), .ZN(n4081)
         );
  AOI22_X1 U5204 ( .A1(n2427), .A2(n4189), .B1(n4081), .B2(n2429), .ZN(n4097)
         );
  AOI22_X1 U5205 ( .A1(n4083), .A2(\DP/ALU0/s_A_SHIFT[3] ), .B1(n4082), .B2(
        \DP/ALU0/s_A_SHIFT[11] ), .ZN(n4084) );
  OAI21_X1 U5206 ( .B1(n45), .B2(n4091), .A(n4084), .ZN(n4085) );
  AOI22_X1 U5207 ( .A1(n2424), .A2(n4086), .B1(n4085), .B2(n2426), .ZN(n4198)
         );
  OAI222_X1 U5208 ( .A1(n4088), .A2(n4092), .B1(n4091), .B2(n25), .C1(n4090), 
        .C2(n4087), .ZN(n4196) );
  OAI222_X1 U5209 ( .A1(n4093), .A2(n4092), .B1(n4091), .B2(n18), .C1(n4090), 
        .C2(n4089), .ZN(n4094) );
  AOI22_X1 U5210 ( .A1(n2424), .A2(n4196), .B1(n4094), .B2(n2426), .ZN(n4095)
         );
  AOI22_X1 U5211 ( .A1(n2427), .A2(n4198), .B1(n4095), .B2(n2429), .ZN(n4190)
         );
  OAI221_X1 U5212 ( .B1(n4098), .B2(n4097), .C1(n4096), .C2(n4190), .A(n2445), 
        .ZN(n4099) );
  OAI211_X1 U5213 ( .C1(n4102), .C2(n4101), .A(n4100), .B(n4099), .ZN(n4109)
         );
  NOR2_X1 U5214 ( .A1(n2362), .A2(n4103), .ZN(n4105) );
  AOI211_X1 U5215 ( .C1(n4106), .C2(n2363), .A(n4105), .B(n4104), .ZN(n4107)
         );
  NOR2_X1 U5216 ( .A1(n4107), .A2(n4111), .ZN(n4108) );
  AOI211_X1 U5217 ( .C1(n4111), .C2(n4110), .A(n4109), .B(n4108), .ZN(n4112)
         );
  AOI21_X1 U5218 ( .B1(n4113), .B2(n4112), .A(n2461), .ZN(\DP/RegALU1/N3 ) );
  AOI22_X1 U5219 ( .A1(n4114), .A2(n2430), .B1(n4164), .B2(
        \DP/ALU0/S_B_LHI[11] ), .ZN(n4122) );
  AOI22_X1 U5220 ( .A1(\DP/ALU0/s_A_SHIFT[11] ), .A2(n4168), .B1(n4152), .B2(
        \DP/ALU0/s_A_SHIFT[27] ), .ZN(n4115) );
  OAI211_X1 U5221 ( .C1(n45), .C2(n4150), .A(n4115), .B(n4124), .ZN(n4174) );
  AOI22_X1 U5222 ( .A1(n2424), .A2(n4174), .B1(n4116), .B2(n4205), .ZN(n4141)
         );
  AOI22_X1 U5223 ( .A1(n2427), .A2(n4141), .B1(n4117), .B2(n2429), .ZN(n4134)
         );
  NOR2_X1 U5224 ( .A1(n38), .A2(n37), .ZN(n4118) );
  AOI211_X1 U5225 ( .C1(n38), .C2(n37), .A(n4118), .B(n4178), .ZN(n4120) );
  NOR3_X1 U5226 ( .A1(n38), .A2(n37), .A3(n4239), .ZN(n4119) );
  AOI211_X1 U5227 ( .C1(n4134), .C2(n4234), .A(n4120), .B(n4119), .ZN(n4121)
         );
  OAI211_X1 U5228 ( .C1(n2396), .C2(n4123), .A(n4122), .B(n4121), .ZN(
        \DP/RegALU1/N30 ) );
  NAND2_X1 U5229 ( .A1(n2424), .A2(n4124), .ZN(n4172) );
  OAI22_X1 U5230 ( .A1(n20), .A2(n4150), .B1(n4125), .B2(n4148), .ZN(n4126) );
  AOI211_X1 U5231 ( .C1(n4152), .C2(\DP/ALU0/s_A_SHIFT[28] ), .A(n4172), .B(
        n4126), .ZN(n4127) );
  AOI21_X1 U5232 ( .B1(n4128), .B2(n4205), .A(n4127), .ZN(n4155) );
  AOI22_X1 U5233 ( .A1(n2427), .A2(n4155), .B1(n4129), .B2(n4223), .ZN(n4147)
         );
  AOI22_X1 U5234 ( .A1(n4130), .A2(n2430), .B1(n4164), .B2(
        \DP/ALU0/S_B_LHI[12] ), .ZN(n4136) );
  NOR2_X1 U5235 ( .A1(n33), .A2(n3), .ZN(n4131) );
  AOI211_X1 U5236 ( .C1(n33), .C2(n3), .A(n4131), .B(n4178), .ZN(n4133) );
  NOR3_X1 U5237 ( .A1(n33), .A2(n3), .A3(n2433), .ZN(n4132) );
  AOI211_X1 U5238 ( .C1(n4134), .C2(n2432), .A(n4133), .B(n4132), .ZN(n4135)
         );
  OAI211_X1 U5239 ( .C1(n4147), .C2(n4175), .A(n4136), .B(n4135), .ZN(
        \DP/RegALU1/N31 ) );
  AOI22_X1 U5240 ( .A1(n4137), .A2(n2430), .B1(n4164), .B2(
        \DP/ALU0/S_B_LHI[13] ), .ZN(n4146) );
  AOI22_X1 U5241 ( .A1(\DP/ALU0/s_A_SHIFT[13] ), .A2(n4168), .B1(n4152), .B2(
        \DP/ALU0/s_A_SHIFT[29] ), .ZN(n4138) );
  OAI21_X1 U5242 ( .B1(n25), .B2(n4150), .A(n4138), .ZN(n4139) );
  OAI22_X1 U5243 ( .A1(n2424), .A2(n4140), .B1(n4139), .B2(n4172), .ZN(n4176)
         );
  AOI22_X1 U5244 ( .A1(n2427), .A2(n4176), .B1(n4141), .B2(n4223), .ZN(n4161)
         );
  NOR2_X1 U5245 ( .A1(n36), .A2(n35), .ZN(n4142) );
  AOI211_X1 U5246 ( .C1(n36), .C2(n35), .A(n4142), .B(n4178), .ZN(n4144) );
  NOR3_X1 U5247 ( .A1(n36), .A2(n35), .A3(n2433), .ZN(n4143) );
  AOI211_X1 U5248 ( .C1(n4234), .C2(n4161), .A(n4144), .B(n4143), .ZN(n4145)
         );
  OAI211_X1 U5249 ( .C1(n4147), .C2(n2396), .A(n4146), .B(n4145), .ZN(
        \DP/RegALU1/N32 ) );
  OAI22_X1 U5250 ( .A1(n22), .A2(n4150), .B1(n4149), .B2(n4148), .ZN(n4151) );
  AOI211_X1 U5251 ( .C1(n4152), .C2(\DP/ALU0/s_A_SHIFT[30] ), .A(n4172), .B(
        n4151), .ZN(n4153) );
  AOI21_X1 U5252 ( .B1(n4154), .B2(n2426), .A(n4153), .ZN(n4156) );
  AOI22_X1 U5253 ( .A1(n2427), .A2(n4156), .B1(n4155), .B2(n4223), .ZN(n4184)
         );
  AOI22_X1 U5254 ( .A1(n4157), .A2(n2430), .B1(n4164), .B2(
        \DP/ALU0/S_B_LHI[14] ), .ZN(n4163) );
  NOR2_X1 U5255 ( .A1(n34), .A2(n2), .ZN(n4158) );
  AOI211_X1 U5256 ( .C1(n34), .C2(n2), .A(n4158), .B(n4178), .ZN(n4160) );
  NOR3_X1 U5257 ( .A1(n34), .A2(n2), .A3(n4239), .ZN(n4159) );
  AOI211_X1 U5258 ( .C1(n2432), .C2(n4161), .A(n4160), .B(n4159), .ZN(n4162)
         );
  OAI211_X1 U5259 ( .C1(n4184), .C2(n4175), .A(n4163), .B(n4162), .ZN(
        \DP/RegALU1/N33 ) );
  AOI22_X1 U5260 ( .A1(n4165), .A2(n2430), .B1(n4164), .B2(
        \DP/ALU0/S_B_LHI[15] ), .ZN(n4183) );
  NOR2_X1 U5261 ( .A1(n56), .A2(n1), .ZN(n4181) );
  AOI22_X1 U5262 ( .A1(n4168), .A2(\DP/ALU0/s_A_SHIFT[15] ), .B1(n4167), .B2(
        n4166), .ZN(n4169) );
  OAI21_X1 U5263 ( .B1(n4171), .B2(n4170), .A(n4169), .ZN(n4173) );
  OAI22_X1 U5264 ( .A1(n2425), .A2(n4174), .B1(n4173), .B2(n4172), .ZN(n4177)
         );
  AOI221_X1 U5265 ( .B1(n2428), .B2(n4177), .C1(n4223), .C2(n4176), .A(n4175), 
        .ZN(n4180) );
  AOI211_X1 U5266 ( .C1(n56), .C2(n1), .A(n4181), .B(n4178), .ZN(n4179) );
  AOI211_X1 U5267 ( .C1(n2434), .C2(n4181), .A(n4180), .B(n4179), .ZN(n4182)
         );
  OAI211_X1 U5268 ( .C1(n4184), .C2(n2396), .A(n4183), .B(n4182), .ZN(
        \DP/RegALU1/N34 ) );
  NAND2_X1 U5269 ( .A1(\DP/ALU0/s_A_LOGIC[1] ), .A2(\DP/ALU0/S_B_LOGIC[1] ), 
        .ZN(n4193) );
  XOR2_X1 U5270 ( .A(\DP/ALU0/s_A_LOGIC[1] ), .B(\DP/ALU0/S_B_LOGIC[1] ), .Z(
        n4185) );
  AOI22_X1 U5271 ( .A1(n4186), .A2(n2430), .B1(n4231), .B2(n4185), .ZN(n4192)
         );
  AOI22_X1 U5272 ( .A1(n2424), .A2(n4188), .B1(n4187), .B2(n2426), .ZN(n4208)
         );
  AOI22_X1 U5273 ( .A1(n2427), .A2(n4208), .B1(n4189), .B2(n4223), .ZN(n4199)
         );
  AOI22_X1 U5274 ( .A1(n4234), .A2(n4199), .B1(n2432), .B2(n4190), .ZN(n4191)
         );
  OAI211_X1 U5275 ( .C1(n2433), .C2(n4193), .A(n4192), .B(n4191), .ZN(
        \DP/RegALU1/N4 ) );
  NAND2_X1 U5276 ( .A1(\DP/ALU0/s_A_LOGIC[2] ), .A2(\DP/ALU0/S_B_LOGIC[2] ), 
        .ZN(n4202) );
  XOR2_X1 U5277 ( .A(\DP/ALU0/s_A_LOGIC[2] ), .B(\DP/ALU0/S_B_LOGIC[2] ), .Z(
        n4194) );
  AOI22_X1 U5278 ( .A1(n4195), .A2(n2430), .B1(n4231), .B2(n4194), .ZN(n4201)
         );
  AOI22_X1 U5279 ( .A1(n2424), .A2(n4197), .B1(n4196), .B2(n4205), .ZN(n4215)
         );
  AOI22_X1 U5280 ( .A1(n2427), .A2(n4215), .B1(n4198), .B2(n2429), .ZN(n4209)
         );
  AOI22_X1 U5281 ( .A1(n2432), .A2(n4199), .B1(n4234), .B2(n4209), .ZN(n4200)
         );
  OAI211_X1 U5282 ( .C1(n2433), .C2(n4202), .A(n4201), .B(n4200), .ZN(
        \DP/RegALU1/N5 ) );
  NAND2_X1 U5283 ( .A1(\DP/ALU0/s_A_LOGIC[3] ), .A2(\DP/ALU0/S_B_LOGIC[3] ), 
        .ZN(n4212) );
  XOR2_X1 U5284 ( .A(\DP/ALU0/s_A_LOGIC[3] ), .B(\DP/ALU0/S_B_LOGIC[3] ), .Z(
        n4203) );
  AOI22_X1 U5285 ( .A1(n4204), .A2(n2430), .B1(n4231), .B2(n4203), .ZN(n4211)
         );
  AOI22_X1 U5286 ( .A1(n2425), .A2(n4207), .B1(n4206), .B2(n2426), .ZN(n4224)
         );
  AOI22_X1 U5287 ( .A1(n2427), .A2(n4224), .B1(n4208), .B2(n2429), .ZN(n4217)
         );
  AOI22_X1 U5288 ( .A1(n2432), .A2(n4209), .B1(n4234), .B2(n4217), .ZN(n4210)
         );
  OAI211_X1 U5289 ( .C1(n4239), .C2(n4212), .A(n4211), .B(n4210), .ZN(
        \DP/RegALU1/N6 ) );
  NAND2_X1 U5290 ( .A1(\DP/ALU0/s_A_LOGIC[4] ), .A2(\DP/ALU0/S_B_LOGIC[4] ), 
        .ZN(n4220) );
  XOR2_X1 U5291 ( .A(\DP/ALU0/s_A_LOGIC[4] ), .B(\DP/ALU0/S_B_LOGIC[4] ), .Z(
        n4213) );
  AOI22_X1 U5292 ( .A1(n4214), .A2(n2430), .B1(n4231), .B2(n4213), .ZN(n4219)
         );
  AOI22_X1 U5293 ( .A1(n2427), .A2(n4216), .B1(n4215), .B2(n2429), .ZN(n4226)
         );
  AOI22_X1 U5294 ( .A1(n2432), .A2(n4217), .B1(n4234), .B2(n4226), .ZN(n4218)
         );
  OAI211_X1 U5295 ( .C1(n4239), .C2(n4220), .A(n4219), .B(n4218), .ZN(
        \DP/RegALU1/N7 ) );
  NAND2_X1 U5296 ( .A1(\DP/ALU0/s_A_LOGIC[5] ), .A2(\DP/ALU0/S_B_LOGIC[5] ), 
        .ZN(n4229) );
  XOR2_X1 U5297 ( .A(\DP/ALU0/s_A_LOGIC[5] ), .B(\DP/ALU0/S_B_LOGIC[5] ), .Z(
        n4221) );
  AOI22_X1 U5298 ( .A1(n4222), .A2(n2430), .B1(n4231), .B2(n4221), .ZN(n4228)
         );
  AOI22_X1 U5299 ( .A1(n2428), .A2(n4225), .B1(n4224), .B2(n2429), .ZN(n4235)
         );
  AOI22_X1 U5300 ( .A1(n2432), .A2(n4226), .B1(n4234), .B2(n4235), .ZN(n4227)
         );
  OAI211_X1 U5301 ( .C1(n2433), .C2(n4229), .A(n4228), .B(n4227), .ZN(
        \DP/RegALU1/N8 ) );
  NAND2_X1 U5302 ( .A1(\DP/ALU0/s_A_LOGIC[6] ), .A2(\DP/ALU0/S_B_LOGIC[6] ), 
        .ZN(n4238) );
  XOR2_X1 U5303 ( .A(\DP/ALU0/s_A_LOGIC[6] ), .B(\DP/ALU0/S_B_LOGIC[6] ), .Z(
        n4230) );
  AOI22_X1 U5304 ( .A1(n4232), .A2(n2430), .B1(n4231), .B2(n4230), .ZN(n4237)
         );
  AOI22_X1 U5305 ( .A1(n2432), .A2(n4235), .B1(n4234), .B2(n4233), .ZN(n4236)
         );
  OAI211_X1 U5306 ( .C1(n2433), .C2(n4238), .A(n4237), .B(n4236), .ZN(
        \DP/RegALU1/N9 ) );
  AND2_X1 U5307 ( .A1(RST), .A2(\DP/RegB_in[7] ), .ZN(\DP/RegB/N10 ) );
  AND2_X1 U5308 ( .A1(RST), .A2(\DP/RegB_in[8] ), .ZN(\DP/RegB/N11 ) );
  AND2_X1 U5309 ( .A1(RST), .A2(\DP/RegB_in[9] ), .ZN(\DP/RegB/N12 ) );
  AND2_X1 U5310 ( .A1(RST), .A2(\DP/RegB_in[10] ), .ZN(\DP/RegB/N13 ) );
  AND2_X1 U5311 ( .A1(RST), .A2(\DP/RegB_in[11] ), .ZN(\DP/RegB/N14 ) );
  AND2_X1 U5312 ( .A1(RST), .A2(\DP/RegB_in[12] ), .ZN(\DP/RegB/N15 ) );
  AND2_X1 U5313 ( .A1(RST), .A2(\DP/RegB_in[13] ), .ZN(\DP/RegB/N16 ) );
  AND2_X1 U5314 ( .A1(RST), .A2(\DP/RegB_in[14] ), .ZN(\DP/RegB/N17 ) );
  AND2_X1 U5315 ( .A1(RST), .A2(\DP/RegB_in[15] ), .ZN(\DP/RegB/N18 ) );
  AND2_X1 U5316 ( .A1(RST), .A2(\DP/RegB_in[16] ), .ZN(\DP/RegB/N19 ) );
  OR2_X1 U5317 ( .A1(n2461), .A2(n66), .ZN(\DP/RegB/N2 ) );
  AND2_X1 U5318 ( .A1(RST), .A2(\DP/RegB_in[17] ), .ZN(\DP/RegB/N20 ) );
  AND2_X1 U5319 ( .A1(RST), .A2(\DP/RegB_in[18] ), .ZN(\DP/RegB/N21 ) );
  AND2_X1 U5320 ( .A1(RST), .A2(\DP/RegB_in[19] ), .ZN(\DP/RegB/N22 ) );
  AND2_X1 U5321 ( .A1(RST), .A2(\DP/RegB_in[20] ), .ZN(\DP/RegB/N23 ) );
  AND2_X1 U5322 ( .A1(RST), .A2(\DP/RegB_in[21] ), .ZN(\DP/RegB/N24 ) );
  AND2_X1 U5323 ( .A1(RST), .A2(\DP/RegB_in[22] ), .ZN(\DP/RegB/N25 ) );
  AND2_X1 U5324 ( .A1(RST), .A2(\DP/RegB_in[23] ), .ZN(\DP/RegB/N26 ) );
  AND2_X1 U5325 ( .A1(RST), .A2(\DP/RegB_in[24] ), .ZN(\DP/RegB/N27 ) );
  AND2_X1 U5326 ( .A1(RST), .A2(\DP/RegB_in[25] ), .ZN(\DP/RegB/N28 ) );
  AND2_X1 U5327 ( .A1(RST), .A2(\DP/RegB_in[26] ), .ZN(\DP/RegB/N29 ) );
  AND2_X1 U5328 ( .A1(RST), .A2(\DP/RegB_in[0] ), .ZN(\DP/RegB/N3 ) );
  AND2_X1 U5329 ( .A1(RST), .A2(\DP/RegB_in[27] ), .ZN(\DP/RegB/N30 ) );
  AND2_X1 U5330 ( .A1(RST), .A2(\DP/RegB_in[28] ), .ZN(\DP/RegB/N31 ) );
  AND2_X1 U5331 ( .A1(RST), .A2(\DP/RegB_in[29] ), .ZN(\DP/RegB/N32 ) );
  AND2_X1 U5332 ( .A1(RST), .A2(\DP/RegB_in[30] ), .ZN(\DP/RegB/N33 ) );
  AND2_X1 U5333 ( .A1(RST), .A2(\DP/RegB_in[31] ), .ZN(\DP/RegB/N34 ) );
  AND2_X1 U5334 ( .A1(RST), .A2(\DP/RegB_in[1] ), .ZN(\DP/RegB/N4 ) );
  AND2_X1 U5335 ( .A1(RST), .A2(\DP/RegB_in[2] ), .ZN(\DP/RegB/N5 ) );
  AND2_X1 U5336 ( .A1(RST), .A2(\DP/RegB_in[3] ), .ZN(\DP/RegB/N6 ) );
  AND2_X1 U5337 ( .A1(RST), .A2(\DP/RegB_in[4] ), .ZN(\DP/RegB/N7 ) );
  AND2_X1 U5338 ( .A1(RST), .A2(\DP/RegB_in[5] ), .ZN(\DP/RegB/N8 ) );
  AND2_X1 U5339 ( .A1(RST), .A2(\DP/RegB_in[6] ), .ZN(\DP/RegB/N9 ) );
  OR4_X1 U5344 ( .A1(\DP/RD1[1] ), .A2(\DP/RD1[0] ), .A3(\DP/RD1[4] ), .A4(
        \DP/RD1[3] ), .ZN(n4240) );
  OAI21_X1 U5345 ( .B1(\DP/RD1[2] ), .B2(n4240), .A(w_RF_WE_EX), .ZN(n4260) );
  OAI22_X1 U5347 ( .A1(n4267), .A2(\DP/RD1[0] ), .B1(n4272), .B2(\DP/RD1[4] ), 
        .ZN(n4242) );
  AOI221_X1 U5348 ( .B1(n4267), .B2(\DP/RD1[0] ), .C1(\DP/RD1[4] ), .C2(n4272), 
        .A(n4242), .ZN(n4243) );
  NOR2_X1 U5352 ( .A1(n4260), .A2(n4246), .ZN(n4255) );
  OAI221_X1 U5354 ( .B1(n104), .B2(n401), .C1(n4272), .C2(n2365), .A(n4247), 
        .ZN(n4252) );
  AOI22_X1 U5355 ( .A1(n103), .A2(n400), .B1(n4267), .B2(\DP/RD2[0] ), .ZN(
        n4248) );
  OAI221_X1 U5356 ( .B1(n103), .B2(n400), .C1(n4267), .C2(\DP/RD2[0] ), .A(
        n4248), .ZN(n4251) );
  AOI22_X1 U5357 ( .A1(n4269), .A2(\DP/RD2[2] ), .B1(n4268), .B2(\DP/RD2[1] ), 
        .ZN(n4249) );
  OAI221_X1 U5358 ( .B1(n4269), .B2(\DP/RD2[2] ), .C1(n4268), .C2(\DP/RD2[1] ), 
        .A(n4249), .ZN(n4250) );
  NOR3_X1 U5360 ( .A1(n4255), .A2(n4254), .A3(n2460), .ZN(\DP/RegFC/N3 ) );
  AND2_X1 U5361 ( .A1(RST), .A2(n4254), .ZN(\DP/RegFC/N4 ) );
  AND2_X1 U5362 ( .A1(RST), .A2(n4255), .ZN(\DP/RegFC/N5 ) );
  OAI22_X1 U5363 ( .A1(n4419), .A2(\DP/RD1[0] ), .B1(n4424), .B2(\DP/RD1[4] ), 
        .ZN(n4256) );
  AOI221_X1 U5364 ( .B1(n4419), .B2(\DP/RD1[0] ), .C1(\DP/RD1[4] ), .C2(n4424), 
        .A(n4256), .ZN(n4257) );
  NOR2_X1 U5368 ( .A1(n4260), .A2(n4261), .ZN(n4265) );
  INV_X1 U5369 ( .A(n4261), .ZN(n4263) );
  NOR2_X1 U5370 ( .A1(n4263), .A2(n4262), .ZN(n4264) );
  NOR3_X1 U5371 ( .A1(n4265), .A2(n4264), .A3(n2461), .ZN(\DP/RegFB/N3 ) );
  AND2_X1 U5372 ( .A1(RST), .A2(n4264), .ZN(\DP/RegFB/N4 ) );
  AND2_X1 U5373 ( .A1(RST), .A2(n4265), .ZN(\DP/RegFB/N5 ) );
  AND2_X1 U5374 ( .A1(IR_OUT[7]), .A2(n4275), .ZN(\DP/RegIMM/N10 ) );
  AND2_X1 U5375 ( .A1(IR_OUT[8]), .A2(n4275), .ZN(\DP/RegIMM/N11 ) );
  NOR2_X1 U5376 ( .A1(n2391), .A2(n4274), .ZN(\DP/RegIMM/N12 ) );
  AND2_X1 U5377 ( .A1(IR_OUT[10]), .A2(n4275), .ZN(\DP/RegIMM/N13 ) );
  NAND2_X1 U5378 ( .A1(n4275), .A2(IR_OUT[11]), .ZN(n584) );
  NAND2_X1 U5379 ( .A1(n4275), .A2(IR_OUT[12]), .ZN(n582) );
  NAND2_X1 U5380 ( .A1(n4275), .A2(IR_OUT[13]), .ZN(n580) );
  NAND2_X1 U5381 ( .A1(n4275), .A2(IR_OUT[14]), .ZN(n578) );
  NAND2_X1 U5382 ( .A1(n4275), .A2(IR_OUT[15]), .ZN(n575) );
  NAND3_X1 U5383 ( .A1(RST), .A2(IR_OUT[15]), .A3(n4266), .ZN(n4271) );
  OAI21_X1 U5384 ( .B1(n4273), .B2(n4419), .A(n4271), .ZN(\DP/RegIMM/N19 ) );
  OAI21_X1 U5385 ( .B1(n4273), .B2(n4420), .A(n4271), .ZN(\DP/RegIMM/N20 ) );
  OAI21_X1 U5386 ( .B1(n4273), .B2(n4421), .A(n4271), .ZN(\DP/RegIMM/N21 ) );
  OAI21_X1 U5387 ( .B1(n4273), .B2(n4422), .A(n4271), .ZN(\DP/RegIMM/N22 ) );
  OAI21_X1 U5388 ( .B1(n4273), .B2(n4424), .A(n4271), .ZN(\DP/RegIMM/N23 ) );
  OAI21_X1 U5389 ( .B1(n4273), .B2(n4267), .A(n4271), .ZN(\DP/RegIMM/N24 ) );
  OAI21_X1 U5390 ( .B1(n4273), .B2(n4268), .A(n4271), .ZN(\DP/RegIMM/N25 ) );
  OAI21_X1 U5391 ( .B1(n4273), .B2(n4269), .A(n4271), .ZN(\DP/RegIMM/N26 ) );
  OAI21_X1 U5392 ( .B1(n4273), .B2(n4270), .A(n4271), .ZN(\DP/RegIMM/N27 ) );
  OAI21_X1 U5393 ( .B1(n4273), .B2(n4272), .A(n4271), .ZN(\DP/RegIMM/N34 ) );
  NOR2_X1 U5394 ( .A1(n2382), .A2(n4274), .ZN(\DP/RegIMM/N4 ) );
  NOR2_X1 U5395 ( .A1(n2390), .A2(n4274), .ZN(\DP/RegIMM/N6 ) );
  AND2_X1 U5396 ( .A1(IR_OUT[4]), .A2(n4275), .ZN(\DP/RegIMM/N7 ) );
  AND2_X1 U5397 ( .A1(IR_OUT[6]), .A2(n4275), .ZN(\DP/RegIMM/N9 ) );
  NOR4_X1 U5398 ( .A1(w_LOAD_SIZE[2]), .A2(n2400), .A3(n2461), .A4(n2369), 
        .ZN(n4287) );
  NAND4_X1 U5399 ( .A1(n202), .A2(RST), .A3(w_LOAD_SIZE[2]), .A4(n2369), .ZN(
        n4276) );
  NAND2_X1 U5400 ( .A1(n4286), .A2(n4276), .ZN(n4308) );
  AND2_X1 U5401 ( .A1(\DP/LOAD8[7] ), .A2(n4308), .ZN(\DP/RegLMD/N10 ) );
  INV_X1 U5402 ( .A(\DP/LOAD16[8] ), .ZN(n4278) );
  INV_X1 U5403 ( .A(n4276), .ZN(n4277) );
  OAI21_X1 U5404 ( .B1(n4286), .B2(n4278), .A(n4288), .ZN(\DP/RegLMD/N11 ) );
  INV_X1 U5405 ( .A(\DP/LOAD16[9] ), .ZN(n4279) );
  OAI21_X1 U5406 ( .B1(n4286), .B2(n4279), .A(n4288), .ZN(\DP/RegLMD/N12 ) );
  INV_X1 U5407 ( .A(\DP/LOAD16[10] ), .ZN(n4280) );
  OAI21_X1 U5408 ( .B1(n4286), .B2(n4280), .A(n4288), .ZN(\DP/RegLMD/N13 ) );
  INV_X1 U5409 ( .A(\DP/LOAD16[11] ), .ZN(n4281) );
  OAI21_X1 U5410 ( .B1(n4286), .B2(n4281), .A(n4288), .ZN(\DP/RegLMD/N14 ) );
  INV_X1 U5411 ( .A(\DP/LOAD16[12] ), .ZN(n4282) );
  OAI21_X1 U5412 ( .B1(n4286), .B2(n4282), .A(n4288), .ZN(\DP/RegLMD/N15 ) );
  INV_X1 U5413 ( .A(\DP/LOAD16[13] ), .ZN(n4283) );
  OAI21_X1 U5414 ( .B1(n4286), .B2(n4283), .A(n4288), .ZN(\DP/RegLMD/N16 ) );
  INV_X1 U5415 ( .A(\DP/LOAD16[14] ), .ZN(n4284) );
  OAI21_X1 U5416 ( .B1(n4286), .B2(n4284), .A(n4288), .ZN(\DP/RegLMD/N17 ) );
  INV_X1 U5417 ( .A(\DP/LOAD16[15] ), .ZN(n4285) );
  OAI21_X1 U5418 ( .B1(n4286), .B2(n4285), .A(n4288), .ZN(\DP/RegLMD/N18 ) );
  NAND3_X1 U5419 ( .A1(n4287), .A2(\DP/LOAD16[15] ), .A3(w_SIGN_LD), .ZN(n4289) );
  AOI21_X1 U5420 ( .B1(n4306), .B2(DRAM_DATA_IN[16]), .A(n4305), .ZN(n4290) );
  INV_X1 U5421 ( .A(n4290), .ZN(\DP/RegLMD/N19 ) );
  AOI21_X1 U5422 ( .B1(n4306), .B2(DRAM_DATA_IN[17]), .A(n4305), .ZN(n4291) );
  INV_X1 U5423 ( .A(n4291), .ZN(\DP/RegLMD/N20 ) );
  AOI21_X1 U5424 ( .B1(n4306), .B2(DRAM_DATA_IN[18]), .A(n4305), .ZN(n4292) );
  INV_X1 U5425 ( .A(n4292), .ZN(\DP/RegLMD/N21 ) );
  AOI21_X1 U5426 ( .B1(n4306), .B2(DRAM_DATA_IN[19]), .A(n4305), .ZN(n4293) );
  INV_X1 U5427 ( .A(n4293), .ZN(\DP/RegLMD/N22 ) );
  AOI21_X1 U5428 ( .B1(n4306), .B2(DRAM_DATA_IN[20]), .A(n4305), .ZN(n4294) );
  INV_X1 U5429 ( .A(n4294), .ZN(\DP/RegLMD/N23 ) );
  AOI21_X1 U5430 ( .B1(n4306), .B2(DRAM_DATA_IN[21]), .A(n4305), .ZN(n4295) );
  INV_X1 U5431 ( .A(n4295), .ZN(\DP/RegLMD/N24 ) );
  AOI21_X1 U5432 ( .B1(n4306), .B2(DRAM_DATA_IN[22]), .A(n4305), .ZN(n4296) );
  INV_X1 U5433 ( .A(n4296), .ZN(\DP/RegLMD/N25 ) );
  AOI21_X1 U5434 ( .B1(n4306), .B2(DRAM_DATA_IN[23]), .A(n4305), .ZN(n4297) );
  INV_X1 U5435 ( .A(n4297), .ZN(\DP/RegLMD/N26 ) );
  AOI21_X1 U5436 ( .B1(n4306), .B2(DRAM_DATA_IN[24]), .A(n4305), .ZN(n4298) );
  INV_X1 U5437 ( .A(n4298), .ZN(\DP/RegLMD/N27 ) );
  AOI21_X1 U5438 ( .B1(n4306), .B2(DRAM_DATA_IN[25]), .A(n4305), .ZN(n4299) );
  INV_X1 U5439 ( .A(n4299), .ZN(\DP/RegLMD/N28 ) );
  AOI21_X1 U5440 ( .B1(n4306), .B2(DRAM_DATA_IN[26]), .A(n4305), .ZN(n4300) );
  INV_X1 U5441 ( .A(n4300), .ZN(\DP/RegLMD/N29 ) );
  AND2_X1 U5442 ( .A1(\DP/LOAD8[0] ), .A2(n4308), .ZN(\DP/RegLMD/N3 ) );
  AOI21_X1 U5443 ( .B1(n4306), .B2(DRAM_DATA_IN[27]), .A(n4305), .ZN(n4301) );
  INV_X1 U5444 ( .A(n4301), .ZN(\DP/RegLMD/N30 ) );
  AOI21_X1 U5445 ( .B1(n4306), .B2(DRAM_DATA_IN[28]), .A(n4305), .ZN(n4302) );
  INV_X1 U5446 ( .A(n4302), .ZN(\DP/RegLMD/N31 ) );
  AOI21_X1 U5447 ( .B1(n4306), .B2(DRAM_DATA_IN[29]), .A(n4305), .ZN(n4303) );
  INV_X1 U5448 ( .A(n4303), .ZN(\DP/RegLMD/N32 ) );
  AOI21_X1 U5449 ( .B1(n4306), .B2(DRAM_DATA_IN[30]), .A(n4305), .ZN(n4304) );
  INV_X1 U5450 ( .A(n4304), .ZN(\DP/RegLMD/N33 ) );
  AOI21_X1 U5451 ( .B1(n4306), .B2(DRAM_DATA_IN[31]), .A(n4305), .ZN(n4307) );
  INV_X1 U5452 ( .A(n4307), .ZN(\DP/RegLMD/N34 ) );
  AND2_X1 U5453 ( .A1(\DP/LOAD8[1] ), .A2(n4308), .ZN(\DP/RegLMD/N4 ) );
  AND2_X1 U5454 ( .A1(\DP/LOAD8[2] ), .A2(n4308), .ZN(\DP/RegLMD/N5 ) );
  AND2_X1 U5455 ( .A1(\DP/LOAD8[3] ), .A2(n4308), .ZN(\DP/RegLMD/N6 ) );
  AND2_X1 U5456 ( .A1(\DP/LOAD8[4] ), .A2(n4308), .ZN(\DP/RegLMD/N7 ) );
  AND2_X1 U5457 ( .A1(\DP/LOAD8[5] ), .A2(n4308), .ZN(\DP/RegLMD/N8 ) );
  AND2_X1 U5458 ( .A1(\DP/LOAD8[6] ), .A2(n4308), .ZN(\DP/RegLMD/N9 ) );
  AND2_X1 U5459 ( .A1(RST), .A2(\DP/RegB_out[7] ), .ZN(\DP/RegME/N10 ) );
  AND2_X1 U5460 ( .A1(RST), .A2(\DP/RegB_out[8] ), .ZN(\DP/RegME/N11 ) );
  AND2_X1 U5461 ( .A1(RST), .A2(\DP/RegB_out[9] ), .ZN(\DP/RegME/N12 ) );
  AND2_X1 U5462 ( .A1(RST), .A2(\DP/RegB_out[10] ), .ZN(\DP/RegME/N13 ) );
  AND2_X1 U5463 ( .A1(RST), .A2(\DP/RegB_out[11] ), .ZN(\DP/RegME/N14 ) );
  AND2_X1 U5464 ( .A1(RST), .A2(\DP/RegB_out[12] ), .ZN(\DP/RegME/N15 ) );
  AND2_X1 U5465 ( .A1(RST), .A2(\DP/RegB_out[13] ), .ZN(\DP/RegME/N16 ) );
  AND2_X1 U5466 ( .A1(RST), .A2(\DP/RegB_out[14] ), .ZN(\DP/RegME/N17 ) );
  AND2_X1 U5467 ( .A1(RST), .A2(\DP/RegB_out[15] ), .ZN(\DP/RegME/N18 ) );
  AND2_X1 U5468 ( .A1(RST), .A2(\DP/RegB_out[16] ), .ZN(\DP/RegME/N19 ) );
  AND2_X1 U5469 ( .A1(RST), .A2(\DP/RegB_out[17] ), .ZN(\DP/RegME/N20 ) );
  AND2_X1 U5470 ( .A1(RST), .A2(\DP/RegB_out[18] ), .ZN(\DP/RegME/N21 ) );
  AND2_X1 U5471 ( .A1(RST), .A2(\DP/RegB_out[19] ), .ZN(\DP/RegME/N22 ) );
  AND2_X1 U5472 ( .A1(RST), .A2(\DP/RegB_out[20] ), .ZN(\DP/RegME/N23 ) );
  AND2_X1 U5473 ( .A1(RST), .A2(\DP/RegB_out[21] ), .ZN(\DP/RegME/N24 ) );
  AND2_X1 U5474 ( .A1(RST), .A2(\DP/RegB_out[22] ), .ZN(\DP/RegME/N25 ) );
  AND2_X1 U5475 ( .A1(RST), .A2(\DP/RegB_out[23] ), .ZN(\DP/RegME/N26 ) );
  AND2_X1 U5476 ( .A1(RST), .A2(\DP/RegB_out[24] ), .ZN(\DP/RegME/N27 ) );
  AND2_X1 U5477 ( .A1(RST), .A2(\DP/RegB_out[25] ), .ZN(\DP/RegME/N28 ) );
  AND2_X1 U5478 ( .A1(RST), .A2(\DP/RegB_out[26] ), .ZN(\DP/RegME/N29 ) );
  AND2_X1 U5479 ( .A1(RST), .A2(\DP/RegB_out[0] ), .ZN(\DP/RegME/N3 ) );
  AND2_X1 U5480 ( .A1(RST), .A2(\DP/RegB_out[27] ), .ZN(\DP/RegME/N30 ) );
  AND2_X1 U5481 ( .A1(RST), .A2(\DP/RegB_out[28] ), .ZN(\DP/RegME/N31 ) );
  AND2_X1 U5482 ( .A1(RST), .A2(\DP/RegB_out[29] ), .ZN(\DP/RegME/N32 ) );
  AND2_X1 U5483 ( .A1(RST), .A2(\DP/RegB_out[30] ), .ZN(\DP/RegME/N33 ) );
  AND2_X1 U5484 ( .A1(RST), .A2(\DP/RegB_out[31] ), .ZN(\DP/RegME/N34 ) );
  AND2_X1 U5485 ( .A1(RST), .A2(\DP/RegB_out[1] ), .ZN(\DP/RegME/N4 ) );
  AND2_X1 U5486 ( .A1(RST), .A2(\DP/RegB_out[2] ), .ZN(\DP/RegME/N5 ) );
  AND2_X1 U5487 ( .A1(RST), .A2(\DP/RegB_out[3] ), .ZN(\DP/RegME/N6 ) );
  AND2_X1 U5488 ( .A1(RST), .A2(\DP/RegB_out[4] ), .ZN(\DP/RegME/N7 ) );
  AND2_X1 U5489 ( .A1(RST), .A2(\DP/RegB_out[5] ), .ZN(\DP/RegME/N8 ) );
  AND2_X1 U5490 ( .A1(RST), .A2(\DP/RegB_out[6] ), .ZN(\DP/RegME/N9 ) );
  NAND3_X1 U5491 ( .A1(IROM_ADDR[0]), .A2(IROM_ADDR[1]), .A3(IROM_ADDR[2]), 
        .ZN(n4399) );
  OAI21_X1 U5497 ( .B1(n4309), .B2(IROM_ADDR[7]), .A(n2437), .ZN(n4311) );
  AOI22_X1 U5498 ( .A1(n2436), .A2(\DP/RegALU2/N10 ), .B1(n2435), .B2(
        \DP/RegA1_out[7] ), .ZN(n4310) );
  OAI21_X1 U5499 ( .B1(n4312), .B2(n4311), .A(n4310), .ZN(\PC/N10 ) );
  AOI22_X1 U5500 ( .A1(n4414), .A2(\DP/RegALU2/N11 ), .B1(n4413), .B2(
        \DP/RegA1_out[8] ), .ZN(n4314) );
  OAI211_X1 U5502 ( .C1(n4312), .C2(IROM_ADDR[8]), .A(n2438), .B(n4315), .ZN(
        n4313) );
  NAND2_X1 U5503 ( .A1(n4314), .A2(n4313), .ZN(\PC/N11 ) );
  OAI21_X1 U5505 ( .B1(n4316), .B2(IROM_ADDR[9]), .A(n2437), .ZN(n4318) );
  AOI22_X1 U5506 ( .A1(n2436), .A2(\DP/RegALU2/N12 ), .B1(n2435), .B2(
        \DP/RegA1_out[9] ), .ZN(n4317) );
  OAI21_X1 U5507 ( .B1(n4319), .B2(n4318), .A(n4317), .ZN(\PC/N12 ) );
  AOI22_X1 U5508 ( .A1(n4414), .A2(\DP/RegALU2/N13 ), .B1(n4413), .B2(
        \DP/RegA1_out[10] ), .ZN(n4321) );
  OAI211_X1 U5510 ( .C1(n4319), .C2(IROM_ADDR[10]), .A(n2438), .B(n4322), .ZN(
        n4320) );
  NAND2_X1 U5511 ( .A1(n4321), .A2(n4320), .ZN(\PC/N13 ) );
  OAI21_X1 U5513 ( .B1(n4323), .B2(IROM_ADDR[11]), .A(n2437), .ZN(n4325) );
  AOI22_X1 U5514 ( .A1(n2436), .A2(\DP/RegALU2/N14 ), .B1(n2435), .B2(
        \DP/RegA1_out[11] ), .ZN(n4324) );
  OAI21_X1 U5515 ( .B1(n4326), .B2(n4325), .A(n4324), .ZN(\PC/N14 ) );
  AOI22_X1 U5516 ( .A1(n4414), .A2(\DP/RegALU2/N15 ), .B1(n4413), .B2(
        \DP/RegA1_out[12] ), .ZN(n4328) );
  OAI211_X1 U5518 ( .C1(n4326), .C2(w_PC_OUT[12]), .A(n2437), .B(n4329), .ZN(
        n4327) );
  NAND2_X1 U5519 ( .A1(n4328), .A2(n4327), .ZN(\PC/N15 ) );
  OAI21_X1 U5521 ( .B1(n4330), .B2(w_PC_OUT[13]), .A(n2438), .ZN(n4332) );
  AOI22_X1 U5522 ( .A1(n4414), .A2(\DP/RegALU2/N16 ), .B1(n4413), .B2(
        \DP/RegA1_out[13] ), .ZN(n4331) );
  OAI21_X1 U5523 ( .B1(n4333), .B2(n4332), .A(n4331), .ZN(\PC/N16 ) );
  AOI22_X1 U5524 ( .A1(n4414), .A2(\DP/RegALU2/N17 ), .B1(n4413), .B2(
        \DP/RegA1_out[14] ), .ZN(n4335) );
  OAI211_X1 U5526 ( .C1(n4333), .C2(w_PC_OUT[14]), .A(n2437), .B(n4336), .ZN(
        n4334) );
  NAND2_X1 U5527 ( .A1(n4335), .A2(n4334), .ZN(\PC/N17 ) );
  OAI21_X1 U5529 ( .B1(n4337), .B2(w_PC_OUT[15]), .A(n2438), .ZN(n4339) );
  AOI22_X1 U5530 ( .A1(n4414), .A2(\DP/RegALU2/N18 ), .B1(n4413), .B2(
        \DP/RegA1_out[15] ), .ZN(n4338) );
  OAI21_X1 U5531 ( .B1(n4340), .B2(n4339), .A(n4338), .ZN(\PC/N18 ) );
  AOI22_X1 U5532 ( .A1(n4414), .A2(\DP/RegALU2/N19 ), .B1(n4413), .B2(
        \DP/RegA1_out[16] ), .ZN(n4342) );
  OAI211_X1 U5534 ( .C1(n4340), .C2(w_PC_OUT[16]), .A(n2437), .B(n4343), .ZN(
        n4341) );
  NAND2_X1 U5535 ( .A1(n4342), .A2(n4341), .ZN(\PC/N19 ) );
  OR2_X1 U5536 ( .A1(w_IF_EN), .A2(n2461), .ZN(\PC/N2 ) );
  OAI21_X1 U5538 ( .B1(n4344), .B2(w_PC_OUT[17]), .A(n2438), .ZN(n4346) );
  AOI22_X1 U5539 ( .A1(n4414), .A2(\DP/RegALU2/N20 ), .B1(n4413), .B2(
        \DP/RegA1_out[17] ), .ZN(n4345) );
  OAI21_X1 U5540 ( .B1(n4347), .B2(n4346), .A(n4345), .ZN(\PC/N20 ) );
  AOI22_X1 U5541 ( .A1(n4414), .A2(\DP/RegALU2/N21 ), .B1(n4413), .B2(
        \DP/RegA1_out[18] ), .ZN(n4349) );
  OAI211_X1 U5543 ( .C1(n4347), .C2(w_PC_OUT[18]), .A(n2437), .B(n4531), .ZN(
        n4348) );
  NAND2_X1 U5544 ( .A1(n4349), .A2(n4348), .ZN(\PC/N21 ) );
  OAI21_X1 U5546 ( .B1(n4351), .B2(w_PC_OUT[19]), .A(n2438), .ZN(n4353) );
  AOI22_X1 U5547 ( .A1(n2436), .A2(\DP/RegALU2/N22 ), .B1(n4413), .B2(
        \DP/RegA1_out[19] ), .ZN(n4352) );
  AOI22_X1 U5549 ( .A1(n2436), .A2(\DP/RegALU2/N23 ), .B1(n2435), .B2(
        \DP/RegA1_out[20] ), .ZN(n4356) );
  NAND2_X1 U5552 ( .A1(n4356), .A2(n4355), .ZN(\PC/N23 ) );
  OAI21_X1 U5554 ( .B1(n4358), .B2(w_PC_OUT[21]), .A(n2438), .ZN(n4360) );
  AOI22_X1 U5555 ( .A1(n2436), .A2(\DP/RegALU2/N24 ), .B1(n4413), .B2(
        \DP/RegA1_out[21] ), .ZN(n4359) );
  OAI21_X1 U5556 ( .B1(n4361), .B2(n4360), .A(n4359), .ZN(\PC/N24 ) );
  AOI22_X1 U5557 ( .A1(n2436), .A2(\DP/RegALU2/N25 ), .B1(n2435), .B2(
        \DP/RegA1_out[22] ), .ZN(n4363) );
  OAI211_X1 U5559 ( .C1(n4361), .C2(w_PC_OUT[22]), .A(n2437), .B(n4364), .ZN(
        n4362) );
  NAND2_X1 U5560 ( .A1(n4363), .A2(n4362), .ZN(\PC/N25 ) );
  OAI21_X1 U5562 ( .B1(n4365), .B2(w_PC_OUT[23]), .A(n2438), .ZN(n4367) );
  AOI22_X1 U5563 ( .A1(n2436), .A2(\DP/RegALU2/N26 ), .B1(n4413), .B2(
        \DP/RegA1_out[23] ), .ZN(n4366) );
  OAI21_X1 U5564 ( .B1(n4368), .B2(n4367), .A(n4366), .ZN(\PC/N26 ) );
  AOI22_X1 U5565 ( .A1(n2436), .A2(\DP/RegALU2/N27 ), .B1(n2435), .B2(
        \DP/RegA1_out[24] ), .ZN(n4370) );
  OAI211_X1 U5567 ( .C1(n4368), .C2(w_PC_OUT[24]), .A(n2437), .B(n4371), .ZN(
        n4369) );
  NAND2_X1 U5568 ( .A1(n4370), .A2(n4369), .ZN(\PC/N27 ) );
  AOI22_X1 U5571 ( .A1(n2436), .A2(\DP/RegALU2/N28 ), .B1(n4413), .B2(
        \DP/RegA1_out[25] ), .ZN(n4373) );
  AOI22_X1 U5573 ( .A1(n2436), .A2(\DP/RegALU2/N29 ), .B1(n2435), .B2(
        \DP/RegA1_out[26] ), .ZN(n4377) );
  NAND2_X1 U5576 ( .A1(n4377), .A2(n4376), .ZN(\PC/N29 ) );
  AOI22_X1 U5577 ( .A1(n2436), .A2(\DP/RegALU2/N3 ), .B1(n4413), .B2(
        \DP/RegA1_out[0] ), .ZN(n4378) );
  OAI21_X1 U5578 ( .B1(IROM_ADDR[0]), .B2(n2381), .A(n4378), .ZN(\PC/N3 ) );
  OAI21_X1 U5580 ( .B1(n4380), .B2(w_PC_OUT[27]), .A(n2438), .ZN(n4382) );
  AOI22_X1 U5581 ( .A1(n2436), .A2(\DP/RegALU2/N30 ), .B1(n2435), .B2(
        \DP/RegA1_out[27] ), .ZN(n4381) );
  OAI21_X1 U5582 ( .B1(n4383), .B2(n4382), .A(n4381), .ZN(\PC/N30 ) );
  AOI22_X1 U5583 ( .A1(n4414), .A2(\DP/RegALU2/N31 ), .B1(n4413), .B2(
        \DP/RegA1_out[28] ), .ZN(n4385) );
  NAND2_X1 U5586 ( .A1(n4385), .A2(n4384), .ZN(\PC/N31 ) );
  OAI21_X1 U5588 ( .B1(n4387), .B2(w_PC_OUT[29]), .A(n2438), .ZN(n4389) );
  AOI22_X1 U5589 ( .A1(n4414), .A2(\DP/RegALU2/N32 ), .B1(n4413), .B2(
        \DP/RegA1_out[29] ), .ZN(n4388) );
  OAI21_X1 U5590 ( .B1(n4390), .B2(n4389), .A(n4388), .ZN(\PC/N32 ) );
  AOI22_X1 U5593 ( .A1(n2436), .A2(\DP/RegALU2/N33 ), .B1(n2435), .B2(
        \DP/RegA1_out[30] ), .ZN(n4391) );
  OAI21_X1 U5594 ( .B1(n2381), .B2(n4392), .A(n4391), .ZN(\PC/N33 ) );
  XOR2_X1 U5595 ( .A(n4393), .B(w_PC_OUT[31]), .Z(n4395) );
  AOI22_X1 U5596 ( .A1(n2436), .A2(\DP/RegALU2/N34 ), .B1(n2435), .B2(
        \DP/RegA1_out[31] ), .ZN(n4394) );
  OAI21_X1 U5597 ( .B1(n4395), .B2(n2381), .A(n4394), .ZN(\PC/N34 ) );
  AOI22_X1 U5598 ( .A1(n2436), .A2(\DP/RegALU2/N4 ), .B1(n2435), .B2(
        \DP/RegA1_out[1] ), .ZN(n4397) );
  NAND2_X1 U5599 ( .A1(IROM_ADDR[0]), .A2(IROM_ADDR[1]), .ZN(n4398) );
  OAI211_X1 U5600 ( .C1(IROM_ADDR[0]), .C2(IROM_ADDR[1]), .A(n2438), .B(n4398), 
        .ZN(n4396) );
  NAND2_X1 U5601 ( .A1(n4397), .A2(n4396), .ZN(\PC/N4 ) );
  AOI22_X1 U5602 ( .A1(n2436), .A2(\DP/RegALU2/N5 ), .B1(n2435), .B2(
        \DP/RegA1_out[2] ), .ZN(n4402) );
  INV_X1 U5603 ( .A(n4398), .ZN(n4400) );
  OAI211_X1 U5604 ( .C1(n4400), .C2(IROM_ADDR[2]), .A(n2438), .B(n4560), .ZN(
        n4401) );
  NAND2_X1 U5605 ( .A1(n4402), .A2(n4401), .ZN(\PC/N5 ) );
  OAI21_X1 U5606 ( .B1(n4403), .B2(IROM_ADDR[3]), .A(n2437), .ZN(n4405) );
  AOI22_X1 U5607 ( .A1(n2436), .A2(\DP/RegALU2/N6 ), .B1(n2435), .B2(
        \DP/RegA1_out[3] ), .ZN(n4404) );
  OAI21_X1 U5608 ( .B1(n4407), .B2(n4405), .A(n4404), .ZN(\PC/N6 ) );
  AOI22_X1 U5609 ( .A1(n2436), .A2(\DP/RegALU2/N7 ), .B1(n2435), .B2(
        \DP/RegA1_out[4] ), .ZN(n4409) );
  OAI211_X1 U5610 ( .C1(n4407), .C2(IROM_ADDR[4]), .A(n2438), .B(n4406), .ZN(
        n4408) );
  NAND2_X1 U5611 ( .A1(n4409), .A2(n4408), .ZN(\PC/N7 ) );
  OAI21_X1 U5612 ( .B1(n4410), .B2(IROM_ADDR[5]), .A(n2438), .ZN(n4412) );
  AOI22_X1 U5613 ( .A1(n2436), .A2(\DP/RegALU2/N8 ), .B1(n2435), .B2(
        \DP/RegA1_out[5] ), .ZN(n4411) );
  OAI21_X1 U5614 ( .B1(n4416), .B2(n4412), .A(n4411), .ZN(\PC/N8 ) );
  AOI22_X1 U5615 ( .A1(n2436), .A2(\DP/RegALU2/N9 ), .B1(n2435), .B2(
        \DP/RegA1_out[6] ), .ZN(n4418) );
  OAI211_X1 U5616 ( .C1(n4416), .C2(IROM_ADDR[6]), .A(n2437), .B(n4415), .ZN(
        n4417) );
  NAND2_X1 U5617 ( .A1(n4418), .A2(n4417), .ZN(\PC/N9 ) );
  AND2_X1 U5618 ( .A1(RST), .A2(\DP/NPC1[7] ), .ZN(\DP/RegNPC1/N10 ) );
  AND2_X1 U5619 ( .A1(RST), .A2(\DP/NPC1[8] ), .ZN(\DP/RegNPC1/N11 ) );
  AND2_X1 U5620 ( .A1(RST), .A2(\DP/NPC1[9] ), .ZN(\DP/RegNPC1/N12 ) );
  AND2_X1 U5621 ( .A1(RST), .A2(\DP/NPC1[10] ), .ZN(\DP/RegNPC1/N13 ) );
  AND2_X1 U5622 ( .A1(RST), .A2(\DP/NPC1[11] ), .ZN(\DP/RegNPC1/N14 ) );
  AND2_X1 U5623 ( .A1(RST), .A2(\DP/NPC1[12] ), .ZN(\DP/RegNPC1/N15 ) );
  AND2_X1 U5624 ( .A1(RST), .A2(\DP/NPC1[13] ), .ZN(\DP/RegNPC1/N16 ) );
  AND2_X1 U5625 ( .A1(RST), .A2(\DP/NPC1[14] ), .ZN(\DP/RegNPC1/N17 ) );
  AND2_X1 U5626 ( .A1(RST), .A2(\DP/NPC1[15] ), .ZN(\DP/RegNPC1/N18 ) );
  AND2_X1 U5627 ( .A1(RST), .A2(\DP/NPC1[16] ), .ZN(\DP/RegNPC1/N19 ) );
  AND2_X1 U5628 ( .A1(RST), .A2(\DP/NPC1[17] ), .ZN(\DP/RegNPC1/N20 ) );
  AND2_X1 U5629 ( .A1(RST), .A2(\DP/NPC1[18] ), .ZN(\DP/RegNPC1/N21 ) );
  AND2_X1 U5630 ( .A1(RST), .A2(\DP/NPC1[19] ), .ZN(\DP/RegNPC1/N22 ) );
  AND2_X1 U5631 ( .A1(RST), .A2(\DP/NPC1[20] ), .ZN(\DP/RegNPC1/N23 ) );
  AND2_X1 U5632 ( .A1(RST), .A2(\DP/NPC1[21] ), .ZN(\DP/RegNPC1/N24 ) );
  AND2_X1 U5633 ( .A1(RST), .A2(\DP/NPC1[22] ), .ZN(\DP/RegNPC1/N25 ) );
  AND2_X1 U5634 ( .A1(RST), .A2(\DP/NPC1[23] ), .ZN(\DP/RegNPC1/N26 ) );
  AND2_X1 U5635 ( .A1(RST), .A2(\DP/NPC1[24] ), .ZN(\DP/RegNPC1/N27 ) );
  AND2_X1 U5636 ( .A1(RST), .A2(\DP/NPC1[25] ), .ZN(\DP/RegNPC1/N28 ) );
  AND2_X1 U5637 ( .A1(RST), .A2(\DP/NPC1[26] ), .ZN(\DP/RegNPC1/N29 ) );
  AND2_X1 U5638 ( .A1(RST), .A2(\DP/NPC1[0] ), .ZN(\DP/RegNPC1/N3 ) );
  AND2_X1 U5639 ( .A1(RST), .A2(\DP/NPC1[27] ), .ZN(\DP/RegNPC1/N30 ) );
  AND2_X1 U5640 ( .A1(RST), .A2(\DP/NPC1[28] ), .ZN(\DP/RegNPC1/N31 ) );
  AND2_X1 U5641 ( .A1(RST), .A2(\DP/NPC1[29] ), .ZN(\DP/RegNPC1/N32 ) );
  AND2_X1 U5642 ( .A1(RST), .A2(\DP/NPC1[30] ), .ZN(\DP/RegNPC1/N33 ) );
  AND2_X1 U5643 ( .A1(RST), .A2(\DP/NPC1[31] ), .ZN(\DP/RegNPC1/N34 ) );
  AND2_X1 U5644 ( .A1(RST), .A2(\DP/NPC1[1] ), .ZN(\DP/RegNPC1/N4 ) );
  AND2_X1 U5645 ( .A1(RST), .A2(\DP/NPC1[2] ), .ZN(\DP/RegNPC1/N5 ) );
  AND2_X1 U5646 ( .A1(RST), .A2(\DP/NPC1[3] ), .ZN(\DP/RegNPC1/N6 ) );
  AND2_X1 U5647 ( .A1(RST), .A2(\DP/NPC1[4] ), .ZN(\DP/RegNPC1/N7 ) );
  AND2_X1 U5648 ( .A1(RST), .A2(\DP/NPC1[5] ), .ZN(\DP/RegNPC1/N8 ) );
  AND2_X1 U5649 ( .A1(RST), .A2(\DP/NPC1[6] ), .ZN(\DP/RegNPC1/N9 ) );
  AND2_X1 U5650 ( .A1(RST), .A2(\DP/NPC2[7] ), .ZN(\DP/RegNPC2/N10 ) );
  AND2_X1 U5651 ( .A1(RST), .A2(\DP/NPC2[8] ), .ZN(\DP/RegNPC2/N11 ) );
  AND2_X1 U5652 ( .A1(RST), .A2(\DP/NPC2[9] ), .ZN(\DP/RegNPC2/N12 ) );
  AND2_X1 U5653 ( .A1(RST), .A2(\DP/NPC2[10] ), .ZN(\DP/RegNPC2/N13 ) );
  AND2_X1 U5654 ( .A1(RST), .A2(\DP/NPC2[11] ), .ZN(\DP/RegNPC2/N14 ) );
  AND2_X1 U5655 ( .A1(RST), .A2(\DP/NPC2[12] ), .ZN(\DP/RegNPC2/N15 ) );
  AND2_X1 U5656 ( .A1(RST), .A2(\DP/NPC2[13] ), .ZN(\DP/RegNPC2/N16 ) );
  AND2_X1 U5657 ( .A1(RST), .A2(\DP/NPC2[14] ), .ZN(\DP/RegNPC2/N17 ) );
  AND2_X1 U5658 ( .A1(RST), .A2(\DP/NPC2[15] ), .ZN(\DP/RegNPC2/N18 ) );
  AND2_X1 U5659 ( .A1(RST), .A2(\DP/NPC2[16] ), .ZN(\DP/RegNPC2/N19 ) );
  AND2_X1 U5660 ( .A1(RST), .A2(\DP/NPC2[17] ), .ZN(\DP/RegNPC2/N20 ) );
  AND2_X1 U5661 ( .A1(RST), .A2(\DP/NPC2[18] ), .ZN(\DP/RegNPC2/N21 ) );
  AND2_X1 U5662 ( .A1(RST), .A2(\DP/NPC2[19] ), .ZN(\DP/RegNPC2/N22 ) );
  AND2_X1 U5663 ( .A1(RST), .A2(\DP/NPC2[20] ), .ZN(\DP/RegNPC2/N23 ) );
  AND2_X1 U5664 ( .A1(RST), .A2(\DP/NPC2[21] ), .ZN(\DP/RegNPC2/N24 ) );
  AND2_X1 U5665 ( .A1(RST), .A2(\DP/NPC2[22] ), .ZN(\DP/RegNPC2/N25 ) );
  AND2_X1 U5666 ( .A1(RST), .A2(\DP/NPC2[23] ), .ZN(\DP/RegNPC2/N26 ) );
  AND2_X1 U5667 ( .A1(RST), .A2(\DP/NPC2[24] ), .ZN(\DP/RegNPC2/N27 ) );
  AND2_X1 U5668 ( .A1(RST), .A2(\DP/NPC2[25] ), .ZN(\DP/RegNPC2/N28 ) );
  AND2_X1 U5669 ( .A1(RST), .A2(\DP/NPC2[26] ), .ZN(\DP/RegNPC2/N29 ) );
  AND2_X1 U5670 ( .A1(RST), .A2(\DP/NPC2[0] ), .ZN(\DP/RegNPC2/N3 ) );
  AND2_X1 U5671 ( .A1(RST), .A2(\DP/NPC2[27] ), .ZN(\DP/RegNPC2/N30 ) );
  AND2_X1 U5672 ( .A1(RST), .A2(\DP/NPC2[28] ), .ZN(\DP/RegNPC2/N31 ) );
  AND2_X1 U5673 ( .A1(RST), .A2(\DP/NPC2[29] ), .ZN(\DP/RegNPC2/N32 ) );
  AND2_X1 U5674 ( .A1(RST), .A2(\DP/NPC2[30] ), .ZN(\DP/RegNPC2/N33 ) );
  AND2_X1 U5675 ( .A1(\DP/NPC2[31] ), .A2(RST), .ZN(\DP/RegNPC2/N34 ) );
  AND2_X1 U5676 ( .A1(RST), .A2(\DP/NPC2[1] ), .ZN(\DP/RegNPC2/N4 ) );
  AND2_X1 U5677 ( .A1(RST), .A2(\DP/NPC2[2] ), .ZN(\DP/RegNPC2/N5 ) );
  AND2_X1 U5678 ( .A1(RST), .A2(\DP/NPC2[3] ), .ZN(\DP/RegNPC2/N6 ) );
  AND2_X1 U5679 ( .A1(RST), .A2(\DP/NPC2[4] ), .ZN(\DP/RegNPC2/N7 ) );
  AND2_X1 U5680 ( .A1(RST), .A2(\DP/NPC2[5] ), .ZN(\DP/RegNPC2/N8 ) );
  AND2_X1 U5681 ( .A1(RST), .A2(\DP/NPC2[6] ), .ZN(\DP/RegNPC2/N9 ) );
  AND2_X1 U5682 ( .A1(RST), .A2(\DP/NPC3[7] ), .ZN(\DP/RegNPC3/N10 ) );
  AND2_X1 U5683 ( .A1(RST), .A2(\DP/NPC3[8] ), .ZN(\DP/RegNPC3/N11 ) );
  AND2_X1 U5684 ( .A1(RST), .A2(\DP/NPC3[9] ), .ZN(\DP/RegNPC3/N12 ) );
  AND2_X1 U5685 ( .A1(RST), .A2(\DP/NPC3[10] ), .ZN(\DP/RegNPC3/N13 ) );
  AND2_X1 U5686 ( .A1(RST), .A2(\DP/NPC3[11] ), .ZN(\DP/RegNPC3/N14 ) );
  AND2_X1 U5687 ( .A1(RST), .A2(\DP/NPC3[12] ), .ZN(\DP/RegNPC3/N15 ) );
  AND2_X1 U5688 ( .A1(RST), .A2(\DP/NPC3[13] ), .ZN(\DP/RegNPC3/N16 ) );
  AND2_X1 U5689 ( .A1(RST), .A2(\DP/NPC3[14] ), .ZN(\DP/RegNPC3/N17 ) );
  AND2_X1 U5690 ( .A1(RST), .A2(\DP/NPC3[15] ), .ZN(\DP/RegNPC3/N18 ) );
  AND2_X1 U5691 ( .A1(RST), .A2(\DP/NPC3[16] ), .ZN(\DP/RegNPC3/N19 ) );
  OR2_X1 U5692 ( .A1(\DP/JL1 ), .A2(n2461), .ZN(\DP/RegNPC3/N2 ) );
  AND2_X1 U5693 ( .A1(RST), .A2(\DP/NPC3[17] ), .ZN(\DP/RegNPC3/N20 ) );
  AND2_X1 U5694 ( .A1(RST), .A2(\DP/NPC3[18] ), .ZN(\DP/RegNPC3/N21 ) );
  AND2_X1 U5695 ( .A1(RST), .A2(\DP/NPC3[19] ), .ZN(\DP/RegNPC3/N22 ) );
  AND2_X1 U5696 ( .A1(RST), .A2(\DP/NPC3[20] ), .ZN(\DP/RegNPC3/N23 ) );
  AND2_X1 U5697 ( .A1(RST), .A2(\DP/NPC3[21] ), .ZN(\DP/RegNPC3/N24 ) );
  AND2_X1 U5698 ( .A1(RST), .A2(\DP/NPC3[22] ), .ZN(\DP/RegNPC3/N25 ) );
  AND2_X1 U5699 ( .A1(RST), .A2(\DP/NPC3[23] ), .ZN(\DP/RegNPC3/N26 ) );
  AND2_X1 U5700 ( .A1(RST), .A2(\DP/NPC3[24] ), .ZN(\DP/RegNPC3/N27 ) );
  AND2_X1 U5701 ( .A1(RST), .A2(\DP/NPC3[25] ), .ZN(\DP/RegNPC3/N28 ) );
  AND2_X1 U5702 ( .A1(RST), .A2(\DP/NPC3[26] ), .ZN(\DP/RegNPC3/N29 ) );
  AND2_X1 U5703 ( .A1(RST), .A2(\DP/NPC3[0] ), .ZN(\DP/RegNPC3/N3 ) );
  AND2_X1 U5704 ( .A1(RST), .A2(\DP/NPC3[27] ), .ZN(\DP/RegNPC3/N30 ) );
  AND2_X1 U5705 ( .A1(RST), .A2(\DP/NPC3[28] ), .ZN(\DP/RegNPC3/N31 ) );
  AND2_X1 U5706 ( .A1(RST), .A2(\DP/NPC3[29] ), .ZN(\DP/RegNPC3/N32 ) );
  AND2_X1 U5707 ( .A1(RST), .A2(\DP/NPC3[30] ), .ZN(\DP/RegNPC3/N33 ) );
  AND2_X1 U5708 ( .A1(RST), .A2(\DP/NPC3[31] ), .ZN(\DP/RegNPC3/N34 ) );
  AND2_X1 U5709 ( .A1(RST), .A2(\DP/NPC3[1] ), .ZN(\DP/RegNPC3/N4 ) );
  AND2_X1 U5710 ( .A1(RST), .A2(\DP/NPC3[2] ), .ZN(\DP/RegNPC3/N5 ) );
  AND2_X1 U5711 ( .A1(RST), .A2(\DP/NPC3[3] ), .ZN(\DP/RegNPC3/N6 ) );
  AND2_X1 U5712 ( .A1(RST), .A2(\DP/NPC3[4] ), .ZN(\DP/RegNPC3/N7 ) );
  AND2_X1 U5713 ( .A1(RST), .A2(\DP/NPC3[5] ), .ZN(\DP/RegNPC3/N8 ) );
  AND2_X1 U5714 ( .A1(RST), .A2(\DP/NPC3[6] ), .ZN(\DP/RegNPC3/N9 ) );
  AND2_X1 U5721 ( .A1(RST), .A2(\DP/RD1[0] ), .ZN(\DP/RegRD2/N3 ) );
  NOR2_X1 U5722 ( .A1(n2460), .A2(n2378), .ZN(\DP/RegRD2/N4 ) );
  NOR2_X1 U5723 ( .A1(n2460), .A2(n2380), .ZN(\DP/RegRD2/N5 ) );
  NOR2_X1 U5724 ( .A1(n2460), .A2(n4635), .ZN(\DP/RegRD2/N6 ) );
  AND2_X1 U5725 ( .A1(RST), .A2(\DP/RD1[4] ), .ZN(\DP/RegRD2/N7 ) );
  AND2_X1 U5726 ( .A1(RST), .A2(\DP/RD2[0] ), .ZN(\DP/RegRD3/N3 ) );
  AND2_X1 U5727 ( .A1(RST), .A2(\DP/RD2[1] ), .ZN(\DP/RegRD3/N4 ) );
  NOR2_X1 U5728 ( .A1(n2460), .A2(n2367), .ZN(\DP/RegRD3/N5 ) );
  NOR2_X1 U5729 ( .A1(n400), .A2(n2460), .ZN(\DP/RegRD3/N6 ) );
  NOR2_X1 U5730 ( .A1(n401), .A2(n2460), .ZN(\DP/RegRD3/N7 ) );
  OAI21_X1 U5731 ( .B1(n204), .B2(n205), .A(n206), .ZN(n4426) );
  AOI21_X1 U5732 ( .B1(n204), .B2(n205), .A(n4426), .ZN(n4427) );
  INV_X1 U5733 ( .A(n4427), .ZN(n4489) );
  AOI22_X1 U5734 ( .A1(\DP/FwdD ), .A2(n4428), .B1(\DP/RegME_out[7] ), .B2(
        n2402), .ZN(n4478) );
  NAND3_X1 U5735 ( .A1(n205), .A2(n204), .A3(n2403), .ZN(n4490) );
  NOR2_X1 U5736 ( .A1(n4478), .A2(n4490), .ZN(n4481) );
  AOI21_X1 U5737 ( .B1(n4482), .B2(\DP/RegME_out[10] ), .A(n4481), .ZN(n4429)
         );
  OAI21_X1 U5738 ( .B1(n4430), .B2(n4484), .A(n4429), .ZN(DRAM_DATA_OUT[10])
         );
  AOI21_X1 U5739 ( .B1(n4482), .B2(\DP/RegME_out[11] ), .A(n4481), .ZN(n4431)
         );
  OAI21_X1 U5740 ( .B1(n4565), .B2(n4484), .A(n4431), .ZN(DRAM_DATA_OUT[11])
         );
  AOI21_X1 U5741 ( .B1(n4482), .B2(\DP/RegME_out[12] ), .A(n4481), .ZN(n4433)
         );
  AOI21_X1 U5743 ( .B1(n4482), .B2(\DP/RegME_out[13] ), .A(n4481), .ZN(n4435)
         );
  OAI21_X1 U5744 ( .B1(n4556), .B2(n4484), .A(n4435), .ZN(DRAM_DATA_OUT[13])
         );
  AOI21_X1 U5745 ( .B1(n4482), .B2(\DP/RegME_out[14] ), .A(n4481), .ZN(n4437)
         );
  OAI21_X1 U5746 ( .B1(n4542), .B2(n4484), .A(n4437), .ZN(DRAM_DATA_OUT[14])
         );
  AOI21_X1 U5747 ( .B1(n4482), .B2(\DP/RegME_out[15] ), .A(n4481), .ZN(n4439)
         );
  OAI21_X1 U5748 ( .B1(n4440), .B2(n4484), .A(n4439), .ZN(DRAM_DATA_OUT[15])
         );
  NAND2_X1 U5749 ( .A1(n4472), .A2(\DP/RegME_out[16] ), .ZN(n4441) );
  OAI211_X1 U5750 ( .C1(n4442), .C2(n4475), .A(n4441), .B(n4473), .ZN(
        DRAM_DATA_OUT[16]) );
  NAND2_X1 U5751 ( .A1(n4472), .A2(\DP/RegME_out[17] ), .ZN(n4443) );
  OAI211_X1 U5752 ( .C1(n4444), .C2(n4475), .A(n4443), .B(n4473), .ZN(
        DRAM_DATA_OUT[17]) );
  NAND2_X1 U5753 ( .A1(n4472), .A2(\DP/RegME_out[18] ), .ZN(n4445) );
  OAI211_X1 U5754 ( .C1(n4756), .C2(n4475), .A(n4445), .B(n4473), .ZN(
        DRAM_DATA_OUT[18]) );
  NAND2_X1 U5755 ( .A1(n4472), .A2(\DP/RegME_out[19] ), .ZN(n4447) );
  OAI211_X1 U5756 ( .C1(n4448), .C2(n4475), .A(n4447), .B(n4473), .ZN(
        DRAM_DATA_OUT[19]) );
  NAND2_X1 U5757 ( .A1(n4472), .A2(\DP/RegME_out[20] ), .ZN(n4449) );
  OAI211_X1 U5758 ( .C1(n4450), .C2(n4475), .A(n4449), .B(n4473), .ZN(
        DRAM_DATA_OUT[20]) );
  NAND2_X1 U5759 ( .A1(n4472), .A2(\DP/RegME_out[21] ), .ZN(n4451) );
  OAI211_X1 U5760 ( .C1(n4554), .C2(n4475), .A(n4451), .B(n4473), .ZN(
        DRAM_DATA_OUT[21]) );
  NAND2_X1 U5761 ( .A1(n4472), .A2(\DP/RegME_out[22] ), .ZN(n4453) );
  OAI211_X1 U5762 ( .C1(n4454), .C2(n4475), .A(n4453), .B(n4473), .ZN(
        DRAM_DATA_OUT[22]) );
  AOI22_X1 U5763 ( .A1(\DP/RegME_out[23] ), .A2(n4472), .B1(n4458), .B2(n4455), 
        .ZN(n4456) );
  NAND2_X1 U5764 ( .A1(n4456), .A2(n4473), .ZN(DRAM_DATA_OUT[23]) );
  AOI22_X1 U5765 ( .A1(\DP/RegME_out[24] ), .A2(n4472), .B1(n4458), .B2(n4457), 
        .ZN(n4459) );
  NAND2_X1 U5766 ( .A1(n4459), .A2(n4473), .ZN(DRAM_DATA_OUT[24]) );
  NAND2_X1 U5767 ( .A1(n4472), .A2(\DP/RegME_out[25] ), .ZN(n4460) );
  OAI211_X1 U5768 ( .C1(n4557), .C2(n4475), .A(n4460), .B(n4473), .ZN(
        DRAM_DATA_OUT[25]) );
  NAND2_X1 U5769 ( .A1(n4472), .A2(\DP/RegME_out[26] ), .ZN(n4462) );
  OAI211_X1 U5770 ( .C1(n4463), .C2(n4475), .A(n4462), .B(n4473), .ZN(
        DRAM_DATA_OUT[26]) );
  NAND2_X1 U5771 ( .A1(n4472), .A2(\DP/RegME_out[27] ), .ZN(n4464) );
  OAI211_X1 U5772 ( .C1(n4550), .C2(n4475), .A(n4464), .B(n4473), .ZN(
        DRAM_DATA_OUT[27]) );
  NAND2_X1 U5773 ( .A1(n4472), .A2(\DP/RegME_out[28] ), .ZN(n4466) );
  NAND2_X1 U5775 ( .A1(n4472), .A2(\DP/RegME_out[29] ), .ZN(n4468) );
  OAI211_X1 U5776 ( .C1(n4469), .C2(n4475), .A(n4468), .B(n4473), .ZN(
        DRAM_DATA_OUT[29]) );
  NAND2_X1 U5777 ( .A1(n4472), .A2(\DP/RegME_out[30] ), .ZN(n4470) );
  NAND2_X1 U5779 ( .A1(n4472), .A2(\DP/RegME_out[31] ), .ZN(n4474) );
  OAI211_X1 U5780 ( .C1(n4549), .C2(n4475), .A(n4474), .B(n4473), .ZN(
        DRAM_DATA_OUT[31]) );
  NAND2_X1 U5781 ( .A1(n4490), .A2(n4489), .ZN(n4488) );
  INV_X1 U5782 ( .A(n4488), .ZN(n4477) );
  NOR2_X1 U5783 ( .A1(n4478), .A2(n4477), .ZN(DRAM_DATA_OUT[7]) );
  AOI21_X1 U5784 ( .B1(n4482), .B2(\DP/RegME_out[8] ), .A(n4481), .ZN(n4479)
         );
  OAI21_X1 U5785 ( .B1(n4548), .B2(n4484), .A(n4479), .ZN(DRAM_DATA_OUT[8]) );
  AOI21_X1 U5786 ( .B1(n4482), .B2(\DP/RegME_out[9] ), .A(n4481), .ZN(n4483)
         );
  OAI21_X1 U5787 ( .B1(n4551), .B2(n4484), .A(n4483), .ZN(DRAM_DATA_OUT[9]) );
  NAND2_X1 U5788 ( .A1(n4486), .A2(n2374), .ZN(n4487) );
  NOR2_X1 U5789 ( .A1(n218), .A2(n4487), .ZN(n2339) );
  NAND2_X1 U5790 ( .A1(\DP/FwdD ), .A2(n4488), .ZN(n4521) );
  AOI21_X1 U5791 ( .B1(n4490), .B2(n4489), .A(\DP/FwdD ), .ZN(n4518) );
  NAND2_X1 U5792 ( .A1(\DP/RegME_out[3] ), .A2(n4518), .ZN(n4491) );
  OAI21_X1 U5793 ( .B1(n4521), .B2(n4492), .A(n4491), .ZN(DRAM_DATA_OUT[3]) );
  NAND2_X1 U5794 ( .A1(\DP/RegME_out[2] ), .A2(n4518), .ZN(n4493) );
  OAI21_X1 U5795 ( .B1(n4521), .B2(n4494), .A(n4493), .ZN(DRAM_DATA_OUT[2]) );
  INV_X1 U5796 ( .A(\DP/A[2] ), .ZN(n4500) );
  OAI221_X1 U5797 ( .B1(n4497), .B2(n4496), .C1(n4497), .C2(
        \DP/ALU0/MULT/SHIFTERi_0/N19 ), .A(n4495), .ZN(n4499) );
  OAI22_X1 U5798 ( .A1(n4515), .A2(n4500), .B1(n4499), .B2(n2439), .ZN(n196)
         );
  NAND2_X1 U5799 ( .A1(\DP/RegME_out[1] ), .A2(n4518), .ZN(n4501) );
  OAI21_X1 U5800 ( .B1(n4521), .B2(n4502), .A(n4501), .ZN(DRAM_DATA_OUT[1]) );
  NAND2_X1 U5801 ( .A1(\DP/RegME_out[0] ), .A2(n4518), .ZN(n4503) );
  OAI21_X1 U5802 ( .B1(n4521), .B2(n4504), .A(n4503), .ZN(DRAM_DATA_OUT[0]) );
  NAND2_X1 U5803 ( .A1(\DP/RegME_out[4] ), .A2(n4518), .ZN(n4505) );
  OAI21_X1 U5804 ( .B1(n4521), .B2(n4561), .A(n4505), .ZN(DRAM_DATA_OUT[4]) );
  INV_X1 U5805 ( .A(\DP/A[4] ), .ZN(n4514) );
  AOI221_X1 U5806 ( .B1(n4511), .B2(n4510), .C1(n4509), .C2(n4508), .A(n4507), 
        .ZN(n4513) );
  OAI22_X1 U5807 ( .A1(n4515), .A2(n4514), .B1(n4513), .B2(n4512), .ZN(n189)
         );
  NAND2_X1 U5808 ( .A1(\DP/RegME_out[5] ), .A2(n4518), .ZN(n4516) );
  OAI21_X1 U5809 ( .B1(n4521), .B2(n4517), .A(n4516), .ZN(DRAM_DATA_OUT[5]) );
  NAND2_X1 U5810 ( .A1(\DP/RegME_out[6] ), .A2(n4518), .ZN(n4519) );
  OAI21_X1 U5811 ( .B1(n4521), .B2(n4520), .A(n4519), .ZN(DRAM_DATA_OUT[6]) );
  INV_X1 U5812 ( .A(n107), .ZN(n4523) );
  AOI221_X1 U5813 ( .B1(n106), .B2(n107), .C1(\DP/A[31] ), .C2(n4523), .A(
        n4522), .ZN(n105) );
  REGISTER_FILE_WIDTH32_LENGTH5 \DP/RF0  ( .CLK(CLK), .RST(RST), .EN(w_WB_EN), 
        .RD1(w_RF_RD1), .RD2(n66), .WR(w_RF_WE), .DATAIN({\DP/RF_DATA[31] , 
        \DP/RF_DATA[30] , \DP/RF_DATA[29] , \DP/RF_DATA[28] , \DP/RF_DATA[27] , 
        \DP/RF_DATA[26] , \DP/RF_DATA[25] , \DP/RF_DATA[24] , \DP/RF_DATA[23] , 
        \DP/RF_DATA[22] , n4539, \DP/RF_DATA[20] , \DP/RF_DATA[19] , 
        \DP/RF_DATA[18] , \DP/RF_DATA[17] , \DP/RF_DATA[16] , \DP/RF_DATA[15] , 
        \DP/RF_DATA[14] , \DP/RF_DATA[13] , \DP/RF_DATA[12] , \DP/RF_DATA[11] , 
        \DP/RF_DATA[10] , \DP/RF_DATA[9] , \DP/RF_DATA[8] , \DP/RF_DATA[7] , 
        \DP/RF_DATA[6] , \DP/RF_DATA[5] , \DP/RF_DATA[4] , \DP/RF_DATA[3] , 
        \DP/RF_DATA[2] , \DP/RF_DATA[1] , \DP/RF_DATA[0] }), .OUT1({
        \DP/RegA_in[31] , \DP/RegA_in[30] , \DP/RegA_in[29] , \DP/RegA_in[28] , 
        \DP/RegA_in[27] , \DP/RegA_in[26] , \DP/RegA_in[25] , \DP/RegA_in[24] , 
        \DP/RegA_in[23] , \DP/RegA_in[22] , \DP/RegA_in[21] , \DP/RegA_in[20] , 
        \DP/RegA_in[19] , \DP/RegA_in[18] , \DP/RegA_in[17] , \DP/RegA_in[16] , 
        \DP/RegA_in[15] , \DP/RegA_in[14] , \DP/RegA_in[13] , \DP/RegA_in[12] , 
        \DP/RegA_in[11] , \DP/RegA_in[10] , \DP/RegA_in[9] , \DP/RegA_in[8] , 
        \DP/RegA_in[7] , \DP/RegA_in[6] , \DP/RegA_in[5] , \DP/RegA_in[4] , 
        \DP/RegA_in[3] , \DP/RegA_in[2] , \DP/RegA_in[1] , \DP/RegA_in[0] }), 
        .OUT2({\DP/RegB_in[31] , \DP/RegB_in[30] , \DP/RegB_in[29] , 
        \DP/RegB_in[28] , \DP/RegB_in[27] , \DP/RegB_in[26] , \DP/RegB_in[25] , 
        \DP/RegB_in[24] , \DP/RegB_in[23] , \DP/RegB_in[22] , \DP/RegB_in[21] , 
        \DP/RegB_in[20] , \DP/RegB_in[19] , \DP/RegB_in[18] , \DP/RegB_in[17] , 
        \DP/RegB_in[16] , \DP/RegB_in[15] , \DP/RegB_in[14] , \DP/RegB_in[13] , 
        \DP/RegB_in[12] , \DP/RegB_in[11] , \DP/RegB_in[10] , \DP/RegB_in[9] , 
        \DP/RegB_in[8] , \DP/RegB_in[7] , \DP/RegB_in[6] , \DP/RegB_in[5] , 
        \DP/RegB_in[4] , \DP/RegB_in[3] , \DP/RegB_in[2] , \DP/RegB_in[1] , 
        \DP/RegB_in[0] }), .ADD_WR({\DP/RF_ADDR[4] , \DP/RF_ADDR[3] , 
        \DP/RF_ADDR[2] , \DP/RF_ADDR[1] , \DP/RF_ADDR[0] }), .ADD_RD1({n104, 
        n103, n102, n101, n100}), .ADD_RD2({n97, n99, n94, n4646, n98}) );
  SNPS_CLOCK_GATE_HIGH_FFD_0 \DP/FFDBRANCH/clk_gate_Q_reg  ( .CLK(CLK), .EN(
        \DP/FFDBRANCH/N2 ), .ENCLK(\DP/FFDBRANCH/net2330 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_12 \DP/RegNPC/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\PC/N2 ), .ENCLK(\DP/RegNPC/net2366 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_11 \DP/RegNPC1/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegNPC1/N2 ), .ENCLK(\DP/RegNPC1/net2366 ), .TE(
        1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_10 \DP/RegA/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegA/N2 ), .ENCLK(\DP/RegA/net2366 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_9 \DP/RegB/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegB/N2 ), .ENCLK(\DP/RegB/net2366 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_7 \DP/RegA1/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegA1/N2 ), .ENCLK(\DP/RegA1/net2366 ), .TE(1'b0)
         );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_6 \DP/RegNPC2/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegNPC2/N2 ), .ENCLK(\DP/RegNPC2/net2366 ), .TE(
        1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_5 \DP/RegALU1/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegALU1/N2 ), .ENCLK(\DP/RegALU1/net2366 ), .TE(
        1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_2 \DP/RegLMD/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(n2461), .ENCLK(\DP/RegLMD/net2366 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_FFD_2 \DP/FFDJL2/clk_gate_Q_reg  ( .CLK(CLK), .EN(
        \DP/FFDJL2/N2 ), .ENCLK(\DP/FFDJL2/net2330 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_REGISTER_GENERIC_WIDTH32_1 \DP/RegNPC3/clk_gate_DOUT_reg  ( 
        .CLK(CLK), .EN(\DP/RegNPC3/N2 ), .ENCLK(\DP/RegNPC3/net2366 ), .TE(
        1'b0) );
  DFF_X2 \DP/FFDJL2/Q_reg  ( .D(\DP/FFDJL2/N3 ), .CK(\DP/FFDJL2/net2330 ), .Q(
        \DP/JL2 ) );
  OAI21_X2 U4631 ( .B1(\DP/JL2 ), .B2(n4444), .A(n3631), .ZN(\DP/RF_DATA[17] )
         );
  OAI21_X2 U4629 ( .B1(\DP/JL2 ), .B2(n4442), .A(n3630), .ZN(\DP/RF_DATA[16] )
         );
  AOI221_X2 U3353 ( .B1(n2471), .B2(n2525), .C1(n2491), .C2(n2525), .A(n2470), 
        .ZN(n2553) );
  CLKBUF_X3 U3241 ( .A(\DP/JL2 ), .Z(n2458) );
  NAND2_X2 U4633 ( .A1(n2459), .A2(\DP/NPC_out[19] ), .ZN(n3633) );
  BUF_X2 U3287 ( .A(\DP/JL2 ), .Z(n2459) );
  AOI21_X2 U3394 ( .B1(IR_OUT[30]), .B2(n2497), .A(n2496), .ZN(n3652) );
  DFF_X1 \CU/cw2_reg[9]  ( .D(\CU/N66 ), .CK(CLK), .Q(n2403), .QN(n206) );
  DFF_X1 \CU/cw2_reg[8]  ( .D(\CU/N65 ), .CK(CLK), .Q(n2399), .QN(n205) );
  DFF_X1 \CU/cw2_reg[4]  ( .D(\CU/N61 ), .CK(CLK), .Q(w_LOAD_SIZE[1]), .QN(
        n2369) );
  DFF_X1 \CU/cw2_reg[3]  ( .D(\CU/N60 ), .CK(CLK), .Q(n2400), .QN(n202) );
  DFF_X1 \DP/RegRD2/DOUT_reg[3]  ( .D(\DP/RegRD2/N6 ), .CK(n2452), .Q(n2385), 
        .QN(n400) );
  DFF_X1 \DP/RegRD2/DOUT_reg[2]  ( .D(\DP/RegRD2/N5 ), .CK(n2452), .Q(
        \DP/RD2[2] ), .QN(n2367) );
  DFF_X1 \DP/RegRD2/DOUT_reg[4]  ( .D(\DP/RegRD2/N7 ), .CK(n2452), .Q(n2365), 
        .QN(n401) );
  DFF_X1 \CU/cw1_reg[12]  ( .D(\CU/N50 ), .CK(CLK), .Q(w_JUMP_LINK), .QN(n2392) );
  DFF_X1 \DP/RegRD1/DOUT_reg[3]  ( .D(\DP/RegRD1/N6 ), .CK(n2452), .Q(
        \DP/RD1[3] ), .QN(n4635) );
  DFF_X1 \DP/RegRD1/DOUT_reg[2]  ( .D(\DP/RegRD1/N5 ), .CK(n2452), .Q(
        \DP/RD1[2] ), .QN(n2380) );
  DFF_X1 \DP/RegRD1/DOUT_reg[1]  ( .D(\DP/RegRD1/N4 ), .CK(n2452), .Q(
        \DP/RD1[1] ), .QN(n2378) );
  DFF_X1 \CU/cw1_reg[17]  ( .D(\CU/N55 ), .CK(CLK), .Q(w_MuxA_SEL), .QN(n2406)
         );
  DFF_X1 \CU/cw1_reg[16]  ( .D(\CU/N54 ), .CK(CLK), .Q(w_MuxB_SEL), .QN(n2407)
         );
  DFF_X1 \DP/FFDFD/Q_reg  ( .D(\DP/FFDFD/N3 ), .CK(\DP/RegNPC1/net2366 ), .Q(
        \DP/FwdD ), .QN(n2402) );
  DFF_X1 \DP/RegALU1/DOUT_reg[24]  ( .D(\DP/RegALU1/N27 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[24] ), .QN(n2393) );
  DFF_X1 \DP/RegFC/DOUT_reg[2]  ( .D(\DP/RegFC/N5 ), .CK(\DP/RegNPC1/net2366 ), 
        .Q(n2398), .QN(n407) );
  DFF_X1 \DP/RegALU1/DOUT_reg[23]  ( .D(\DP/RegALU1/N26 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[23] ), .QN(n2366) );
  DFF_X1 \DP/RegFC/DOUT_reg[1]  ( .D(\DP/RegFC/N4 ), .CK(\DP/RegNPC1/net2366 ), 
        .Q(\DP/FwdC[1] ), .QN(n2401) );
  DFF_X1 \CU/aluOpcode1_reg[4]  ( .D(\CU/N79 ), .CK(CLK), .Q(w_ALU_OPCODE[4]), 
        .QN(n2376) );
  DFF_X2 \DP/RegALU1/DOUT_reg[21]  ( .D(\DP/RegALU1/N24 ), .CK(
        \DP/RegALU1/net2366 ), .Q(\DP/RegALU1_out[21] ) );
  DFF_X2 \PC/DOUT_reg[28]  ( .D(\PC/N31 ), .CK(\DP/RegNPC/net2366 ), .Q(
        w_PC_OUT[28]) );
  DFF_X2 \DP/RegFC/DOUT_reg[0]  ( .D(\DP/RegFC/N3 ), .CK(\DP/RegNPC1/net2366 ), 
        .Q(n2370), .QN(n406) );
  DFF_X2 \DP/RegFB/DOUT_reg[2]  ( .D(\DP/RegFB/N5 ), .CK(\DP/RegNPC1/net2366 ), 
        .QN(n405) );
  DFFRS_X1 \DP/RegALU1/DOUT_reg[20]  ( .D(\DP/RegALU1/N23 ), .CK(
        \DP/RegALU1/net2366 ), .RN(1'b1), .SN(1'b1), .Q(\DP/RegALU1_out[20] )
         );
  DFF_X1 \CU/aluOpcode1_reg[1]  ( .D(\CU/N76 ), .CK(CLK), .Q(n2373), .QN(n4744) );
  DFF_X2 \CU/cw3_reg[1]  ( .D(\CU/N70 ), .CK(CLK), .Q(n2360), .QN(n200) );
  DFF_X2 \DP/RegNPC/DOUT_reg[31]  ( .D(n4530), .CK(\DP/RegNPC/net2366 ), .Q(
        \DP/NPC1[31] ) );
  DFF_X2 \PC/DOUT_reg[31]  ( .D(\PC/N34 ), .CK(n2456), .Q(w_PC_OUT[31]) );
  CLKBUF_X1 U3065 ( .A(n3615), .Z(n4524) );
  INV_X1 U3068 ( .A(n2464), .ZN(n4525) );
  OAI21_X1 U3071 ( .B1(\DP/JL2 ), .B2(n4448), .A(n3633), .ZN(\DP/RF_DATA[19] )
         );
  INV_X2 U3073 ( .A(n4175), .ZN(n4234) );
  CLKBUF_X1 U3093 ( .A(n2469), .Z(n4526) );
  AND2_X1 U3154 ( .A1(n2487), .A2(n2481), .ZN(n2502) );
  NAND2_X1 U3168 ( .A1(n2527), .A2(n2394), .ZN(n4527) );
  AND2_X1 U3169 ( .A1(n2514), .A2(n4793), .ZN(n4528) );
  NOR3_X1 U3170 ( .A1(n4708), .A2(n2550), .A3(n4707), .ZN(n2514) );
  CLKBUF_X1 U3171 ( .A(n2566), .Z(n4529) );
  OAI21_X1 U3172 ( .B1(n4395), .B2(n2381), .A(n4394), .ZN(n4530) );
  OR2_X2 U3173 ( .A1(n4315), .A2(n4787), .ZN(n4531) );
  CLKBUF_X1 U3174 ( .A(\CU/JUMP2 ), .Z(n4532) );
  INV_X1 U3175 ( .A(IROM_ADDR[4]), .ZN(n4917) );
  INV_X1 U3176 ( .A(IR_OUT[29]), .ZN(n4818) );
  NOR2_X1 U3177 ( .A1(IR_OUT[29]), .A2(IR_OUT[31]), .ZN(n4819) );
  AND2_X1 U3178 ( .A1(n4854), .A2(w_PC_OUT[13]), .ZN(n4333) );
  OAI21_X1 U3180 ( .B1(n4899), .B2(w_PC_OUT[25]), .A(n4801), .ZN(n4800) );
  NOR2_X1 U3181 ( .A1(n4375), .A2(n4802), .ZN(n4801) );
  NAND2_X1 U3182 ( .A1(n4856), .A2(w_PC_OUT[12]), .ZN(n4855) );
  OR2_X1 U3183 ( .A1(n4531), .A2(n4869), .ZN(n4393) );
  NOR2_X1 U3184 ( .A1(n4531), .A2(n4836), .ZN(n4835) );
  NOR2_X1 U3190 ( .A1(n4531), .A2(n4839), .ZN(n4380) );
  OAI21_X1 U3191 ( .B1(n4531), .B2(n4827), .A(n4834), .ZN(n4833) );
  AND2_X1 U3194 ( .A1(n4316), .A2(IROM_ADDR[9]), .ZN(n4319) );
  AND2_X1 U3200 ( .A1(n4316), .A2(n4665), .ZN(n4375) );
  NAND2_X1 U3207 ( .A1(n4316), .A2(n4849), .ZN(n4322) );
  AND2_X1 U3226 ( .A1(n4316), .A2(n4803), .ZN(n4669) );
  CLKBUF_X2 U3235 ( .A(n4399), .Z(n4560) );
  AND2_X1 U3236 ( .A1(n4853), .A2(w_PC_OUT[17]), .ZN(n4347) );
  CLKBUF_X1 U3237 ( .A(n3653), .Z(n4533) );
  AND3_X1 U3238 ( .A1(n4547), .A2(n4528), .A3(n2553), .ZN(n3653) );
  CLKBUF_X1 U3240 ( .A(n4789), .Z(n4534) );
  INV_X1 U3242 ( .A(n4536), .ZN(n4535) );
  AND3_X1 U3250 ( .A1(n3653), .A2(n2515), .A3(n2505), .ZN(n3615) );
  AND2_X1 U3253 ( .A1(n2530), .A2(n4753), .ZN(n2525) );
  INV_X2 U3259 ( .A(n2434), .ZN(n2433) );
  NAND2_X1 U3260 ( .A1(n4546), .A2(n4616), .ZN(n2530) );
  INV_X1 U3261 ( .A(n2547), .ZN(n2462) );
  AND2_X2 U3262 ( .A1(n2547), .A2(n4710), .ZN(n2528) );
  INV_X1 U3281 ( .A(n2553), .ZN(n4790) );
  NAND2_X1 U3283 ( .A1(n2479), .A2(n4678), .ZN(n4677) );
  AND2_X1 U3300 ( .A1(n2479), .A2(n4676), .ZN(n2546) );
  AND2_X1 U3306 ( .A1(n2479), .A2(n4673), .ZN(n4710) );
  AND2_X1 U3309 ( .A1(n2479), .A2(n4674), .ZN(n2526) );
  NAND2_X1 U3312 ( .A1(n4826), .A2(n4715), .ZN(n2478) );
  NOR3_X1 U3313 ( .A1(IR_OUT[30]), .A2(n4814), .A3(n2397), .ZN(n4715) );
  INV_X1 U3314 ( .A(n4818), .ZN(n4814) );
  NOR3_X1 U3315 ( .A1(n2533), .A2(n4792), .A3(n4790), .ZN(n2504) );
  AND2_X2 U3316 ( .A1(n4671), .A2(n4670), .ZN(n2479) );
  BUF_X2 U3318 ( .A(n200), .Z(n2449) );
  NOR2_X1 U3319 ( .A1(IR_OUT[30]), .A2(IR_OUT[27]), .ZN(n4678) );
  CLKBUF_X1 U3321 ( .A(IR_OUT[27]), .Z(n4559) );
  CLKBUF_X1 U3323 ( .A(n2530), .Z(n4566) );
  CLKBUF_X1 U3330 ( .A(n2508), .Z(n4555) );
  AND2_X2 U3335 ( .A1(n4537), .A2(n4538), .ZN(n4546) );
  BUF_X1 U3337 ( .A(\DP/RF_DATA[21] ), .Z(n4539) );
  OAI21_X1 U3338 ( .B1(n4452), .B2(\DP/JL2 ), .A(n3636), .ZN(\DP/RF_DATA[21] )
         );
  OR2_X1 U3340 ( .A1(n4438), .A2(n2458), .ZN(n4543) );
  AOI21_X1 U3341 ( .B1(\DP/RegLMD_out[14] ), .B2(n2448), .A(n4541), .ZN(n4438)
         );
  INV_X1 U3343 ( .A(n4544), .ZN(n4541) );
  CLKBUF_X1 U3344 ( .A(n4438), .Z(n4542) );
  NAND2_X1 U3345 ( .A1(n3628), .A2(n4543), .ZN(\DP/RF_DATA[14] ) );
  NAND2_X1 U3346 ( .A1(\DP/RegALU2_out[14] ), .A2(n200), .ZN(n4544) );
  INV_X2 U3347 ( .A(n200), .ZN(n2448) );
  INV_X2 U3349 ( .A(n2387), .ZN(n2446) );
  AND2_X1 U3354 ( .A1(n2387), .A2(n4545), .ZN(n4073) );
  NAND2_X2 U3356 ( .A1(n4074), .A2(n4072), .ZN(n4545) );
  OR2_X2 U3357 ( .A1(n3577), .A2(\DP/ALU0/N88 ), .ZN(n2387) );
  NOR2_X2 U3358 ( .A1(n3575), .A2(n3576), .ZN(n3577) );
  NAND3_X1 U3365 ( .A1(n4546), .A2(n4536), .A3(IR_OUT[29]), .ZN(n2467) );
  AND2_X2 U3366 ( .A1(n4546), .A2(n4536), .ZN(n4826) );
  NAND3_X1 U3367 ( .A1(n4546), .A2(n4536), .A3(IR_OUT[20]), .ZN(n4424) );
  NOR2_X1 U3382 ( .A1(n4789), .A2(n66), .ZN(n4547) );
  BUF_X1 U3383 ( .A(n4480), .Z(n4548) );
  BUF_X1 U3385 ( .A(n4476), .Z(n4549) );
  BUF_X2 U3395 ( .A(n4465), .Z(n4550) );
  BUF_X2 U3396 ( .A(n4485), .Z(n4551) );
  NAND2_X4 U3402 ( .A1(n4690), .A2(n3644), .ZN(\DP/RF_DATA[30] ) );
  INV_X1 U3423 ( .A(w_RF_RD1), .ZN(n4552) );
  NAND2_X1 U3427 ( .A1(n4552), .A2(RST), .ZN(\DP/RegA/N2 ) );
  BUF_X2 U3428 ( .A(n2483), .Z(n4553) );
  NAND2_X1 U3430 ( .A1(n4422), .A2(n2385), .ZN(n4661) );
  AND2_X1 U3435 ( .A1(n4662), .A2(n4661), .ZN(n4660) );
  BUF_X2 U3438 ( .A(n4452), .Z(n4554) );
  AOI21_X1 U3447 ( .B1(n2477), .B2(IR_OUT[27]), .A(n2478), .ZN(n2516) );
  NAND2_X1 U3459 ( .A1(n2527), .A2(n2394), .ZN(n2477) );
  NAND2_X1 U3461 ( .A1(n4574), .A2(n2372), .ZN(n2510) );
  NAND3_X1 U3475 ( .A1(n2566), .A2(n2510), .A3(n2531), .ZN(n4792) );
  BUF_X2 U3629 ( .A(n4436), .Z(n4556) );
  NAND2_X2 U3793 ( .A1(n4672), .A2(n3642), .ZN(\DP/RF_DATA[29] ) );
  BUF_X2 U3796 ( .A(n4461), .Z(n4557) );
  NAND2_X2 U3865 ( .A1(n2387), .A2(n4558), .ZN(n4178) );
  AND2_X2 U4012 ( .A1(RST), .A2(\DP/ALU0/s_LOGIC[2] ), .ZN(n4558) );
  AOI21_X1 U4313 ( .B1(n4619), .B2(n4617), .A(n4562), .ZN(\DP/FFDBRANCH/N3 )
         );
  NAND2_X2 U4316 ( .A1(n4615), .A2(n4614), .ZN(n4613) );
  NAND2_X1 U4353 ( .A1(n4613), .A2(n4598), .ZN(n4597) );
  BUF_X2 U4356 ( .A(n4506), .Z(n4561) );
  OR2_X2 U4445 ( .A1(n4815), .A2(n2461), .ZN(n4562) );
  NAND3_X1 U4529 ( .A1(n4656), .A2(n4660), .A3(n4563), .ZN(n3620) );
  INV_X2 U4540 ( .A(n4564), .ZN(n4563) );
  NOR2_X2 U4550 ( .A1(n4421), .A2(\DP/RD2[2] ), .ZN(n4564) );
  NAND2_X2 U4554 ( .A1(n3643), .A2(n4640), .ZN(\DP/RF_DATA[2] ) );
  BUF_X2 U4558 ( .A(n4432), .Z(n4565) );
  NAND2_X2 U4561 ( .A1(n3646), .A2(n4683), .ZN(\DP/RF_DATA[3] ) );
  NAND2_X2 U4564 ( .A1(n3637), .A2(n4685), .ZN(\DP/RF_DATA[22] ) );
  NAND2_X2 U4565 ( .A1(n3645), .A2(n4682), .ZN(\DP/RF_DATA[31] ) );
  NAND2_X2 U4566 ( .A1(n3651), .A2(n4687), .ZN(\DP/RF_DATA[9] ) );
  NAND2_X2 U4567 ( .A1(n3650), .A2(n4681), .ZN(\DP/RF_DATA[8] ) );
  INV_X2 U4568 ( .A(n2445), .ZN(n1110) );
  NAND2_X2 U4594 ( .A1(n2445), .A2(n4567), .ZN(n2396) );
  NOR2_X2 U4595 ( .A1(n2461), .A2(n4098), .ZN(n4567) );
  NAND2_X2 U4596 ( .A1(n4742), .A2(n4568), .ZN(n2445) );
  NAND2_X2 U4597 ( .A1(n4486), .A2(n2374), .ZN(n4568) );
  OR2_X2 U4599 ( .A1(n4743), .A2(n3810), .ZN(n4742) );
  NAND3_X1 U4600 ( .A1(n4735), .A2(n4734), .A3(n4246), .ZN(n4732) );
  NAND4_X2 U4601 ( .A1(n4243), .A2(n4733), .A3(n4739), .A4(n4569), .ZN(n4246)
         );
  AND2_X2 U4602 ( .A1(n4736), .A2(n4570), .ZN(n4569) );
  INV_X2 U4603 ( .A(n4571), .ZN(n4570) );
  OAI22_X2 U4604 ( .A1(n102), .A2(n2380), .B1(n4269), .B2(\DP/RD1[2] ), .ZN(
        n4571) );
  NOR3_X1 U4605 ( .A1(n2466), .A2(n2465), .A3(n2388), .ZN(n4574) );
  OR3_X1 U4606 ( .A1(n2466), .A2(n2465), .A3(n4572), .ZN(n4709) );
  NAND2_X1 U4609 ( .A1(n4573), .A2(n224), .ZN(n4572) );
  INV_X1 U4614 ( .A(n2388), .ZN(n4573) );
  INV_X1 U4621 ( .A(n4574), .ZN(n4576) );
  NOR2_X2 U4623 ( .A1(n2572), .A2(n4575), .ZN(n2579) );
  NAND2_X2 U4625 ( .A1(n4577), .A2(n4576), .ZN(n4575) );
  NAND2_X2 U4627 ( .A1(n2575), .A2(n2574), .ZN(n4577) );
  NOR2_X1 U4634 ( .A1(n2530), .A2(n224), .ZN(n2527) );
  NAND2_X2 U4636 ( .A1(n4579), .A2(n4578), .ZN(\DP/RF_DATA[7] ) );
  NAND2_X2 U4639 ( .A1(\DP/JL2 ), .A2(\DP/NPC_out[7] ), .ZN(n4578) );
  NAND2_X2 U4641 ( .A1(n4428), .A2(n4580), .ZN(n4579) );
  INV_X2 U4648 ( .A(\DP/JL2 ), .ZN(n4580) );
  NAND2_X2 U4650 ( .A1(n4698), .A2(n4581), .ZN(n4428) );
  NAND2_X2 U4652 ( .A1(n2448), .A2(\DP/RegLMD_out[7] ), .ZN(n4581) );
  NAND2_X2 U4654 ( .A1(n4701), .A2(n3640), .ZN(\DP/RF_DATA[27] ) );
  NOR2_X2 U4656 ( .A1(n2539), .A2(IR_OUT[4]), .ZN(n2556) );
  NAND2_X2 U4658 ( .A1(n2517), .A2(n4582), .ZN(n2571) );
  NOR2_X2 U4660 ( .A1(n2539), .A2(n4587), .ZN(n4582) );
  OAI22_X2 U4662 ( .A1(n4589), .A2(n4585), .B1(n2522), .B2(n4583), .ZN(n4590)
         );
  INV_X2 U4664 ( .A(n4584), .ZN(n4583) );
  NOR2_X2 U4665 ( .A1(n2523), .A2(n4593), .ZN(n4584) );
  INV_X2 U4666 ( .A(n4586), .ZN(n4585) );
  NOR3_X2 U4668 ( .A1(n2539), .A2(n4593), .A3(n4587), .ZN(n4586) );
  NAND2_X2 U4670 ( .A1(n4588), .A2(IR_OUT[5]), .ZN(n4587) );
  INV_X2 U4682 ( .A(IR_OUT[4]), .ZN(n4588) );
  INV_X2 U4716 ( .A(n2517), .ZN(n4589) );
  INV_X2 U4754 ( .A(n4590), .ZN(n2541) );
  OAI21_X2 U4758 ( .B1(n2571), .B2(n4593), .A(n4591), .ZN(n2540) );
  INV_X2 U4785 ( .A(n4592), .ZN(n4591) );
  NOR3_X2 U4819 ( .A1(n2522), .A2(n2523), .A3(n4593), .ZN(n4592) );
  INV_X2 U5194 ( .A(n4594), .ZN(n4593) );
  INV_X1 U5340 ( .A(IR_OUT[0]), .ZN(n4594) );
  NAND3_X1 U5341 ( .A1(n4430), .A2(n4438), .A3(n4595), .ZN(n4785) );
  NOR2_X2 U5342 ( .A1(n4613), .A2(n4596), .ZN(n4595) );
  INV_X2 U5343 ( .A(n4463), .ZN(n4596) );
  NAND2_X2 U5346 ( .A1(n3626), .A2(n4597), .ZN(\DP/RF_DATA[12] ) );
  INV_X2 U5349 ( .A(\DP/JL2 ), .ZN(n4598) );
  NAND2_X2 U5350 ( .A1(n3662), .A2(n4599), .ZN(\DP/RegA1/N15 ) );
  NAND2_X2 U5351 ( .A1(n4613), .A2(n4600), .ZN(n4599) );
  INV_X2 U5353 ( .A(n3693), .ZN(n4600) );
  NAND2_X2 U5359 ( .A1(n3452), .A2(n4601), .ZN(\DP/B[12] ) );
  NOR2_X2 U5365 ( .A1(n4605), .A2(n4602), .ZN(n4601) );
  INV_X2 U5366 ( .A(n4603), .ZN(n4602) );
  NAND2_X2 U5367 ( .A1(n4613), .A2(n4604), .ZN(n4603) );
  INV_X2 U5492 ( .A(n2418), .ZN(n4604) );
  INV_X2 U5493 ( .A(n3453), .ZN(n4605) );
  NAND2_X1 U5494 ( .A1(n2773), .A2(n4606), .ZN(\DP/A[12] ) );
  NOR2_X1 U5495 ( .A1(n4610), .A2(n4607), .ZN(n4606) );
  INV_X1 U5496 ( .A(n4608), .ZN(n4607) );
  NAND2_X1 U5501 ( .A1(n4613), .A2(n4609), .ZN(n4608) );
  INV_X1 U5504 ( .A(n2413), .ZN(n4609) );
  INV_X1 U5509 ( .A(n2774), .ZN(n4610) );
  NAND2_X2 U5512 ( .A1(n4433), .A2(n4611), .ZN(DRAM_DATA_OUT[12]) );
  NAND2_X2 U5517 ( .A1(n4613), .A2(n4612), .ZN(n4611) );
  INV_X2 U5520 ( .A(n4484), .ZN(n4612) );
  NAND2_X1 U5525 ( .A1(\DP/RegALU2_out[12] ), .A2(n200), .ZN(n4614) );
  NAND2_X2 U5528 ( .A1(n2448), .A2(\DP/RegLMD_out[12] ), .ZN(n4615) );
  INV_X2 U5533 ( .A(n4309), .ZN(n4415) );
  NAND2_X2 U5537 ( .A1(n4309), .A2(n4751), .ZN(n4315) );
  AND2_X2 U5542 ( .A1(n4416), .A2(IROM_ADDR[6]), .ZN(n4309) );
  AND2_X2 U5545 ( .A1(n4410), .A2(IROM_ADDR[5]), .ZN(n4416) );
  NOR2_X1 U5548 ( .A1(\CU/JUMP1 ), .A2(n2388), .ZN(n4616) );
  NOR2_X1 U5550 ( .A1(w_JUMP_LINK), .A2(n4618), .ZN(n4617) );
  NAND2_X1 U5551 ( .A1(n208), .A2(n207), .ZN(n4618) );
  XNOR2_X1 U5553 ( .A(n4621), .B(n4620), .ZN(n4619) );
  INV_X1 U5558 ( .A(w_JUMP_EQ), .ZN(n4620) );
  OAI21_X1 U5561 ( .B1(n4622), .B2(n3654), .A(n4746), .ZN(n4621) );
  NOR2_X1 U5566 ( .A1(n4778), .A2(n4749), .ZN(n4622) );
  INV_X1 U5569 ( .A(n4239), .ZN(n2434) );
  NAND2_X2 U5570 ( .A1(n2387), .A2(n4624), .ZN(n4239) );
  CLKBUF_X1 U5572 ( .A(n2387), .Z(n4623) );
  NOR2_X1 U5574 ( .A1(n4626), .A2(n4625), .ZN(n4624) );
  INV_X1 U5575 ( .A(RST), .ZN(n4625) );
  INV_X1 U5579 ( .A(\DP/ALU0/s_LOGIC[3] ), .ZN(n4626) );
  NAND2_X2 U5584 ( .A1(n3623), .A2(n4627), .ZN(\DP/RF_DATA[0] ) );
  NAND2_X2 U5585 ( .A1(n4629), .A2(n4628), .ZN(n4627) );
  INV_X2 U5587 ( .A(n2459), .ZN(n4628) );
  INV_X2 U5591 ( .A(n4504), .ZN(n4629) );
  NAND2_X2 U5592 ( .A1(n3647), .A2(n4630), .ZN(\DP/RF_DATA[4] ) );
  NAND2_X2 U5715 ( .A1(n4632), .A2(n4631), .ZN(n4630) );
  INV_X2 U5716 ( .A(\DP/JL2 ), .ZN(n4631) );
  INV_X2 U5717 ( .A(n4506), .ZN(n4632) );
  NAND4_X2 U5718 ( .A1(n4639), .A2(n4638), .A3(n4257), .A4(n4633), .ZN(n4261)
         );
  NOR2_X2 U5719 ( .A1(n4637), .A2(n4634), .ZN(n4633) );
  OAI22_X2 U5720 ( .A1(n4636), .A2(n4635), .B1(n4421), .B2(\DP/RD1[2] ), .ZN(
        n4634) );
  INV_X2 U5742 ( .A(n4422), .ZN(n4636) );
  OAI22_X2 U5774 ( .A1(n96), .A2(n2378), .B1(n4420), .B2(\DP/RD1[1] ), .ZN(
        n4637) );
  INV_X2 U5778 ( .A(n4420), .ZN(n96) );
  OR2_X2 U5814 ( .A1(n94), .A2(n2380), .ZN(n4638) );
  NAND2_X2 U5815 ( .A1(n99), .A2(n4635), .ZN(n4639) );
  INV_X1 U5816 ( .A(n4854), .ZN(n4329) );
  INV_X1 U5817 ( .A(n4853), .ZN(n4343) );
  NAND2_X1 U5818 ( .A1(n4642), .A2(n4641), .ZN(n4640) );
  INV_X1 U5819 ( .A(\DP/JL2 ), .ZN(n4641) );
  INV_X1 U5820 ( .A(n4494), .ZN(n4642) );
  NOR2_X2 U5821 ( .A1(n4822), .A2(n4655), .ZN(n2576) );
  OAI21_X2 U5822 ( .B1(n584), .B2(n4655), .A(n4643), .ZN(\DP/RegRD1/N3 ) );
  NAND2_X2 U5823 ( .A1(n4653), .A2(n4644), .ZN(n4643) );
  INV_X2 U5824 ( .A(n4419), .ZN(n4644) );
  OAI21_X2 U5825 ( .B1(n582), .B2(n4655), .A(n4645), .ZN(\DP/RegRD1/N4 ) );
  NAND2_X2 U5826 ( .A1(n4653), .A2(n4646), .ZN(n4645) );
  INV_X2 U5827 ( .A(n4420), .ZN(n4646) );
  OAI21_X2 U5828 ( .B1(n580), .B2(n4655), .A(n4647), .ZN(\DP/RegRD1/N5 ) );
  NAND2_X2 U5829 ( .A1(n4653), .A2(n4648), .ZN(n4647) );
  INV_X2 U5830 ( .A(n4421), .ZN(n4648) );
  OAI21_X2 U5831 ( .B1(n578), .B2(n4655), .A(n4649), .ZN(\DP/RegRD1/N6 ) );
  NAND2_X2 U5832 ( .A1(n4653), .A2(n4650), .ZN(n4649) );
  INV_X2 U5833 ( .A(n4422), .ZN(n4650) );
  OAI21_X2 U5834 ( .B1(n575), .B2(n4655), .A(n4651), .ZN(\DP/RegRD1/N7 ) );
  NAND2_X2 U5835 ( .A1(n4653), .A2(n4652), .ZN(n4651) );
  INV_X2 U5836 ( .A(n4424), .ZN(n4652) );
  NOR2_X2 U5837 ( .A1(n4726), .A2(n4654), .ZN(n4653) );
  INV_X2 U5838 ( .A(RST), .ZN(n4654) );
  INV_X2 U5839 ( .A(n4726), .ZN(n4655) );
  AND2_X2 U5840 ( .A1(n2502), .A2(n2525), .ZN(n4726) );
  INV_X2 U5841 ( .A(n4422), .ZN(n99) );
  INV_X2 U5842 ( .A(n4657), .ZN(n4656) );
  OAI211_X2 U5843 ( .C1(n4422), .C2(n2385), .A(n3616), .B(n4658), .ZN(n4657)
         );
  INV_X2 U5844 ( .A(n4659), .ZN(n4658) );
  OAI21_X2 U5845 ( .B1(n4419), .B2(\DP/RD2[0] ), .A(n4247), .ZN(n4659) );
  NAND2_X2 U5846 ( .A1(n4815), .A2(IR_OUT[19]), .ZN(n4422) );
  OR2_X2 U5847 ( .A1(n4420), .A2(\DP/RD2[1] ), .ZN(n4662) );
  NAND2_X2 U5848 ( .A1(n4815), .A2(n4718), .ZN(n4420) );
  OAI21_X1 U5849 ( .B1(n4316), .B2(w_PC_OUT[20]), .A(n4663), .ZN(n4668) );
  INV_X2 U5850 ( .A(n4664), .ZN(n4663) );
  OAI21_X2 U5851 ( .B1(n4803), .B2(w_PC_OUT[20]), .A(n2437), .ZN(n4664) );
  INV_X2 U5852 ( .A(n4666), .ZN(n4665) );
  NAND2_X2 U5853 ( .A1(n4803), .A2(n4831), .ZN(n4666) );
  AND2_X2 U5854 ( .A1(n4669), .A2(n4872), .ZN(n4368) );
  NAND2_X2 U5855 ( .A1(n4667), .A2(n4357), .ZN(n4355) );
  INV_X2 U5856 ( .A(n4668), .ZN(n4667) );
  OAI21_X2 U5857 ( .B1(n4353), .B2(n4669), .A(n4352), .ZN(\PC/N22 ) );
  INV_X1 U5858 ( .A(n2465), .ZN(n2509) );
  OR2_X1 U5859 ( .A1(n2479), .A2(n2371), .ZN(n2465) );
  NOR2_X1 U5860 ( .A1(\CU/JUMP2 ), .A2(n2394), .ZN(n4670) );
  NOR2_X1 U5861 ( .A1(\CU/JUMP3 ), .A2(\CU/JUMP1 ), .ZN(n4671) );
  OR2_X2 U5862 ( .A1(n4469), .A2(\DP/JL2 ), .ZN(n4672) );
  INV_X2 U5863 ( .A(IR_OUT[30]), .ZN(n4673) );
  NOR2_X2 U5864 ( .A1(IR_OUT[31]), .A2(n2371), .ZN(n4674) );
  NOR2_X2 U5865 ( .A1(n2466), .A2(n4675), .ZN(n2471) );
  INV_X2 U5866 ( .A(n2546), .ZN(n4675) );
  INV_X2 U5867 ( .A(n2371), .ZN(n4676) );
  NOR2_X2 U5868 ( .A1(n2488), .A2(n4677), .ZN(n2501) );
  AND2_X1 U5869 ( .A1(n2530), .A2(n4846), .ZN(n2574) );
  NOR3_X2 U5870 ( .A1(n4315), .A2(n4787), .A3(n4868), .ZN(n4358) );
  NOR3_X2 U5871 ( .A1(n4315), .A2(n4787), .A3(n4679), .ZN(n4361) );
  NAND2_X2 U5872 ( .A1(n4680), .A2(w_PC_OUT[21]), .ZN(n4679) );
  INV_X2 U5873 ( .A(n4868), .ZN(n4680) );
  OR2_X1 U5874 ( .A1(n4480), .A2(\DP/JL2 ), .ZN(n4681) );
  OR2_X1 U5875 ( .A1(n4476), .A2(\DP/JL2 ), .ZN(n4682) );
  INV_X1 U5876 ( .A(n4684), .ZN(n4683) );
  NOR2_X1 U5877 ( .A1(n4492), .A2(\DP/JL2 ), .ZN(n4684) );
  INV_X1 U5878 ( .A(n4686), .ZN(n4685) );
  NOR2_X1 U5879 ( .A1(n4454), .A2(\DP/JL2 ), .ZN(n4686) );
  OR2_X1 U5880 ( .A1(n4485), .A2(\DP/JL2 ), .ZN(n4687) );
  NAND4_X2 U5881 ( .A1(n4469), .A2(n4465), .A3(n4774), .A4(n4695), .ZN(n3588)
         );
  NAND2_X2 U5882 ( .A1(n3683), .A2(n4688), .ZN(\DP/RegA1/N33 ) );
  INV_X2 U5883 ( .A(n4689), .ZN(n4688) );
  NOR2_X2 U5884 ( .A1(n2423), .A2(n4695), .ZN(n4689) );
  OR2_X1 U5885 ( .A1(n4695), .A2(\DP/JL2 ), .ZN(n4690) );
  NAND2_X2 U5886 ( .A1(n3560), .A2(n4691), .ZN(n3561) );
  OR2_X2 U5887 ( .A1(n4695), .A2(n2417), .ZN(n4691) );
  NAND3_X1 U5888 ( .A1(n3370), .A2(n3371), .A3(n4692), .ZN(\DP/A[30] ) );
  OR2_X2 U5889 ( .A1(n4695), .A2(n2412), .ZN(n4692) );
  NAND2_X2 U5890 ( .A1(n4473), .A2(n4693), .ZN(DRAM_DATA_OUT[30]) );
  NOR2_X2 U5891 ( .A1(n4697), .A2(n4694), .ZN(n4693) );
  NOR2_X2 U5892 ( .A1(n4475), .A2(n4695), .ZN(n4694) );
  AOI21_X1 U5893 ( .B1(n2449), .B2(\DP/RegALU2_out[30] ), .A(n4696), .ZN(n4695) );
  AND2_X1 U5894 ( .A1(n2360), .A2(\DP/RegLMD_out[30] ), .ZN(n4696) );
  INV_X2 U5895 ( .A(n4470), .ZN(n4697) );
  NAND2_X2 U5896 ( .A1(n4723), .A2(n3648), .ZN(\DP/RF_DATA[5] ) );
  INV_X1 U5897 ( .A(n4428), .ZN(n3657) );
  NAND2_X1 U5898 ( .A1(\DP/RegALU2_out[7] ), .A2(n200), .ZN(n4698) );
  NAND2_X1 U5899 ( .A1(n3639), .A2(n4699), .ZN(\DP/RF_DATA[26] ) );
  OR2_X1 U5900 ( .A1(n2458), .A2(n4463), .ZN(n4699) );
  NAND2_X1 U5901 ( .A1(n3635), .A2(n4700), .ZN(\DP/RF_DATA[20] ) );
  OR2_X1 U5902 ( .A1(n2458), .A2(n4450), .ZN(n4700) );
  OR2_X1 U5903 ( .A1(n4465), .A2(n2458), .ZN(n4701) );
  NAND2_X1 U5904 ( .A1(n3625), .A2(n4702), .ZN(\DP/RF_DATA[11] ) );
  OR2_X1 U5905 ( .A1(n4432), .A2(n2458), .ZN(n4702) );
  NAND2_X2 U5906 ( .A1(n3634), .A2(n4703), .ZN(\DP/RF_DATA[1] ) );
  OR2_X2 U5907 ( .A1(n2459), .A2(n4502), .ZN(n4703) );
  NAND2_X2 U5908 ( .A1(n3629), .A2(n4704), .ZN(\DP/RF_DATA[15] ) );
  OR2_X2 U5909 ( .A1(n4440), .A2(n2459), .ZN(n4704) );
  NAND2_X2 U5910 ( .A1(n3627), .A2(n4705), .ZN(\DP/RF_DATA[13] ) );
  OR2_X2 U5911 ( .A1(n4436), .A2(n2459), .ZN(n4705) );
  NAND2_X2 U5912 ( .A1(n3638), .A2(n4706), .ZN(\DP/RF_DATA[25] ) );
  OR2_X2 U5913 ( .A1(n4461), .A2(n2459), .ZN(n4706) );
  AND2_X1 U5914 ( .A1(n2528), .A2(n2525), .ZN(n4707) );
  NOR2_X1 U5915 ( .A1(n2506), .A2(n4526), .ZN(n2550) );
  INV_X1 U5916 ( .A(n4709), .ZN(n4708) );
  NAND2_X1 U5917 ( .A1(n2508), .A2(n224), .ZN(n2506) );
  INV_X1 U5918 ( .A(n2530), .ZN(n2508) );
  BUF_X2 U5919 ( .A(n4816), .Z(n4711) );
  NAND2_X1 U5920 ( .A1(n4716), .A2(n4826), .ZN(n2487) );
  INV_X2 U5921 ( .A(n4826), .ZN(n4816) );
  NOR2_X1 U5922 ( .A1(n4722), .A2(n4712), .ZN(n3616) );
  NOR2_X1 U5923 ( .A1(n4713), .A2(n4826), .ZN(n4712) );
  INV_X1 U5924 ( .A(n4762), .ZN(n4713) );
  NAND2_X2 U5925 ( .A1(n4815), .A2(n4714), .ZN(\DP/FFDJL2/N2 ) );
  INV_X2 U5926 ( .A(\DP/RegNPC2/N2 ), .ZN(n4714) );
  INV_X2 U5927 ( .A(n4819), .ZN(n4716) );
  NAND2_X2 U5928 ( .A1(n4826), .A2(n4717), .ZN(n4419) );
  INV_X2 U5929 ( .A(n4758), .ZN(n4717) );
  INV_X2 U5930 ( .A(n4759), .ZN(n4718) );
  NOR2_X2 U5931 ( .A1(n4816), .A2(n2377), .ZN(n2512) );
  NOR2_X2 U5932 ( .A1(n4816), .A2(n2460), .ZN(n4275) );
  NOR2_X2 U5933 ( .A1(n4711), .A2(n4719), .ZN(n2519) );
  NAND2_X2 U5934 ( .A1(n4721), .A2(n4720), .ZN(n4719) );
  INV_X2 U5935 ( .A(n2382), .ZN(n4720) );
  INV_X2 U5936 ( .A(IR_OUT[2]), .ZN(n4721) );
  OAI21_X2 U5937 ( .B1(n2523), .B2(n4711), .A(n2349), .ZN(n2350) );
  OR2_X2 U5938 ( .A1(n4761), .A2(n4760), .ZN(n4722) );
  CLKBUF_X3 U5939 ( .A(n4826), .Z(n4815) );
  OR2_X1 U5940 ( .A1(n2459), .A2(n4517), .ZN(n4723) );
  NAND2_X2 U5941 ( .A1(n3624), .A2(n4724), .ZN(\DP/RF_DATA[10] ) );
  OR2_X2 U5942 ( .A1(n4430), .A2(n2458), .ZN(n4724) );
  NAND2_X2 U5943 ( .A1(n3649), .A2(n4725), .ZN(\DP/RF_DATA[6] ) );
  OR2_X2 U5944 ( .A1(n2458), .A2(n4520), .ZN(n4725) );
  NAND2_X1 U5945 ( .A1(n2485), .A2(n2511), .ZN(n66) );
  NAND2_X1 U5946 ( .A1(n4726), .A2(n4824), .ZN(n2485) );
  NOR2_X1 U5947 ( .A1(n4731), .A2(n4727), .ZN(n2355) );
  NAND4_X1 U5948 ( .A1(n4730), .A2(n2514), .A3(n4729), .A4(n2515), .ZN(n4727)
         );
  AND2_X1 U5949 ( .A1(n3652), .A2(n4728), .ZN(n2515) );
  NAND2_X1 U5950 ( .A1(n2502), .A2(n4555), .ZN(n4728) );
  NOR2_X1 U5951 ( .A1(n2354), .A2(n2516), .ZN(n4729) );
  INV_X1 U5952 ( .A(n2346), .ZN(n4730) );
  NOR2_X1 U5953 ( .A1(n2352), .A2(n2537), .ZN(n4731) );
  NOR2_X1 U5954 ( .A1(n4732), .A2(n4251), .ZN(n4254) );
  OR2_X1 U5955 ( .A1(n103), .A2(n4635), .ZN(n4733) );
  INV_X1 U5956 ( .A(n4250), .ZN(n4734) );
  INV_X1 U5957 ( .A(n4252), .ZN(n4735) );
  AOI22_X1 U5958 ( .A1(n4738), .A2(n4737), .B1(\DP/RD1[1] ), .B2(n4268), .ZN(
        n4736) );
  INV_X1 U5959 ( .A(\DP/RD1[3] ), .ZN(n4737) );
  INV_X1 U5960 ( .A(n4270), .ZN(n4738) );
  NAND2_X1 U5961 ( .A1(n101), .A2(n2378), .ZN(n4739) );
  INV_X2 U5962 ( .A(n4742), .ZN(n2341) );
  CLKBUF_X1 U5963 ( .A(n1110), .Z(n4740) );
  NAND2_X1 U5964 ( .A1(n2445), .A2(n4741), .ZN(n4175) );
  AND2_X2 U5965 ( .A1(RST), .A2(n4098), .ZN(n4741) );
  NAND2_X2 U5966 ( .A1(n4745), .A2(n4744), .ZN(n4743) );
  INV_X2 U5967 ( .A(w_ALU_OPCODE[2]), .ZN(n4745) );
  NOR2_X1 U5968 ( .A1(n4748), .A2(n4747), .ZN(n4746) );
  INV_X1 U5969 ( .A(n3609), .ZN(n4747) );
  INV_X1 U5970 ( .A(n3610), .ZN(n4748) );
  NAND4_X1 U5971 ( .A1(n4777), .A2(n4781), .A3(n4786), .A4(n4750), .ZN(n4749)
         );
  NOR3_X1 U5972 ( .A1(n3579), .A2(n4457), .A3(n4455), .ZN(n4750) );
  INV_X2 U5973 ( .A(n4315), .ZN(n4316) );
  NAND3_X1 U5974 ( .A1(n4309), .A2(n4751), .A3(n4797), .ZN(n4364) );
  AND2_X2 U5975 ( .A1(n4309), .A2(IROM_ADDR[7]), .ZN(n4312) );
  AND2_X2 U5976 ( .A1(IROM_ADDR[7]), .A2(IROM_ADDR[8]), .ZN(n4751) );
  NOR2_X2 U5977 ( .A1(n4907), .A2(n4752), .ZN(n4906) );
  INV_X2 U5978 ( .A(w_PC_OUT[25]), .ZN(n4752) );
  INV_X2 U5979 ( .A(n2372), .ZN(n4753) );
  INV_X2 U5980 ( .A(n4909), .ZN(n4908) );
  NOR2_X2 U5981 ( .A1(n4754), .A2(n4909), .ZN(n4898) );
  INV_X2 U5982 ( .A(n4914), .ZN(n4754) );
  AND2_X2 U5983 ( .A1(w_PC_OUT[27]), .A2(w_PC_OUT[28]), .ZN(n4914) );
  OAI21_X2 U5984 ( .B1(n2459), .B2(n4446), .A(n3632), .ZN(\DP/RF_DATA[18] ) );
  AOI21_X2 U5985 ( .B1(\DP/RegLMD_out[18] ), .B2(n2448), .A(n4755), .ZN(n4446)
         );
  INV_X2 U5986 ( .A(n4757), .ZN(n4755) );
  CLKBUF_X1 U5987 ( .A(n4446), .Z(n4756) );
  NAND2_X1 U5988 ( .A1(\DP/RegALU2_out[18] ), .A2(n200), .ZN(n4757) );
  INV_X2 U5989 ( .A(IR_OUT[16]), .ZN(n4758) );
  INV_X2 U5990 ( .A(IR_OUT[17]), .ZN(n4759) );
  NOR2_X2 U5991 ( .A1(n4764), .A2(IR_OUT[16]), .ZN(n4760) );
  NOR2_X2 U5992 ( .A1(n4763), .A2(IR_OUT[17]), .ZN(n4761) );
  NAND2_X2 U5993 ( .A1(n4764), .A2(n4763), .ZN(n4762) );
  INV_X2 U5994 ( .A(\DP/RD2[1] ), .ZN(n4763) );
  INV_X2 U5995 ( .A(\DP/RD2[0] ), .ZN(n4764) );
  CLKBUF_X1 U5996 ( .A(n4419), .Z(n4765) );
  NAND2_X2 U5997 ( .A1(n3681), .A2(n4766), .ZN(\DP/RegA1/N31 ) );
  OR2_X2 U5998 ( .A1(n3693), .A2(n4774), .ZN(n4766) );
  NAND2_X2 U5999 ( .A1(n3641), .A2(n4767), .ZN(\DP/RF_DATA[28] ) );
  OR2_X2 U6000 ( .A1(n4774), .A2(\DP/JL2 ), .ZN(n4767) );
  NAND2_X1 U6001 ( .A1(n3326), .A2(n4768), .ZN(\DP/A[28] ) );
  NOR2_X1 U6002 ( .A1(n4770), .A2(n4769), .ZN(n4768) );
  NOR2_X1 U6003 ( .A1(n4774), .A2(n2412), .ZN(n4769) );
  INV_X1 U6004 ( .A(n3327), .ZN(n4770) );
  NAND2_X2 U6005 ( .A1(n3547), .A2(n4771), .ZN(n3548) );
  OR2_X2 U6006 ( .A1(n4774), .A2(n2417), .ZN(n4771) );
  NAND2_X2 U6007 ( .A1(n4473), .A2(n4772), .ZN(DRAM_DATA_OUT[28]) );
  NOR2_X2 U6008 ( .A1(n4776), .A2(n4773), .ZN(n4772) );
  NOR2_X2 U6009 ( .A1(n4475), .A2(n4774), .ZN(n4773) );
  AOI21_X1 U6010 ( .B1(n2449), .B2(\DP/RegALU2_out[28] ), .A(n4775), .ZN(n4774) );
  AND2_X1 U6011 ( .A1(n2360), .A2(\DP/RegLMD_out[28] ), .ZN(n4775) );
  INV_X2 U6012 ( .A(n4466), .ZN(n4776) );
  INV_X1 U6013 ( .A(n3583), .ZN(n4781) );
  AND2_X2 U6014 ( .A1(n4783), .A2(n4784), .ZN(n4777) );
  NAND3_X1 U6015 ( .A1(n4782), .A2(n4779), .A3(n4780), .ZN(n4778) );
  INV_X1 U6016 ( .A(n3582), .ZN(n4779) );
  INV_X1 U6017 ( .A(n4785), .ZN(n4780) );
  NOR2_X1 U6018 ( .A1(n3588), .A2(n3587), .ZN(n4782) );
  AND2_X1 U6019 ( .A1(n4436), .A2(n4446), .ZN(n4783) );
  AND2_X1 U6020 ( .A1(n4432), .A2(n4461), .ZN(n4784) );
  AND2_X1 U6021 ( .A1(n4442), .A2(n4444), .ZN(n4786) );
  INV_X2 U6022 ( .A(n4808), .ZN(n4787) );
  NAND2_X1 U6023 ( .A1(n2514), .A2(n4793), .ZN(n2533) );
  NAND2_X1 U6024 ( .A1(n4788), .A2(n2553), .ZN(n2486) );
  NOR2_X1 U6025 ( .A1(n2533), .A2(n4534), .ZN(n4788) );
  NAND2_X1 U6026 ( .A1(n4791), .A2(n2500), .ZN(n4789) );
  INV_X1 U6027 ( .A(n4792), .ZN(n4791) );
  INV_X1 U6028 ( .A(n4794), .ZN(n4793) );
  NOR2_X1 U6029 ( .A1(n2569), .A2(n224), .ZN(n4794) );
  AND2_X1 U6030 ( .A1(n4316), .A2(n4795), .ZN(n4390) );
  AND2_X1 U6031 ( .A1(n4316), .A2(n4799), .ZN(n4853) );
  AND2_X1 U6032 ( .A1(n4316), .A2(n4847), .ZN(n4854) );
  NOR2_X2 U6033 ( .A1(n4891), .A2(n4796), .ZN(n4795) );
  INV_X2 U6034 ( .A(n4797), .ZN(n4796) );
  INV_X2 U6035 ( .A(n4798), .ZN(n4797) );
  NAND2_X2 U6036 ( .A1(n4799), .A2(n4852), .ZN(n4798) );
  AND2_X2 U6037 ( .A1(n4813), .A2(n4847), .ZN(n4799) );
  INV_X2 U6038 ( .A(n4899), .ZN(n4371) );
  NAND2_X2 U6039 ( .A1(n4800), .A2(n4373), .ZN(\PC/N28 ) );
  INV_X2 U6040 ( .A(n2437), .ZN(n4802) );
  NAND2_X1 U6041 ( .A1(n4316), .A2(n4806), .ZN(n4336) );
  INV_X2 U6042 ( .A(n4804), .ZN(n4803) );
  NAND2_X2 U6043 ( .A1(n4808), .A2(n4805), .ZN(n4804) );
  INV_X2 U6044 ( .A(n4883), .ZN(n4805) );
  INV_X2 U6045 ( .A(n4807), .ZN(n4806) );
  NAND2_X2 U6046 ( .A1(n4847), .A2(n4812), .ZN(n4807) );
  NOR2_X2 U6047 ( .A1(n4809), .A2(n4811), .ZN(n4808) );
  NAND3_X1 U6048 ( .A1(n4847), .A2(n4812), .A3(n4810), .ZN(n4809) );
  INV_X2 U6049 ( .A(n4865), .ZN(n4810) );
  INV_X2 U6050 ( .A(n4861), .ZN(n4811) );
  INV_X2 U6051 ( .A(n4858), .ZN(n4812) );
  NOR2_X2 U6052 ( .A1(n4364), .A2(n4900), .ZN(n4899) );
  NOR2_X2 U6053 ( .A1(n4862), .A2(n4858), .ZN(n4813) );
  CLKBUF_X1 U6054 ( .A(n4816), .Z(n4817) );
  NAND2_X2 U6055 ( .A1(n4815), .A2(IR_OUT[21]), .ZN(n4267) );
  NAND2_X2 U6056 ( .A1(n4815), .A2(IR_OUT[25]), .ZN(n4272) );
  OR2_X2 U6057 ( .A1(n4816), .A2(n4820), .ZN(n2539) );
  INV_X2 U6058 ( .A(IR_OUT[3]), .ZN(n4820) );
  NAND2_X2 U6059 ( .A1(n4826), .A2(IR_OUT[23]), .ZN(n4269) );
  NAND2_X2 U6060 ( .A1(n4815), .A2(IR_OUT[22]), .ZN(n4268) );
  NAND2_X2 U6061 ( .A1(n4815), .A2(IR_OUT[24]), .ZN(n4270) );
  NAND2_X2 U6062 ( .A1(n4815), .A2(IR_OUT[18]), .ZN(n4421) );
  OR2_X2 U6063 ( .A1(n4817), .A2(n4821), .ZN(n2347) );
  NAND2_X2 U6064 ( .A1(IR_OUT[4]), .A2(IR_OUT[3]), .ZN(n4821) );
  NOR2_X2 U6065 ( .A1(n4823), .A2(n4817), .ZN(n4822) );
  INV_X2 U6066 ( .A(n2513), .ZN(n4823) );
  NOR2_X2 U6067 ( .A1(n4825), .A2(n4817), .ZN(n4824) );
  NOR2_X2 U6068 ( .A1(n2475), .A2(n2513), .ZN(n4825) );
  NAND2_X2 U6069 ( .A1(n4872), .A2(n4828), .ZN(n4827) );
  AND2_X2 U6070 ( .A1(n4906), .A2(n4829), .ZN(n4828) );
  AND2_X2 U6071 ( .A1(n2437), .A2(n4830), .ZN(n4829) );
  INV_X2 U6072 ( .A(n4883), .ZN(n4830) );
  INV_X2 U6073 ( .A(n4832), .ZN(n4831) );
  NAND2_X2 U6074 ( .A1(n4872), .A2(n4906), .ZN(n4832) );
  NAND2_X1 U6075 ( .A1(n4379), .A2(n4833), .ZN(n4376) );
  NAND2_X1 U6076 ( .A1(n2437), .A2(w_PC_OUT[26]), .ZN(n4834) );
  INV_X2 U6077 ( .A(n4835), .ZN(n4845) );
  NAND2_X2 U6078 ( .A1(n4884), .A2(n4837), .ZN(n4836) );
  NOR2_X2 U6079 ( .A1(n4868), .A2(n4838), .ZN(n4837) );
  NAND2_X2 U6080 ( .A1(n2437), .A2(w_PC_OUT[27]), .ZN(n4838) );
  NAND2_X2 U6081 ( .A1(n4884), .A2(n4840), .ZN(n4839) );
  INV_X2 U6082 ( .A(n4868), .ZN(n4840) );
  AND2_X2 U6083 ( .A1(n4358), .A2(n4841), .ZN(n4383) );
  INV_X2 U6084 ( .A(n4842), .ZN(n4841) );
  NAND2_X2 U6085 ( .A1(n4884), .A2(w_PC_OUT[27]), .ZN(n4842) );
  NAND2_X1 U6086 ( .A1(n4386), .A2(n4843), .ZN(n4384) );
  NAND2_X1 U6087 ( .A1(n4845), .A2(n4844), .ZN(n4843) );
  NAND2_X1 U6088 ( .A1(n2437), .A2(w_PC_OUT[28]), .ZN(n4844) );
  INV_X2 U6089 ( .A(n224), .ZN(n4846) );
  NOR2_X2 U6090 ( .A1(n4855), .A2(n4848), .ZN(n4847) );
  INV_X2 U6091 ( .A(n4849), .ZN(n4848) );
  AND2_X2 U6092 ( .A1(IROM_ADDR[9]), .A2(IROM_ADDR[10]), .ZN(n4849) );
  INV_X2 U6093 ( .A(n4387), .ZN(n4386) );
  NOR2_X2 U6094 ( .A1(n4364), .A2(n4850), .ZN(n4387) );
  OR2_X2 U6095 ( .A1(n4897), .A2(n4851), .ZN(n4850) );
  OR2_X2 U6096 ( .A1(n4896), .A2(n4900), .ZN(n4851) );
  NOR2_X2 U6097 ( .A1(n4878), .A2(n4865), .ZN(n4852) );
  NOR2_X2 U6098 ( .A1(n4322), .A2(n4857), .ZN(n4326) );
  INV_X2 U6099 ( .A(n4857), .ZN(n4856) );
  INV_X1 U6100 ( .A(n4322), .ZN(n4323) );
  INV_X2 U6101 ( .A(IROM_ADDR[11]), .ZN(n4857) );
  NAND2_X2 U6102 ( .A1(n4859), .A2(w_PC_OUT[14]), .ZN(n4858) );
  INV_X2 U6103 ( .A(n4860), .ZN(n4859) );
  INV_X2 U6104 ( .A(n4329), .ZN(n4330) );
  INV_X1 U6105 ( .A(w_PC_OUT[13]), .ZN(n4860) );
  INV_X2 U6106 ( .A(n4862), .ZN(n4861) );
  NOR2_X2 U6107 ( .A1(n4336), .A2(n4864), .ZN(n4340) );
  NAND2_X2 U6108 ( .A1(n4863), .A2(w_PC_OUT[16]), .ZN(n4862) );
  INV_X2 U6109 ( .A(n4864), .ZN(n4863) );
  INV_X1 U6110 ( .A(n4336), .ZN(n4337) );
  INV_X2 U6111 ( .A(w_PC_OUT[15]), .ZN(n4864) );
  NAND2_X2 U6112 ( .A1(n4866), .A2(w_PC_OUT[18]), .ZN(n4865) );
  INV_X2 U6113 ( .A(n4867), .ZN(n4866) );
  INV_X2 U6114 ( .A(n4343), .ZN(n4344) );
  INV_X1 U6115 ( .A(w_PC_OUT[17]), .ZN(n4867) );
  INV_X2 U6116 ( .A(n4870), .ZN(n4868) );
  NAND2_X2 U6117 ( .A1(n4874), .A2(n4870), .ZN(n4869) );
  AND2_X2 U6118 ( .A1(n4873), .A2(n4871), .ZN(n4870) );
  INV_X2 U6119 ( .A(n4883), .ZN(n4871) );
  AND2_X2 U6120 ( .A1(n4875), .A2(n4873), .ZN(n4872) );
  INV_X2 U6121 ( .A(n4877), .ZN(n4873) );
  AND2_X2 U6122 ( .A1(n4903), .A2(n4875), .ZN(n4874) );
  INV_X2 U6123 ( .A(n4876), .ZN(n4875) );
  INV_X2 U6124 ( .A(n4885), .ZN(n4876) );
  INV_X2 U6125 ( .A(n4881), .ZN(n4877) );
  NAND2_X2 U6126 ( .A1(n4880), .A2(n4879), .ZN(n4878) );
  INV_X2 U6127 ( .A(n4883), .ZN(n4879) );
  AND2_X2 U6128 ( .A1(n4881), .A2(n4888), .ZN(n4880) );
  INV_X2 U6129 ( .A(n4882), .ZN(n4881) );
  INV_X1 U6130 ( .A(n4531), .ZN(n4351) );
  INV_X2 U6131 ( .A(w_PC_OUT[20]), .ZN(n4882) );
  INV_X2 U6132 ( .A(w_PC_OUT[19]), .ZN(n4883) );
  AND2_X2 U6133 ( .A1(n4904), .A2(n4885), .ZN(n4884) );
  INV_X2 U6134 ( .A(n4886), .ZN(n4885) );
  NAND2_X2 U6135 ( .A1(n4888), .A2(n4887), .ZN(n4886) );
  INV_X2 U6136 ( .A(n4902), .ZN(n4887) );
  AND2_X2 U6137 ( .A1(w_PC_OUT[21]), .A2(w_PC_OUT[22]), .ZN(n4888) );
  INV_X2 U6138 ( .A(n4358), .ZN(n4357) );
  NAND2_X1 U6139 ( .A1(n4393), .A2(n4889), .ZN(n4392) );
  INV_X1 U6140 ( .A(n4890), .ZN(n4889) );
  NOR2_X1 U6141 ( .A1(n4390), .A2(w_PC_OUT[30]), .ZN(n4890) );
  NAND2_X2 U6142 ( .A1(n4893), .A2(n4892), .ZN(n4891) );
  NOR2_X2 U6143 ( .A1(n4894), .A2(n4902), .ZN(n4892) );
  INV_X2 U6144 ( .A(n4895), .ZN(n4893) );
  INV_X2 U6145 ( .A(n4912), .ZN(n4894) );
  INV_X2 U6146 ( .A(n4904), .ZN(n4895) );
  INV_X1 U6147 ( .A(w_PC_OUT[25]), .ZN(n4896) );
  INV_X1 U6148 ( .A(n4898), .ZN(n4897) );
  NAND2_X2 U6149 ( .A1(n4901), .A2(w_PC_OUT[24]), .ZN(n4900) );
  INV_X2 U6150 ( .A(n4902), .ZN(n4901) );
  INV_X2 U6151 ( .A(n4364), .ZN(n4365) );
  INV_X1 U6152 ( .A(w_PC_OUT[23]), .ZN(n4902) );
  AND2_X2 U6153 ( .A1(n4910), .A2(n4904), .ZN(n4903) );
  INV_X2 U6154 ( .A(n4905), .ZN(n4904) );
  NAND2_X2 U6155 ( .A1(n4906), .A2(n4908), .ZN(n4905) );
  INV_X2 U6156 ( .A(w_PC_OUT[24]), .ZN(n4907) );
  INV_X2 U6157 ( .A(w_PC_OUT[26]), .ZN(n4909) );
  INV_X2 U6158 ( .A(n4380), .ZN(n4379) );
  INV_X2 U6159 ( .A(n4911), .ZN(n4910) );
  NAND2_X2 U6160 ( .A1(n4912), .A2(w_PC_OUT[30]), .ZN(n4911) );
  INV_X2 U6161 ( .A(n4913), .ZN(n4912) );
  NAND2_X2 U6162 ( .A1(n4914), .A2(w_PC_OUT[29]), .ZN(n4913) );
  INV_X1 U6163 ( .A(n4406), .ZN(n4410) );
  NAND2_X1 U6164 ( .A1(n4916), .A2(n4915), .ZN(n4406) );
  INV_X1 U6165 ( .A(n4399), .ZN(n4915) );
  NOR2_X2 U6166 ( .A1(n4560), .A2(n4918), .ZN(n4407) );
  NOR2_X2 U6167 ( .A1(n4918), .A2(n4917), .ZN(n4916) );
  INV_X2 U6168 ( .A(n4560), .ZN(n4403) );
  INV_X1 U6169 ( .A(IROM_ADDR[3]), .ZN(n4918) );
endmodule

